module Rob(
  input         clk,
  input         reset,
  input         io_dis_valids_0,
  input         io_dis_valids_1,
  input         io_dis_uops_0_valid,
  input  [1:0]  io_dis_uops_0_iw_state,
  input  [8:0]  io_dis_uops_0_uopc,
  input  [31:0] io_dis_uops_0_inst,
  input  [39:0] io_dis_uops_0_pc,
  input  [7:0]  io_dis_uops_0_fu_code,
  input  [3:0]  io_dis_uops_0_ctrl_br_type,
  input  [1:0]  io_dis_uops_0_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_0_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_0_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_0_ctrl_op_fcn,
  input         io_dis_uops_0_ctrl_fcn_dw,
  input         io_dis_uops_0_ctrl_rf_wen,
  input  [2:0]  io_dis_uops_0_ctrl_csr_cmd,
  input         io_dis_uops_0_ctrl_is_load,
  input         io_dis_uops_0_ctrl_is_sta,
  input         io_dis_uops_0_ctrl_is_std,
  input  [1:0]  io_dis_uops_0_wakeup_delay,
  input         io_dis_uops_0_allocate_brtag,
  input         io_dis_uops_0_is_br_or_jmp,
  input         io_dis_uops_0_is_jump,
  input         io_dis_uops_0_is_jal,
  input         io_dis_uops_0_is_ret,
  input         io_dis_uops_0_is_call,
  input  [7:0]  io_dis_uops_0_br_mask,
  input  [2:0]  io_dis_uops_0_br_tag,
  input         io_dis_uops_0_br_prediction_bpd_predict_val,
  input         io_dis_uops_0_br_prediction_bpd_predict_taken,
  input         io_dis_uops_0_br_prediction_btb_hit,
  input         io_dis_uops_0_br_prediction_btb_predicted,
  input         io_dis_uops_0_br_prediction_is_br_or_jalr,
  input         io_dis_uops_0_stat_brjmp_mispredicted,
  input         io_dis_uops_0_stat_btb_made_pred,
  input         io_dis_uops_0_stat_btb_mispredicted,
  input         io_dis_uops_0_stat_bpd_made_pred,
  input         io_dis_uops_0_stat_bpd_mispredicted,
  input  [2:0]  io_dis_uops_0_fetch_pc_lob,
  input  [19:0] io_dis_uops_0_imm_packed,
  input  [11:0] io_dis_uops_0_csr_addr,
  input  [5:0]  io_dis_uops_0_rob_idx,
  input  [3:0]  io_dis_uops_0_ldq_idx,
  input  [3:0]  io_dis_uops_0_stq_idx,
  input  [4:0]  io_dis_uops_0_brob_idx,
  input  [6:0]  io_dis_uops_0_pdst,
  input  [6:0]  io_dis_uops_0_pop1,
  input  [6:0]  io_dis_uops_0_pop2,
  input  [6:0]  io_dis_uops_0_pop3,
  input         io_dis_uops_0_prs1_busy,
  input         io_dis_uops_0_prs2_busy,
  input         io_dis_uops_0_prs3_busy,
  input  [6:0]  io_dis_uops_0_stale_pdst,
  input         io_dis_uops_0_exception,
  input  [63:0] io_dis_uops_0_exc_cause,
  input         io_dis_uops_0_bypassable,
  input  [3:0]  io_dis_uops_0_mem_cmd,
  input  [2:0]  io_dis_uops_0_mem_typ,
  input         io_dis_uops_0_is_fence,
  input         io_dis_uops_0_is_fencei,
  input         io_dis_uops_0_is_store,
  input         io_dis_uops_0_is_amo,
  input         io_dis_uops_0_is_load,
  input         io_dis_uops_0_is_unique,
  input         io_dis_uops_0_flush_on_commit,
  input  [5:0]  io_dis_uops_0_ldst,
  input  [5:0]  io_dis_uops_0_lrs1,
  input  [5:0]  io_dis_uops_0_lrs2,
  input  [5:0]  io_dis_uops_0_lrs3,
  input         io_dis_uops_0_ldst_val,
  input  [1:0]  io_dis_uops_0_dst_rtype,
  input  [1:0]  io_dis_uops_0_lrs1_rtype,
  input  [1:0]  io_dis_uops_0_lrs2_rtype,
  input         io_dis_uops_0_frs3_en,
  input         io_dis_uops_0_fp_val,
  input         io_dis_uops_0_fp_single,
  input         io_dis_uops_0_xcpt_if,
  input         io_dis_uops_0_replay_if,
  input  [63:0] io_dis_uops_0_debug_wdata,
  input  [31:0] io_dis_uops_0_debug_events_fetch_seq,
  input         io_dis_uops_1_valid,
  input  [1:0]  io_dis_uops_1_iw_state,
  input  [8:0]  io_dis_uops_1_uopc,
  input  [31:0] io_dis_uops_1_inst,
  input  [39:0] io_dis_uops_1_pc,
  input  [7:0]  io_dis_uops_1_fu_code,
  input  [3:0]  io_dis_uops_1_ctrl_br_type,
  input  [1:0]  io_dis_uops_1_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_1_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_1_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_1_ctrl_op_fcn,
  input         io_dis_uops_1_ctrl_fcn_dw,
  input         io_dis_uops_1_ctrl_rf_wen,
  input  [2:0]  io_dis_uops_1_ctrl_csr_cmd,
  input         io_dis_uops_1_ctrl_is_load,
  input         io_dis_uops_1_ctrl_is_sta,
  input         io_dis_uops_1_ctrl_is_std,
  input  [1:0]  io_dis_uops_1_wakeup_delay,
  input         io_dis_uops_1_allocate_brtag,
  input         io_dis_uops_1_is_br_or_jmp,
  input         io_dis_uops_1_is_jump,
  input         io_dis_uops_1_is_jal,
  input         io_dis_uops_1_is_ret,
  input         io_dis_uops_1_is_call,
  input  [7:0]  io_dis_uops_1_br_mask,
  input  [2:0]  io_dis_uops_1_br_tag,
  input         io_dis_uops_1_br_prediction_bpd_predict_val,
  input         io_dis_uops_1_br_prediction_bpd_predict_taken,
  input         io_dis_uops_1_br_prediction_btb_hit,
  input         io_dis_uops_1_br_prediction_btb_predicted,
  input         io_dis_uops_1_br_prediction_is_br_or_jalr,
  input         io_dis_uops_1_stat_brjmp_mispredicted,
  input         io_dis_uops_1_stat_btb_made_pred,
  input         io_dis_uops_1_stat_btb_mispredicted,
  input         io_dis_uops_1_stat_bpd_made_pred,
  input         io_dis_uops_1_stat_bpd_mispredicted,
  input  [2:0]  io_dis_uops_1_fetch_pc_lob,
  input  [19:0] io_dis_uops_1_imm_packed,
  input  [11:0] io_dis_uops_1_csr_addr,
  input  [5:0]  io_dis_uops_1_rob_idx,
  input  [3:0]  io_dis_uops_1_ldq_idx,
  input  [3:0]  io_dis_uops_1_stq_idx,
  input  [4:0]  io_dis_uops_1_brob_idx,
  input  [6:0]  io_dis_uops_1_pdst,
  input  [6:0]  io_dis_uops_1_pop1,
  input  [6:0]  io_dis_uops_1_pop2,
  input  [6:0]  io_dis_uops_1_pop3,
  input         io_dis_uops_1_prs1_busy,
  input         io_dis_uops_1_prs2_busy,
  input         io_dis_uops_1_prs3_busy,
  input  [6:0]  io_dis_uops_1_stale_pdst,
  input         io_dis_uops_1_exception,
  input  [63:0] io_dis_uops_1_exc_cause,
  input         io_dis_uops_1_bypassable,
  input  [3:0]  io_dis_uops_1_mem_cmd,
  input  [2:0]  io_dis_uops_1_mem_typ,
  input         io_dis_uops_1_is_fence,
  input         io_dis_uops_1_is_fencei,
  input         io_dis_uops_1_is_store,
  input         io_dis_uops_1_is_amo,
  input         io_dis_uops_1_is_load,
  input         io_dis_uops_1_is_unique,
  input         io_dis_uops_1_flush_on_commit,
  input  [5:0]  io_dis_uops_1_ldst,
  input  [5:0]  io_dis_uops_1_lrs1,
  input  [5:0]  io_dis_uops_1_lrs2,
  input  [5:0]  io_dis_uops_1_lrs3,
  input         io_dis_uops_1_ldst_val,
  input  [1:0]  io_dis_uops_1_dst_rtype,
  input  [1:0]  io_dis_uops_1_lrs1_rtype,
  input  [1:0]  io_dis_uops_1_lrs2_rtype,
  input         io_dis_uops_1_frs3_en,
  input         io_dis_uops_1_fp_val,
  input         io_dis_uops_1_fp_single,
  input         io_dis_uops_1_xcpt_if,
  input         io_dis_uops_1_replay_if,
  input  [63:0] io_dis_uops_1_debug_wdata,
  input  [31:0] io_dis_uops_1_debug_events_fetch_seq,
  input         io_dis_has_br_or_jalr_in_packet,
  input         io_dis_partial_stall,
  input         io_dis_new_packet,
  output [5:0]  io_curr_rob_tail,
  input         io_wb_resps_0_valid,
  input         io_wb_resps_0_bits_uop_valid,
  input  [1:0]  io_wb_resps_0_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_0_bits_uop_uopc,
  input  [31:0] io_wb_resps_0_bits_uop_inst,
  input  [39:0] io_wb_resps_0_bits_uop_pc,
  input  [7:0]  io_wb_resps_0_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_0_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_0_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_0_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_0_bits_uop_ctrl_is_load,
  input         io_wb_resps_0_bits_uop_ctrl_is_sta,
  input         io_wb_resps_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_0_bits_uop_wakeup_delay,
  input         io_wb_resps_0_bits_uop_allocate_brtag,
  input         io_wb_resps_0_bits_uop_is_br_or_jmp,
  input         io_wb_resps_0_bits_uop_is_jump,
  input         io_wb_resps_0_bits_uop_is_jal,
  input         io_wb_resps_0_bits_uop_is_ret,
  input         io_wb_resps_0_bits_uop_is_call,
  input  [7:0]  io_wb_resps_0_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_0_bits_uop_br_tag,
  input         io_wb_resps_0_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_0_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_0_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_0_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_0_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_0_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_0_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_0_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_0_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_0_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_0_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_0_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_0_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_0_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_0_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_0_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_0_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_0_bits_uop_pdst,
  input  [6:0]  io_wb_resps_0_bits_uop_pop1,
  input  [6:0]  io_wb_resps_0_bits_uop_pop2,
  input  [6:0]  io_wb_resps_0_bits_uop_pop3,
  input         io_wb_resps_0_bits_uop_prs1_busy,
  input         io_wb_resps_0_bits_uop_prs2_busy,
  input         io_wb_resps_0_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_0_bits_uop_stale_pdst,
  input         io_wb_resps_0_bits_uop_exception,
  input  [63:0] io_wb_resps_0_bits_uop_exc_cause,
  input         io_wb_resps_0_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_0_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_0_bits_uop_mem_typ,
  input         io_wb_resps_0_bits_uop_is_fence,
  input         io_wb_resps_0_bits_uop_is_fencei,
  input         io_wb_resps_0_bits_uop_is_store,
  input         io_wb_resps_0_bits_uop_is_amo,
  input         io_wb_resps_0_bits_uop_is_load,
  input         io_wb_resps_0_bits_uop_is_unique,
  input         io_wb_resps_0_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_0_bits_uop_ldst,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs3,
  input         io_wb_resps_0_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_0_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_0_bits_uop_lrs2_rtype,
  input         io_wb_resps_0_bits_uop_frs3_en,
  input         io_wb_resps_0_bits_uop_fp_val,
  input         io_wb_resps_0_bits_uop_fp_single,
  input         io_wb_resps_0_bits_uop_xcpt_if,
  input         io_wb_resps_0_bits_uop_replay_if,
  input  [63:0] io_wb_resps_0_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_0_bits_uop_debug_events_fetch_seq,
  input  [64:0] io_wb_resps_0_bits_data,
  input         io_wb_resps_0_bits_fflags_valid,
  input         io_wb_resps_0_bits_fflags_bits_uop_valid,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_0_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_0_bits_fflags_bits_uop_inst,
  input  [39:0] io_wb_resps_0_bits_fflags_bits_uop_pc,
  input  [7:0]  io_wb_resps_0_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_wakeup_delay,
  input         io_wb_resps_0_bits_fflags_bits_uop_allocate_brtag,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_br_or_jmp,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_jump,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_ret,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_call,
  input  [7:0]  io_wb_resps_0_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_br_tag,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_0_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_0_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pop1,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pop2,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pop3,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_0_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_0_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_0_bits_fflags_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_mem_typ,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_store,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_load,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_0_bits_fflags_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_0_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_0_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_0_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_0_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_0_bits_fflags_bits_uop_xcpt_if,
  input         io_wb_resps_0_bits_fflags_bits_uop_replay_if,
  input  [63:0] io_wb_resps_0_bits_fflags_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_0_bits_fflags_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_flags,
  input         io_wb_resps_1_valid,
  input         io_wb_resps_1_bits_uop_valid,
  input  [1:0]  io_wb_resps_1_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_1_bits_uop_uopc,
  input  [31:0] io_wb_resps_1_bits_uop_inst,
  input  [39:0] io_wb_resps_1_bits_uop_pc,
  input  [7:0]  io_wb_resps_1_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_1_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_1_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_1_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_1_bits_uop_ctrl_is_load,
  input         io_wb_resps_1_bits_uop_ctrl_is_sta,
  input         io_wb_resps_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_1_bits_uop_wakeup_delay,
  input         io_wb_resps_1_bits_uop_allocate_brtag,
  input         io_wb_resps_1_bits_uop_is_br_or_jmp,
  input         io_wb_resps_1_bits_uop_is_jump,
  input         io_wb_resps_1_bits_uop_is_jal,
  input         io_wb_resps_1_bits_uop_is_ret,
  input         io_wb_resps_1_bits_uop_is_call,
  input  [7:0]  io_wb_resps_1_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_1_bits_uop_br_tag,
  input         io_wb_resps_1_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_1_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_1_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_1_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_1_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_1_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_1_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_1_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_1_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_1_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_1_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_1_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_1_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_1_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_1_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_1_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_1_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_1_bits_uop_pdst,
  input  [6:0]  io_wb_resps_1_bits_uop_pop1,
  input  [6:0]  io_wb_resps_1_bits_uop_pop2,
  input  [6:0]  io_wb_resps_1_bits_uop_pop3,
  input         io_wb_resps_1_bits_uop_prs1_busy,
  input         io_wb_resps_1_bits_uop_prs2_busy,
  input         io_wb_resps_1_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_1_bits_uop_stale_pdst,
  input         io_wb_resps_1_bits_uop_exception,
  input  [63:0] io_wb_resps_1_bits_uop_exc_cause,
  input         io_wb_resps_1_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_1_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_1_bits_uop_mem_typ,
  input         io_wb_resps_1_bits_uop_is_fence,
  input         io_wb_resps_1_bits_uop_is_fencei,
  input         io_wb_resps_1_bits_uop_is_store,
  input         io_wb_resps_1_bits_uop_is_amo,
  input         io_wb_resps_1_bits_uop_is_load,
  input         io_wb_resps_1_bits_uop_is_unique,
  input         io_wb_resps_1_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_1_bits_uop_ldst,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs3,
  input         io_wb_resps_1_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_1_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_1_bits_uop_lrs2_rtype,
  input         io_wb_resps_1_bits_uop_frs3_en,
  input         io_wb_resps_1_bits_uop_fp_val,
  input         io_wb_resps_1_bits_uop_fp_single,
  input         io_wb_resps_1_bits_uop_xcpt_if,
  input         io_wb_resps_1_bits_uop_replay_if,
  input  [63:0] io_wb_resps_1_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_1_bits_uop_debug_events_fetch_seq,
  input  [64:0] io_wb_resps_1_bits_data,
  input         io_wb_resps_1_bits_fflags_valid,
  input         io_wb_resps_1_bits_fflags_bits_uop_valid,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_1_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_1_bits_fflags_bits_uop_inst,
  input  [39:0] io_wb_resps_1_bits_fflags_bits_uop_pc,
  input  [7:0]  io_wb_resps_1_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_wakeup_delay,
  input         io_wb_resps_1_bits_fflags_bits_uop_allocate_brtag,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_br_or_jmp,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_jump,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_ret,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_call,
  input  [7:0]  io_wb_resps_1_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_br_tag,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_1_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_1_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pop1,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pop2,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pop3,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_1_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_1_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_1_bits_fflags_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_mem_typ,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_store,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_load,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_1_bits_fflags_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_1_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_1_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_1_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_1_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_1_bits_fflags_bits_uop_xcpt_if,
  input         io_wb_resps_1_bits_fflags_bits_uop_replay_if,
  input  [63:0] io_wb_resps_1_bits_fflags_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_1_bits_fflags_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_flags,
  input         io_wb_resps_2_valid,
  input         io_wb_resps_2_bits_uop_valid,
  input  [1:0]  io_wb_resps_2_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_2_bits_uop_uopc,
  input  [31:0] io_wb_resps_2_bits_uop_inst,
  input  [39:0] io_wb_resps_2_bits_uop_pc,
  input  [7:0]  io_wb_resps_2_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_2_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_2_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_2_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_2_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_2_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_2_bits_uop_ctrl_is_load,
  input         io_wb_resps_2_bits_uop_ctrl_is_sta,
  input         io_wb_resps_2_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_2_bits_uop_wakeup_delay,
  input         io_wb_resps_2_bits_uop_allocate_brtag,
  input         io_wb_resps_2_bits_uop_is_br_or_jmp,
  input         io_wb_resps_2_bits_uop_is_jump,
  input         io_wb_resps_2_bits_uop_is_jal,
  input         io_wb_resps_2_bits_uop_is_ret,
  input         io_wb_resps_2_bits_uop_is_call,
  input  [7:0]  io_wb_resps_2_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_2_bits_uop_br_tag,
  input         io_wb_resps_2_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_2_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_2_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_2_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_2_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_2_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_2_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_2_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_2_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_2_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_2_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_2_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_2_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_2_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_2_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_2_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_2_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_2_bits_uop_pdst,
  input  [6:0]  io_wb_resps_2_bits_uop_pop1,
  input  [6:0]  io_wb_resps_2_bits_uop_pop2,
  input  [6:0]  io_wb_resps_2_bits_uop_pop3,
  input         io_wb_resps_2_bits_uop_prs1_busy,
  input         io_wb_resps_2_bits_uop_prs2_busy,
  input         io_wb_resps_2_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_2_bits_uop_stale_pdst,
  input         io_wb_resps_2_bits_uop_exception,
  input  [63:0] io_wb_resps_2_bits_uop_exc_cause,
  input         io_wb_resps_2_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_2_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_2_bits_uop_mem_typ,
  input         io_wb_resps_2_bits_uop_is_fence,
  input         io_wb_resps_2_bits_uop_is_fencei,
  input         io_wb_resps_2_bits_uop_is_store,
  input         io_wb_resps_2_bits_uop_is_amo,
  input         io_wb_resps_2_bits_uop_is_load,
  input         io_wb_resps_2_bits_uop_is_unique,
  input         io_wb_resps_2_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_2_bits_uop_ldst,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs3,
  input         io_wb_resps_2_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_2_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_2_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_2_bits_uop_lrs2_rtype,
  input         io_wb_resps_2_bits_uop_frs3_en,
  input         io_wb_resps_2_bits_uop_fp_val,
  input         io_wb_resps_2_bits_uop_fp_single,
  input         io_wb_resps_2_bits_uop_xcpt_if,
  input         io_wb_resps_2_bits_uop_replay_if,
  input  [63:0] io_wb_resps_2_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_2_bits_uop_debug_events_fetch_seq,
  input  [64:0] io_wb_resps_2_bits_data,
  input         io_wb_resps_2_bits_fflags_valid,
  input         io_wb_resps_2_bits_fflags_bits_uop_valid,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_2_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_2_bits_fflags_bits_uop_inst,
  input  [39:0] io_wb_resps_2_bits_fflags_bits_uop_pc,
  input  [7:0]  io_wb_resps_2_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_wakeup_delay,
  input         io_wb_resps_2_bits_fflags_bits_uop_allocate_brtag,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_br_or_jmp,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_jump,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_ret,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_call,
  input  [7:0]  io_wb_resps_2_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_br_tag,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_2_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_2_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pop1,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pop2,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pop3,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_2_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_2_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_2_bits_fflags_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_mem_typ,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_store,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_load,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_2_bits_fflags_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_2_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_2_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_2_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_2_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_2_bits_fflags_bits_uop_xcpt_if,
  input         io_wb_resps_2_bits_fflags_bits_uop_replay_if,
  input  [63:0] io_wb_resps_2_bits_fflags_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_2_bits_fflags_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_flags,
  input         io_debug_wb_valids_0,
  input         io_debug_wb_valids_1,
  input         io_debug_wb_valids_2,
  input  [63:0] io_debug_wb_wdata_0,
  input  [63:0] io_debug_wb_wdata_1,
  input  [63:0] io_debug_wb_wdata_2,
  input         io_fflags_0_valid,
  input         io_fflags_0_bits_uop_valid,
  input  [1:0]  io_fflags_0_bits_uop_iw_state,
  input  [8:0]  io_fflags_0_bits_uop_uopc,
  input  [31:0] io_fflags_0_bits_uop_inst,
  input  [39:0] io_fflags_0_bits_uop_pc,
  input  [7:0]  io_fflags_0_bits_uop_fu_code,
  input  [3:0]  io_fflags_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_fflags_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_fflags_0_bits_uop_ctrl_op_fcn,
  input         io_fflags_0_bits_uop_ctrl_fcn_dw,
  input         io_fflags_0_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_csr_cmd,
  input         io_fflags_0_bits_uop_ctrl_is_load,
  input         io_fflags_0_bits_uop_ctrl_is_sta,
  input         io_fflags_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_fflags_0_bits_uop_wakeup_delay,
  input         io_fflags_0_bits_uop_allocate_brtag,
  input         io_fflags_0_bits_uop_is_br_or_jmp,
  input         io_fflags_0_bits_uop_is_jump,
  input         io_fflags_0_bits_uop_is_jal,
  input         io_fflags_0_bits_uop_is_ret,
  input         io_fflags_0_bits_uop_is_call,
  input  [7:0]  io_fflags_0_bits_uop_br_mask,
  input  [2:0]  io_fflags_0_bits_uop_br_tag,
  input         io_fflags_0_bits_uop_br_prediction_bpd_predict_val,
  input         io_fflags_0_bits_uop_br_prediction_bpd_predict_taken,
  input         io_fflags_0_bits_uop_br_prediction_btb_hit,
  input         io_fflags_0_bits_uop_br_prediction_btb_predicted,
  input         io_fflags_0_bits_uop_br_prediction_is_br_or_jalr,
  input         io_fflags_0_bits_uop_stat_brjmp_mispredicted,
  input         io_fflags_0_bits_uop_stat_btb_made_pred,
  input         io_fflags_0_bits_uop_stat_btb_mispredicted,
  input         io_fflags_0_bits_uop_stat_bpd_made_pred,
  input         io_fflags_0_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_fflags_0_bits_uop_fetch_pc_lob,
  input  [19:0] io_fflags_0_bits_uop_imm_packed,
  input  [11:0] io_fflags_0_bits_uop_csr_addr,
  input  [5:0]  io_fflags_0_bits_uop_rob_idx,
  input  [3:0]  io_fflags_0_bits_uop_ldq_idx,
  input  [3:0]  io_fflags_0_bits_uop_stq_idx,
  input  [4:0]  io_fflags_0_bits_uop_brob_idx,
  input  [6:0]  io_fflags_0_bits_uop_pdst,
  input  [6:0]  io_fflags_0_bits_uop_pop1,
  input  [6:0]  io_fflags_0_bits_uop_pop2,
  input  [6:0]  io_fflags_0_bits_uop_pop3,
  input         io_fflags_0_bits_uop_prs1_busy,
  input         io_fflags_0_bits_uop_prs2_busy,
  input         io_fflags_0_bits_uop_prs3_busy,
  input  [6:0]  io_fflags_0_bits_uop_stale_pdst,
  input         io_fflags_0_bits_uop_exception,
  input  [63:0] io_fflags_0_bits_uop_exc_cause,
  input         io_fflags_0_bits_uop_bypassable,
  input  [3:0]  io_fflags_0_bits_uop_mem_cmd,
  input  [2:0]  io_fflags_0_bits_uop_mem_typ,
  input         io_fflags_0_bits_uop_is_fence,
  input         io_fflags_0_bits_uop_is_fencei,
  input         io_fflags_0_bits_uop_is_store,
  input         io_fflags_0_bits_uop_is_amo,
  input         io_fflags_0_bits_uop_is_load,
  input         io_fflags_0_bits_uop_is_unique,
  input         io_fflags_0_bits_uop_flush_on_commit,
  input  [5:0]  io_fflags_0_bits_uop_ldst,
  input  [5:0]  io_fflags_0_bits_uop_lrs1,
  input  [5:0]  io_fflags_0_bits_uop_lrs2,
  input  [5:0]  io_fflags_0_bits_uop_lrs3,
  input         io_fflags_0_bits_uop_ldst_val,
  input  [1:0]  io_fflags_0_bits_uop_dst_rtype,
  input  [1:0]  io_fflags_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_fflags_0_bits_uop_lrs2_rtype,
  input         io_fflags_0_bits_uop_frs3_en,
  input         io_fflags_0_bits_uop_fp_val,
  input         io_fflags_0_bits_uop_fp_single,
  input         io_fflags_0_bits_uop_xcpt_if,
  input         io_fflags_0_bits_uop_replay_if,
  input  [63:0] io_fflags_0_bits_uop_debug_wdata,
  input  [31:0] io_fflags_0_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_1_valid,
  input         io_fflags_1_bits_uop_valid,
  input  [1:0]  io_fflags_1_bits_uop_iw_state,
  input  [8:0]  io_fflags_1_bits_uop_uopc,
  input  [31:0] io_fflags_1_bits_uop_inst,
  input  [39:0] io_fflags_1_bits_uop_pc,
  input  [7:0]  io_fflags_1_bits_uop_fu_code,
  input  [3:0]  io_fflags_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_fflags_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_fflags_1_bits_uop_ctrl_op_fcn,
  input         io_fflags_1_bits_uop_ctrl_fcn_dw,
  input         io_fflags_1_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_csr_cmd,
  input         io_fflags_1_bits_uop_ctrl_is_load,
  input         io_fflags_1_bits_uop_ctrl_is_sta,
  input         io_fflags_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_fflags_1_bits_uop_wakeup_delay,
  input         io_fflags_1_bits_uop_allocate_brtag,
  input         io_fflags_1_bits_uop_is_br_or_jmp,
  input         io_fflags_1_bits_uop_is_jump,
  input         io_fflags_1_bits_uop_is_jal,
  input         io_fflags_1_bits_uop_is_ret,
  input         io_fflags_1_bits_uop_is_call,
  input  [7:0]  io_fflags_1_bits_uop_br_mask,
  input  [2:0]  io_fflags_1_bits_uop_br_tag,
  input         io_fflags_1_bits_uop_br_prediction_bpd_predict_val,
  input         io_fflags_1_bits_uop_br_prediction_bpd_predict_taken,
  input         io_fflags_1_bits_uop_br_prediction_btb_hit,
  input         io_fflags_1_bits_uop_br_prediction_btb_predicted,
  input         io_fflags_1_bits_uop_br_prediction_is_br_or_jalr,
  input         io_fflags_1_bits_uop_stat_brjmp_mispredicted,
  input         io_fflags_1_bits_uop_stat_btb_made_pred,
  input         io_fflags_1_bits_uop_stat_btb_mispredicted,
  input         io_fflags_1_bits_uop_stat_bpd_made_pred,
  input         io_fflags_1_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_fflags_1_bits_uop_fetch_pc_lob,
  input  [19:0] io_fflags_1_bits_uop_imm_packed,
  input  [11:0] io_fflags_1_bits_uop_csr_addr,
  input  [5:0]  io_fflags_1_bits_uop_rob_idx,
  input  [3:0]  io_fflags_1_bits_uop_ldq_idx,
  input  [3:0]  io_fflags_1_bits_uop_stq_idx,
  input  [4:0]  io_fflags_1_bits_uop_brob_idx,
  input  [6:0]  io_fflags_1_bits_uop_pdst,
  input  [6:0]  io_fflags_1_bits_uop_pop1,
  input  [6:0]  io_fflags_1_bits_uop_pop2,
  input  [6:0]  io_fflags_1_bits_uop_pop3,
  input         io_fflags_1_bits_uop_prs1_busy,
  input         io_fflags_1_bits_uop_prs2_busy,
  input         io_fflags_1_bits_uop_prs3_busy,
  input  [6:0]  io_fflags_1_bits_uop_stale_pdst,
  input         io_fflags_1_bits_uop_exception,
  input  [63:0] io_fflags_1_bits_uop_exc_cause,
  input         io_fflags_1_bits_uop_bypassable,
  input  [3:0]  io_fflags_1_bits_uop_mem_cmd,
  input  [2:0]  io_fflags_1_bits_uop_mem_typ,
  input         io_fflags_1_bits_uop_is_fence,
  input         io_fflags_1_bits_uop_is_fencei,
  input         io_fflags_1_bits_uop_is_store,
  input         io_fflags_1_bits_uop_is_amo,
  input         io_fflags_1_bits_uop_is_load,
  input         io_fflags_1_bits_uop_is_unique,
  input         io_fflags_1_bits_uop_flush_on_commit,
  input  [5:0]  io_fflags_1_bits_uop_ldst,
  input  [5:0]  io_fflags_1_bits_uop_lrs1,
  input  [5:0]  io_fflags_1_bits_uop_lrs2,
  input  [5:0]  io_fflags_1_bits_uop_lrs3,
  input         io_fflags_1_bits_uop_ldst_val,
  input  [1:0]  io_fflags_1_bits_uop_dst_rtype,
  input  [1:0]  io_fflags_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_fflags_1_bits_uop_lrs2_rtype,
  input         io_fflags_1_bits_uop_frs3_en,
  input         io_fflags_1_bits_uop_fp_val,
  input         io_fflags_1_bits_uop_fp_single,
  input         io_fflags_1_bits_uop_xcpt_if,
  input         io_fflags_1_bits_uop_replay_if,
  input  [63:0] io_fflags_1_bits_uop_debug_wdata,
  input  [31:0] io_fflags_1_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_fflags_1_bits_flags,
  input         io_lxcpt_valid,
  input         io_lxcpt_bits_uop_valid,
  input  [1:0]  io_lxcpt_bits_uop_iw_state,
  input  [8:0]  io_lxcpt_bits_uop_uopc,
  input  [31:0] io_lxcpt_bits_uop_inst,
  input  [39:0] io_lxcpt_bits_uop_pc,
  input  [7:0]  io_lxcpt_bits_uop_fu_code,
  input  [3:0]  io_lxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_lxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_lxcpt_bits_uop_ctrl_op_fcn,
  input         io_lxcpt_bits_uop_ctrl_fcn_dw,
  input         io_lxcpt_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_csr_cmd,
  input         io_lxcpt_bits_uop_ctrl_is_load,
  input         io_lxcpt_bits_uop_ctrl_is_sta,
  input         io_lxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_lxcpt_bits_uop_wakeup_delay,
  input         io_lxcpt_bits_uop_allocate_brtag,
  input         io_lxcpt_bits_uop_is_br_or_jmp,
  input         io_lxcpt_bits_uop_is_jump,
  input         io_lxcpt_bits_uop_is_jal,
  input         io_lxcpt_bits_uop_is_ret,
  input         io_lxcpt_bits_uop_is_call,
  input  [7:0]  io_lxcpt_bits_uop_br_mask,
  input  [2:0]  io_lxcpt_bits_uop_br_tag,
  input         io_lxcpt_bits_uop_br_prediction_bpd_predict_val,
  input         io_lxcpt_bits_uop_br_prediction_bpd_predict_taken,
  input         io_lxcpt_bits_uop_br_prediction_btb_hit,
  input         io_lxcpt_bits_uop_br_prediction_btb_predicted,
  input         io_lxcpt_bits_uop_br_prediction_is_br_or_jalr,
  input         io_lxcpt_bits_uop_stat_brjmp_mispredicted,
  input         io_lxcpt_bits_uop_stat_btb_made_pred,
  input         io_lxcpt_bits_uop_stat_btb_mispredicted,
  input         io_lxcpt_bits_uop_stat_bpd_made_pred,
  input         io_lxcpt_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_lxcpt_bits_uop_fetch_pc_lob,
  input  [19:0] io_lxcpt_bits_uop_imm_packed,
  input  [11:0] io_lxcpt_bits_uop_csr_addr,
  input  [5:0]  io_lxcpt_bits_uop_rob_idx,
  input  [3:0]  io_lxcpt_bits_uop_ldq_idx,
  input  [3:0]  io_lxcpt_bits_uop_stq_idx,
  input  [4:0]  io_lxcpt_bits_uop_brob_idx,
  input  [6:0]  io_lxcpt_bits_uop_pdst,
  input  [6:0]  io_lxcpt_bits_uop_pop1,
  input  [6:0]  io_lxcpt_bits_uop_pop2,
  input  [6:0]  io_lxcpt_bits_uop_pop3,
  input         io_lxcpt_bits_uop_prs1_busy,
  input         io_lxcpt_bits_uop_prs2_busy,
  input         io_lxcpt_bits_uop_prs3_busy,
  input  [6:0]  io_lxcpt_bits_uop_stale_pdst,
  input         io_lxcpt_bits_uop_exception,
  input  [63:0] io_lxcpt_bits_uop_exc_cause,
  input         io_lxcpt_bits_uop_bypassable,
  input  [3:0]  io_lxcpt_bits_uop_mem_cmd,
  input  [2:0]  io_lxcpt_bits_uop_mem_typ,
  input         io_lxcpt_bits_uop_is_fence,
  input         io_lxcpt_bits_uop_is_fencei,
  input         io_lxcpt_bits_uop_is_store,
  input         io_lxcpt_bits_uop_is_amo,
  input         io_lxcpt_bits_uop_is_load,
  input         io_lxcpt_bits_uop_is_unique,
  input         io_lxcpt_bits_uop_flush_on_commit,
  input  [5:0]  io_lxcpt_bits_uop_ldst,
  input  [5:0]  io_lxcpt_bits_uop_lrs1,
  input  [5:0]  io_lxcpt_bits_uop_lrs2,
  input  [5:0]  io_lxcpt_bits_uop_lrs3,
  input         io_lxcpt_bits_uop_ldst_val,
  input  [1:0]  io_lxcpt_bits_uop_dst_rtype,
  input  [1:0]  io_lxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_lxcpt_bits_uop_lrs2_rtype,
  input         io_lxcpt_bits_uop_frs3_en,
  input         io_lxcpt_bits_uop_fp_val,
  input         io_lxcpt_bits_uop_fp_single,
  input         io_lxcpt_bits_uop_xcpt_if,
  input         io_lxcpt_bits_uop_replay_if,
  input  [63:0] io_lxcpt_bits_uop_debug_wdata,
  input  [31:0] io_lxcpt_bits_uop_debug_events_fetch_seq,
  input  [3:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  input         io_bxcpt_valid,
  input         io_bxcpt_bits_uop_valid,
  input  [1:0]  io_bxcpt_bits_uop_iw_state,
  input  [8:0]  io_bxcpt_bits_uop_uopc,
  input  [31:0] io_bxcpt_bits_uop_inst,
  input  [39:0] io_bxcpt_bits_uop_pc,
  input  [7:0]  io_bxcpt_bits_uop_fu_code,
  input  [3:0]  io_bxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_bxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bxcpt_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bxcpt_bits_uop_ctrl_op_fcn,
  input         io_bxcpt_bits_uop_ctrl_fcn_dw,
  input         io_bxcpt_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_bxcpt_bits_uop_ctrl_csr_cmd,
  input         io_bxcpt_bits_uop_ctrl_is_load,
  input         io_bxcpt_bits_uop_ctrl_is_sta,
  input         io_bxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_bxcpt_bits_uop_wakeup_delay,
  input         io_bxcpt_bits_uop_allocate_brtag,
  input         io_bxcpt_bits_uop_is_br_or_jmp,
  input         io_bxcpt_bits_uop_is_jump,
  input         io_bxcpt_bits_uop_is_jal,
  input         io_bxcpt_bits_uop_is_ret,
  input         io_bxcpt_bits_uop_is_call,
  input  [7:0]  io_bxcpt_bits_uop_br_mask,
  input  [2:0]  io_bxcpt_bits_uop_br_tag,
  input         io_bxcpt_bits_uop_br_prediction_bpd_predict_val,
  input         io_bxcpt_bits_uop_br_prediction_bpd_predict_taken,
  input         io_bxcpt_bits_uop_br_prediction_btb_hit,
  input         io_bxcpt_bits_uop_br_prediction_btb_predicted,
  input         io_bxcpt_bits_uop_br_prediction_is_br_or_jalr,
  input         io_bxcpt_bits_uop_stat_brjmp_mispredicted,
  input         io_bxcpt_bits_uop_stat_btb_made_pred,
  input         io_bxcpt_bits_uop_stat_btb_mispredicted,
  input         io_bxcpt_bits_uop_stat_bpd_made_pred,
  input         io_bxcpt_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_bxcpt_bits_uop_fetch_pc_lob,
  input  [19:0] io_bxcpt_bits_uop_imm_packed,
  input  [11:0] io_bxcpt_bits_uop_csr_addr,
  input  [5:0]  io_bxcpt_bits_uop_rob_idx,
  input  [3:0]  io_bxcpt_bits_uop_ldq_idx,
  input  [3:0]  io_bxcpt_bits_uop_stq_idx,
  input  [4:0]  io_bxcpt_bits_uop_brob_idx,
  input  [6:0]  io_bxcpt_bits_uop_pdst,
  input  [6:0]  io_bxcpt_bits_uop_pop1,
  input  [6:0]  io_bxcpt_bits_uop_pop2,
  input  [6:0]  io_bxcpt_bits_uop_pop3,
  input         io_bxcpt_bits_uop_prs1_busy,
  input         io_bxcpt_bits_uop_prs2_busy,
  input         io_bxcpt_bits_uop_prs3_busy,
  input  [6:0]  io_bxcpt_bits_uop_stale_pdst,
  input         io_bxcpt_bits_uop_exception,
  input  [63:0] io_bxcpt_bits_uop_exc_cause,
  input         io_bxcpt_bits_uop_bypassable,
  input  [3:0]  io_bxcpt_bits_uop_mem_cmd,
  input  [2:0]  io_bxcpt_bits_uop_mem_typ,
  input         io_bxcpt_bits_uop_is_fence,
  input         io_bxcpt_bits_uop_is_fencei,
  input         io_bxcpt_bits_uop_is_store,
  input         io_bxcpt_bits_uop_is_amo,
  input         io_bxcpt_bits_uop_is_load,
  input         io_bxcpt_bits_uop_is_unique,
  input         io_bxcpt_bits_uop_flush_on_commit,
  input  [5:0]  io_bxcpt_bits_uop_ldst,
  input  [5:0]  io_bxcpt_bits_uop_lrs1,
  input  [5:0]  io_bxcpt_bits_uop_lrs2,
  input  [5:0]  io_bxcpt_bits_uop_lrs3,
  input         io_bxcpt_bits_uop_ldst_val,
  input  [1:0]  io_bxcpt_bits_uop_dst_rtype,
  input  [1:0]  io_bxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_bxcpt_bits_uop_lrs2_rtype,
  input         io_bxcpt_bits_uop_frs3_en,
  input         io_bxcpt_bits_uop_fp_val,
  input         io_bxcpt_bits_uop_fp_single,
  input         io_bxcpt_bits_uop_xcpt_if,
  input         io_bxcpt_bits_uop_replay_if,
  input  [63:0] io_bxcpt_bits_uop_debug_wdata,
  input  [31:0] io_bxcpt_bits_uop_debug_events_fetch_seq,
  input  [3:0]  io_bxcpt_bits_cause,
  input  [39:0] io_bxcpt_bits_badvaddr,
  input         io_cxcpt_valid,
  input         io_cxcpt_bits_uop_valid,
  input  [1:0]  io_cxcpt_bits_uop_iw_state,
  input  [8:0]  io_cxcpt_bits_uop_uopc,
  input  [31:0] io_cxcpt_bits_uop_inst,
  input  [39:0] io_cxcpt_bits_uop_pc,
  input  [7:0]  io_cxcpt_bits_uop_fu_code,
  input  [3:0]  io_cxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_cxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_cxcpt_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_cxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_cxcpt_bits_uop_ctrl_op_fcn,
  input         io_cxcpt_bits_uop_ctrl_fcn_dw,
  input         io_cxcpt_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_cxcpt_bits_uop_ctrl_csr_cmd,
  input         io_cxcpt_bits_uop_ctrl_is_load,
  input         io_cxcpt_bits_uop_ctrl_is_sta,
  input         io_cxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_cxcpt_bits_uop_wakeup_delay,
  input         io_cxcpt_bits_uop_allocate_brtag,
  input         io_cxcpt_bits_uop_is_br_or_jmp,
  input         io_cxcpt_bits_uop_is_jump,
  input         io_cxcpt_bits_uop_is_jal,
  input         io_cxcpt_bits_uop_is_ret,
  input         io_cxcpt_bits_uop_is_call,
  input  [7:0]  io_cxcpt_bits_uop_br_mask,
  input  [2:0]  io_cxcpt_bits_uop_br_tag,
  input         io_cxcpt_bits_uop_br_prediction_bpd_predict_val,
  input         io_cxcpt_bits_uop_br_prediction_bpd_predict_taken,
  input         io_cxcpt_bits_uop_br_prediction_btb_hit,
  input         io_cxcpt_bits_uop_br_prediction_btb_predicted,
  input         io_cxcpt_bits_uop_br_prediction_is_br_or_jalr,
  input         io_cxcpt_bits_uop_stat_brjmp_mispredicted,
  input         io_cxcpt_bits_uop_stat_btb_made_pred,
  input         io_cxcpt_bits_uop_stat_btb_mispredicted,
  input         io_cxcpt_bits_uop_stat_bpd_made_pred,
  input         io_cxcpt_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_cxcpt_bits_uop_fetch_pc_lob,
  input  [19:0] io_cxcpt_bits_uop_imm_packed,
  input  [11:0] io_cxcpt_bits_uop_csr_addr,
  input  [5:0]  io_cxcpt_bits_uop_rob_idx,
  input  [3:0]  io_cxcpt_bits_uop_ldq_idx,
  input  [3:0]  io_cxcpt_bits_uop_stq_idx,
  input  [4:0]  io_cxcpt_bits_uop_brob_idx,
  input  [6:0]  io_cxcpt_bits_uop_pdst,
  input  [6:0]  io_cxcpt_bits_uop_pop1,
  input  [6:0]  io_cxcpt_bits_uop_pop2,
  input  [6:0]  io_cxcpt_bits_uop_pop3,
  input         io_cxcpt_bits_uop_prs1_busy,
  input         io_cxcpt_bits_uop_prs2_busy,
  input         io_cxcpt_bits_uop_prs3_busy,
  input  [6:0]  io_cxcpt_bits_uop_stale_pdst,
  input         io_cxcpt_bits_uop_exception,
  input  [63:0] io_cxcpt_bits_uop_exc_cause,
  input         io_cxcpt_bits_uop_bypassable,
  input  [3:0]  io_cxcpt_bits_uop_mem_cmd,
  input  [2:0]  io_cxcpt_bits_uop_mem_typ,
  input         io_cxcpt_bits_uop_is_fence,
  input         io_cxcpt_bits_uop_is_fencei,
  input         io_cxcpt_bits_uop_is_store,
  input         io_cxcpt_bits_uop_is_amo,
  input         io_cxcpt_bits_uop_is_load,
  input         io_cxcpt_bits_uop_is_unique,
  input         io_cxcpt_bits_uop_flush_on_commit,
  input  [5:0]  io_cxcpt_bits_uop_ldst,
  input  [5:0]  io_cxcpt_bits_uop_lrs1,
  input  [5:0]  io_cxcpt_bits_uop_lrs2,
  input  [5:0]  io_cxcpt_bits_uop_lrs3,
  input         io_cxcpt_bits_uop_ldst_val,
  input  [1:0]  io_cxcpt_bits_uop_dst_rtype,
  input  [1:0]  io_cxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_cxcpt_bits_uop_lrs2_rtype,
  input         io_cxcpt_bits_uop_frs3_en,
  input         io_cxcpt_bits_uop_fp_val,
  input         io_cxcpt_bits_uop_fp_single,
  input         io_cxcpt_bits_uop_xcpt_if,
  input         io_cxcpt_bits_uop_replay_if,
  input  [63:0] io_cxcpt_bits_uop_debug_wdata,
  input  [31:0] io_cxcpt_bits_uop_debug_events_fetch_seq,
  input  [3:0]  io_cxcpt_bits_cause,
  input  [39:0] io_cxcpt_bits_badvaddr,
  output        io_com_valids_0,
  output        io_com_valids_1,
  output        io_com_uops_0_valid,
  output [1:0]  io_com_uops_0_iw_state,
  output [8:0]  io_com_uops_0_uopc,
  output [31:0] io_com_uops_0_inst,
  output [39:0] io_com_uops_0_pc,
  output [7:0]  io_com_uops_0_fu_code,
  output [3:0]  io_com_uops_0_ctrl_br_type,
  output [1:0]  io_com_uops_0_ctrl_op1_sel,
  output [2:0]  io_com_uops_0_ctrl_op2_sel,
  output [2:0]  io_com_uops_0_ctrl_imm_sel,
  output [3:0]  io_com_uops_0_ctrl_op_fcn,
  output        io_com_uops_0_ctrl_fcn_dw,
  output        io_com_uops_0_ctrl_rf_wen,
  output [2:0]  io_com_uops_0_ctrl_csr_cmd,
  output        io_com_uops_0_ctrl_is_load,
  output        io_com_uops_0_ctrl_is_sta,
  output        io_com_uops_0_ctrl_is_std,
  output [1:0]  io_com_uops_0_wakeup_delay,
  output        io_com_uops_0_allocate_brtag,
  output        io_com_uops_0_is_br_or_jmp,
  output        io_com_uops_0_is_jump,
  output        io_com_uops_0_is_jal,
  output        io_com_uops_0_is_ret,
  output        io_com_uops_0_is_call,
  output [7:0]  io_com_uops_0_br_mask,
  output [2:0]  io_com_uops_0_br_tag,
  output        io_com_uops_0_br_prediction_bpd_predict_val,
  output        io_com_uops_0_br_prediction_bpd_predict_taken,
  output        io_com_uops_0_br_prediction_btb_hit,
  output        io_com_uops_0_br_prediction_btb_predicted,
  output        io_com_uops_0_br_prediction_is_br_or_jalr,
  output        io_com_uops_0_stat_brjmp_mispredicted,
  output        io_com_uops_0_stat_btb_made_pred,
  output        io_com_uops_0_stat_btb_mispredicted,
  output        io_com_uops_0_stat_bpd_made_pred,
  output        io_com_uops_0_stat_bpd_mispredicted,
  output [2:0]  io_com_uops_0_fetch_pc_lob,
  output [19:0] io_com_uops_0_imm_packed,
  output [11:0] io_com_uops_0_csr_addr,
  output [5:0]  io_com_uops_0_rob_idx,
  output [3:0]  io_com_uops_0_ldq_idx,
  output [3:0]  io_com_uops_0_stq_idx,
  output [4:0]  io_com_uops_0_brob_idx,
  output [6:0]  io_com_uops_0_pdst,
  output [6:0]  io_com_uops_0_pop1,
  output [6:0]  io_com_uops_0_pop2,
  output [6:0]  io_com_uops_0_pop3,
  output        io_com_uops_0_prs1_busy,
  output        io_com_uops_0_prs2_busy,
  output        io_com_uops_0_prs3_busy,
  output [6:0]  io_com_uops_0_stale_pdst,
  output        io_com_uops_0_exception,
  output [63:0] io_com_uops_0_exc_cause,
  output        io_com_uops_0_bypassable,
  output [3:0]  io_com_uops_0_mem_cmd,
  output [2:0]  io_com_uops_0_mem_typ,
  output        io_com_uops_0_is_fence,
  output        io_com_uops_0_is_fencei,
  output        io_com_uops_0_is_store,
  output        io_com_uops_0_is_amo,
  output        io_com_uops_0_is_load,
  output        io_com_uops_0_is_unique,
  output        io_com_uops_0_flush_on_commit,
  output [5:0]  io_com_uops_0_ldst,
  output [5:0]  io_com_uops_0_lrs1,
  output [5:0]  io_com_uops_0_lrs2,
  output [5:0]  io_com_uops_0_lrs3,
  output        io_com_uops_0_ldst_val,
  output [1:0]  io_com_uops_0_dst_rtype,
  output [1:0]  io_com_uops_0_lrs1_rtype,
  output [1:0]  io_com_uops_0_lrs2_rtype,
  output        io_com_uops_0_frs3_en,
  output        io_com_uops_0_fp_val,
  output        io_com_uops_0_fp_single,
  output        io_com_uops_0_xcpt_if,
  output        io_com_uops_0_replay_if,
  output [63:0] io_com_uops_0_debug_wdata,
  output [31:0] io_com_uops_0_debug_events_fetch_seq,
  output        io_com_uops_1_valid,
  output [1:0]  io_com_uops_1_iw_state,
  output [8:0]  io_com_uops_1_uopc,
  output [31:0] io_com_uops_1_inst,
  output [39:0] io_com_uops_1_pc,
  output [7:0]  io_com_uops_1_fu_code,
  output [3:0]  io_com_uops_1_ctrl_br_type,
  output [1:0]  io_com_uops_1_ctrl_op1_sel,
  output [2:0]  io_com_uops_1_ctrl_op2_sel,
  output [2:0]  io_com_uops_1_ctrl_imm_sel,
  output [3:0]  io_com_uops_1_ctrl_op_fcn,
  output        io_com_uops_1_ctrl_fcn_dw,
  output        io_com_uops_1_ctrl_rf_wen,
  output [2:0]  io_com_uops_1_ctrl_csr_cmd,
  output        io_com_uops_1_ctrl_is_load,
  output        io_com_uops_1_ctrl_is_sta,
  output        io_com_uops_1_ctrl_is_std,
  output [1:0]  io_com_uops_1_wakeup_delay,
  output        io_com_uops_1_allocate_brtag,
  output        io_com_uops_1_is_br_or_jmp,
  output        io_com_uops_1_is_jump,
  output        io_com_uops_1_is_jal,
  output        io_com_uops_1_is_ret,
  output        io_com_uops_1_is_call,
  output [7:0]  io_com_uops_1_br_mask,
  output [2:0]  io_com_uops_1_br_tag,
  output        io_com_uops_1_br_prediction_bpd_predict_val,
  output        io_com_uops_1_br_prediction_bpd_predict_taken,
  output        io_com_uops_1_br_prediction_btb_hit,
  output        io_com_uops_1_br_prediction_btb_predicted,
  output        io_com_uops_1_br_prediction_is_br_or_jalr,
  output        io_com_uops_1_stat_brjmp_mispredicted,
  output        io_com_uops_1_stat_btb_made_pred,
  output        io_com_uops_1_stat_btb_mispredicted,
  output        io_com_uops_1_stat_bpd_made_pred,
  output        io_com_uops_1_stat_bpd_mispredicted,
  output [2:0]  io_com_uops_1_fetch_pc_lob,
  output [19:0] io_com_uops_1_imm_packed,
  output [11:0] io_com_uops_1_csr_addr,
  output [5:0]  io_com_uops_1_rob_idx,
  output [3:0]  io_com_uops_1_ldq_idx,
  output [3:0]  io_com_uops_1_stq_idx,
  output [4:0]  io_com_uops_1_brob_idx,
  output [6:0]  io_com_uops_1_pdst,
  output [6:0]  io_com_uops_1_pop1,
  output [6:0]  io_com_uops_1_pop2,
  output [6:0]  io_com_uops_1_pop3,
  output        io_com_uops_1_prs1_busy,
  output        io_com_uops_1_prs2_busy,
  output        io_com_uops_1_prs3_busy,
  output [6:0]  io_com_uops_1_stale_pdst,
  output        io_com_uops_1_exception,
  output [63:0] io_com_uops_1_exc_cause,
  output        io_com_uops_1_bypassable,
  output [3:0]  io_com_uops_1_mem_cmd,
  output [2:0]  io_com_uops_1_mem_typ,
  output        io_com_uops_1_is_fence,
  output        io_com_uops_1_is_fencei,
  output        io_com_uops_1_is_store,
  output        io_com_uops_1_is_amo,
  output        io_com_uops_1_is_load,
  output        io_com_uops_1_is_unique,
  output        io_com_uops_1_flush_on_commit,
  output [5:0]  io_com_uops_1_ldst,
  output [5:0]  io_com_uops_1_lrs1,
  output [5:0]  io_com_uops_1_lrs2,
  output [5:0]  io_com_uops_1_lrs3,
  output        io_com_uops_1_ldst_val,
  output [1:0]  io_com_uops_1_dst_rtype,
  output [1:0]  io_com_uops_1_lrs1_rtype,
  output [1:0]  io_com_uops_1_lrs2_rtype,
  output        io_com_uops_1_frs3_en,
  output        io_com_uops_1_fp_val,
  output        io_com_uops_1_fp_single,
  output        io_com_uops_1_xcpt_if,
  output        io_com_uops_1_replay_if,
  output [63:0] io_com_uops_1_debug_wdata,
  output [31:0] io_com_uops_1_debug_events_fetch_seq,
  output        io_com_fflags_val,
  output [4:0]  io_com_fflags,
  output        io_com_st_mask_0,
  output        io_com_st_mask_1,
  output        io_com_ld_mask_0,
  output        io_com_ld_mask_1,
  input         io_lsu_clr_bsy_valid,
  input  [5:0]  io_lsu_clr_bsy_rob_idx,
  output        io_com_load_is_at_rob_head,
  output        io_com_exception,
  output [63:0] io_com_exc_cause,
  output        io_com_handling_exc,
  output        io_com_rbk_valids_0,
  output        io_com_rbk_valids_1,
  output [63:0] io_com_badvaddr,
  input         io_brinfo_valid,
  input         io_brinfo_mispredict,
  input  [7:0]  io_brinfo_mask,
  input  [2:0]  io_brinfo_tag,
  input  [7:0]  io_brinfo_exe_mask,
  input  [5:0]  io_brinfo_rob_idx,
  input  [3:0]  io_brinfo_ldq_idx,
  input  [3:0]  io_brinfo_stq_idx,
  input         io_brinfo_taken,
  input         io_brinfo_is_jr,
  input         io_brinfo_btb_made_pred,
  input         io_brinfo_btb_mispredict,
  input         io_brinfo_bpd_made_pred,
  input         io_brinfo_bpd_mispredict,
  input  [5:0]  io_get_pc_rob_idx,
  output [39:0] io_get_pc_curr_pc,
  output [4:0]  io_get_pc_curr_brob_idx,
  output        io_get_pc_next_val,
  output [39:0] io_get_pc_next_pc,
  output        io_lsu_misspec,
  output        io_flush_take_pc,
  output [39:0] io_flush_pc,
  output        io_flush_pipeline,
  output        io_flush_brob,
  output        io_empty,
  output        io_ready,
  output        io_brob_deallocate_valid,
  output [4:0]  io_brob_deallocate_bits_brob_idx,
  output [1:0]  io_debug_state,
  output [5:0]  io_debug_rob_head,
  output        io_debug_xcpt_val,
  output        io_debug_xcpt_uop_valid,
  output [1:0]  io_debug_xcpt_uop_iw_state,
  output [8:0]  io_debug_xcpt_uop_uopc,
  output [31:0] io_debug_xcpt_uop_inst,
  output [39:0] io_debug_xcpt_uop_pc,
  output [7:0]  io_debug_xcpt_uop_fu_code,
  output [3:0]  io_debug_xcpt_uop_ctrl_br_type,
  output [1:0]  io_debug_xcpt_uop_ctrl_op1_sel,
  output [2:0]  io_debug_xcpt_uop_ctrl_op2_sel,
  output [2:0]  io_debug_xcpt_uop_ctrl_imm_sel,
  output [3:0]  io_debug_xcpt_uop_ctrl_op_fcn,
  output        io_debug_xcpt_uop_ctrl_fcn_dw,
  output        io_debug_xcpt_uop_ctrl_rf_wen,
  output [2:0]  io_debug_xcpt_uop_ctrl_csr_cmd,
  output        io_debug_xcpt_uop_ctrl_is_load,
  output        io_debug_xcpt_uop_ctrl_is_sta,
  output        io_debug_xcpt_uop_ctrl_is_std,
  output [1:0]  io_debug_xcpt_uop_wakeup_delay,
  output        io_debug_xcpt_uop_allocate_brtag,
  output        io_debug_xcpt_uop_is_br_or_jmp,
  output        io_debug_xcpt_uop_is_jump,
  output        io_debug_xcpt_uop_is_jal,
  output        io_debug_xcpt_uop_is_ret,
  output        io_debug_xcpt_uop_is_call,
  output [7:0]  io_debug_xcpt_uop_br_mask,
  output [2:0]  io_debug_xcpt_uop_br_tag,
  output        io_debug_xcpt_uop_br_prediction_bpd_predict_val,
  output        io_debug_xcpt_uop_br_prediction_bpd_predict_taken,
  output        io_debug_xcpt_uop_br_prediction_btb_hit,
  output        io_debug_xcpt_uop_br_prediction_btb_predicted,
  output        io_debug_xcpt_uop_br_prediction_is_br_or_jalr,
  output        io_debug_xcpt_uop_stat_brjmp_mispredicted,
  output        io_debug_xcpt_uop_stat_btb_made_pred,
  output        io_debug_xcpt_uop_stat_btb_mispredicted,
  output        io_debug_xcpt_uop_stat_bpd_made_pred,
  output        io_debug_xcpt_uop_stat_bpd_mispredicted,
  output [2:0]  io_debug_xcpt_uop_fetch_pc_lob,
  output [19:0] io_debug_xcpt_uop_imm_packed,
  output [11:0] io_debug_xcpt_uop_csr_addr,
  output [5:0]  io_debug_xcpt_uop_rob_idx,
  output [3:0]  io_debug_xcpt_uop_ldq_idx,
  output [3:0]  io_debug_xcpt_uop_stq_idx,
  output [4:0]  io_debug_xcpt_uop_brob_idx,
  output [6:0]  io_debug_xcpt_uop_pdst,
  output [6:0]  io_debug_xcpt_uop_pop1,
  output [6:0]  io_debug_xcpt_uop_pop2,
  output [6:0]  io_debug_xcpt_uop_pop3,
  output        io_debug_xcpt_uop_prs1_busy,
  output        io_debug_xcpt_uop_prs2_busy,
  output        io_debug_xcpt_uop_prs3_busy,
  output [6:0]  io_debug_xcpt_uop_stale_pdst,
  output        io_debug_xcpt_uop_exception,
  output [63:0] io_debug_xcpt_uop_exc_cause,
  output        io_debug_xcpt_uop_bypassable,
  output [3:0]  io_debug_xcpt_uop_mem_cmd,
  output [2:0]  io_debug_xcpt_uop_mem_typ,
  output        io_debug_xcpt_uop_is_fence,
  output        io_debug_xcpt_uop_is_fencei,
  output        io_debug_xcpt_uop_is_store,
  output        io_debug_xcpt_uop_is_amo,
  output        io_debug_xcpt_uop_is_load,
  output        io_debug_xcpt_uop_is_unique,
  output        io_debug_xcpt_uop_flush_on_commit,
  output [5:0]  io_debug_xcpt_uop_ldst,
  output [5:0]  io_debug_xcpt_uop_lrs1,
  output [5:0]  io_debug_xcpt_uop_lrs2,
  output [5:0]  io_debug_xcpt_uop_lrs3,
  output        io_debug_xcpt_uop_ldst_val,
  output [1:0]  io_debug_xcpt_uop_dst_rtype,
  output [1:0]  io_debug_xcpt_uop_lrs1_rtype,
  output [1:0]  io_debug_xcpt_uop_lrs2_rtype,
  output        io_debug_xcpt_uop_frs3_en,
  output        io_debug_xcpt_uop_fp_val,
  output        io_debug_xcpt_uop_fp_single,
  output        io_debug_xcpt_uop_xcpt_if,
  output        io_debug_xcpt_uop_replay_if,
  output [63:0] io_debug_xcpt_uop_debug_wdata,
  output [31:0] io_debug_xcpt_uop_debug_events_fetch_seq,
  output [63:0] io_debug_xcpt_badvaddr,
  input  [63:0] io_debug_tsc
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_262;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_261;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [63:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [63:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [63:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [63:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [63:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [63:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [63:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [63:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [63:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [63:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [63:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [63:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [63:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [63:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [63:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [63:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [63:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [63:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [63:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [63:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [63:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [63:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [63:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [63:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [63:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [63:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [63:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [63:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [63:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [63:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [63:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [63:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [63:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [63:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [63:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [63:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [63:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [63:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [63:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [63:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [63:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [63:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [63:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [63:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [63:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [63:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [63:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [63:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [63:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [63:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [63:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [63:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [63:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [63:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [63:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [63:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [63:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [63:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [63:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [63:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [63:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [63:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [63:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [63:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [63:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [63:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [63:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [63:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [63:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [63:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [63:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [63:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [63:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [63:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [63:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [63:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [63:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [63:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [63:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [63:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [63:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [63:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [63:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [63:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [63:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [63:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [63:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [63:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [63:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [63:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [63:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [63:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [63:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [63:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [63:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [63:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [63:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [31:0] _RAND_2862;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [63:0] _RAND_2865;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [63:0] _RAND_2889;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [63:0] _RAND_2895;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2905;
  reg [31:0] _RAND_2906;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [63:0] _RAND_2943;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2958;
  reg [31:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [63:0] _RAND_2967;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [63:0] _RAND_2973;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [31:0] _RAND_3003;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [63:0] _RAND_3021;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [63:0] _RAND_3045;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [63:0] _RAND_3051;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3055;
  reg [31:0] _RAND_3056;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3069;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [63:0] _RAND_3099;
  reg [31:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [63:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [63:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
  reg [31:0] _RAND_3140;
  reg [31:0] _RAND_3141;
  reg [31:0] _RAND_3142;
  reg [31:0] _RAND_3143;
  reg [31:0] _RAND_3144;
  reg [31:0] _RAND_3145;
  reg [31:0] _RAND_3146;
  reg [31:0] _RAND_3147;
  reg [31:0] _RAND_3148;
  reg [31:0] _RAND_3149;
  reg [31:0] _RAND_3150;
  reg [31:0] _RAND_3151;
  reg [31:0] _RAND_3152;
  reg [31:0] _RAND_3153;
  reg [31:0] _RAND_3154;
  reg [31:0] _RAND_3155;
  reg [31:0] _RAND_3156;
  reg [31:0] _RAND_3157;
  reg [31:0] _RAND_3158;
  reg [31:0] _RAND_3159;
  reg [31:0] _RAND_3160;
  reg [31:0] _RAND_3161;
  reg [31:0] _RAND_3162;
  reg [31:0] _RAND_3163;
  reg [31:0] _RAND_3164;
  reg [31:0] _RAND_3165;
  reg [31:0] _RAND_3166;
  reg [31:0] _RAND_3167;
  reg [31:0] _RAND_3168;
  reg [31:0] _RAND_3169;
  reg [31:0] _RAND_3170;
  reg [31:0] _RAND_3171;
  reg [31:0] _RAND_3172;
  reg [31:0] _RAND_3173;
  reg [31:0] _RAND_3174;
  reg [31:0] _RAND_3175;
  reg [31:0] _RAND_3176;
  reg [63:0] _RAND_3177;
  reg [31:0] _RAND_3178;
  reg [31:0] _RAND_3179;
  reg [31:0] _RAND_3180;
  reg [31:0] _RAND_3181;
  reg [31:0] _RAND_3182;
  reg [31:0] _RAND_3183;
  reg [31:0] _RAND_3184;
  reg [31:0] _RAND_3185;
  reg [31:0] _RAND_3186;
  reg [31:0] _RAND_3187;
  reg [31:0] _RAND_3188;
  reg [31:0] _RAND_3189;
  reg [31:0] _RAND_3190;
  reg [31:0] _RAND_3191;
  reg [31:0] _RAND_3192;
  reg [31:0] _RAND_3193;
  reg [31:0] _RAND_3194;
  reg [31:0] _RAND_3195;
  reg [31:0] _RAND_3196;
  reg [31:0] _RAND_3197;
  reg [31:0] _RAND_3198;
  reg [31:0] _RAND_3199;
  reg [31:0] _RAND_3200;
  reg [63:0] _RAND_3201;
  reg [31:0] _RAND_3202;
  reg [31:0] _RAND_3203;
  reg [31:0] _RAND_3204;
  reg [31:0] _RAND_3205;
  reg [31:0] _RAND_3206;
  reg [63:0] _RAND_3207;
  reg [31:0] _RAND_3208;
  reg [31:0] _RAND_3209;
  reg [31:0] _RAND_3210;
  reg [31:0] _RAND_3211;
  reg [31:0] _RAND_3212;
  reg [31:0] _RAND_3213;
  reg [31:0] _RAND_3214;
  reg [31:0] _RAND_3215;
  reg [31:0] _RAND_3216;
  reg [31:0] _RAND_3217;
  reg [31:0] _RAND_3218;
  reg [31:0] _RAND_3219;
  reg [31:0] _RAND_3220;
  reg [31:0] _RAND_3221;
  reg [31:0] _RAND_3222;
  reg [31:0] _RAND_3223;
  reg [31:0] _RAND_3224;
  reg [31:0] _RAND_3225;
  reg [31:0] _RAND_3226;
  reg [31:0] _RAND_3227;
  reg [31:0] _RAND_3228;
  reg [31:0] _RAND_3229;
  reg [31:0] _RAND_3230;
  reg [31:0] _RAND_3231;
  reg [31:0] _RAND_3232;
  reg [31:0] _RAND_3233;
  reg [31:0] _RAND_3234;
  reg [31:0] _RAND_3235;
  reg [31:0] _RAND_3236;
  reg [31:0] _RAND_3237;
  reg [31:0] _RAND_3238;
  reg [31:0] _RAND_3239;
  reg [31:0] _RAND_3240;
  reg [31:0] _RAND_3241;
  reg [31:0] _RAND_3242;
  reg [31:0] _RAND_3243;
  reg [31:0] _RAND_3244;
  reg [31:0] _RAND_3245;
  reg [31:0] _RAND_3246;
  reg [31:0] _RAND_3247;
  reg [31:0] _RAND_3248;
  reg [31:0] _RAND_3249;
  reg [31:0] _RAND_3250;
  reg [31:0] _RAND_3251;
  reg [31:0] _RAND_3252;
  reg [31:0] _RAND_3253;
  reg [31:0] _RAND_3254;
  reg [63:0] _RAND_3255;
  reg [31:0] _RAND_3256;
  reg [31:0] _RAND_3257;
  reg [31:0] _RAND_3258;
  reg [31:0] _RAND_3259;
  reg [31:0] _RAND_3260;
  reg [31:0] _RAND_3261;
  reg [31:0] _RAND_3262;
  reg [31:0] _RAND_3263;
  reg [31:0] _RAND_3264;
  reg [31:0] _RAND_3265;
  reg [31:0] _RAND_3266;
  reg [31:0] _RAND_3267;
  reg [31:0] _RAND_3268;
  reg [31:0] _RAND_3269;
  reg [31:0] _RAND_3270;
  reg [31:0] _RAND_3271;
  reg [31:0] _RAND_3272;
  reg [31:0] _RAND_3273;
  reg [31:0] _RAND_3274;
  reg [31:0] _RAND_3275;
  reg [31:0] _RAND_3276;
  reg [31:0] _RAND_3277;
  reg [31:0] _RAND_3278;
  reg [63:0] _RAND_3279;
  reg [31:0] _RAND_3280;
  reg [31:0] _RAND_3281;
  reg [31:0] _RAND_3282;
  reg [31:0] _RAND_3283;
  reg [31:0] _RAND_3284;
  reg [63:0] _RAND_3285;
  reg [31:0] _RAND_3286;
  reg [31:0] _RAND_3287;
  reg [31:0] _RAND_3288;
  reg [31:0] _RAND_3289;
  reg [31:0] _RAND_3290;
  reg [31:0] _RAND_3291;
  reg [31:0] _RAND_3292;
  reg [31:0] _RAND_3293;
  reg [31:0] _RAND_3294;
  reg [31:0] _RAND_3295;
  reg [31:0] _RAND_3296;
  reg [31:0] _RAND_3297;
  reg [31:0] _RAND_3298;
  reg [31:0] _RAND_3299;
  reg [31:0] _RAND_3300;
  reg [31:0] _RAND_3301;
  reg [31:0] _RAND_3302;
  reg [31:0] _RAND_3303;
  reg [31:0] _RAND_3304;
  reg [31:0] _RAND_3305;
  reg [31:0] _RAND_3306;
  reg [31:0] _RAND_3307;
  reg [31:0] _RAND_3308;
  reg [31:0] _RAND_3309;
  reg [31:0] _RAND_3310;
  reg [31:0] _RAND_3311;
  reg [31:0] _RAND_3312;
  reg [31:0] _RAND_3313;
  reg [31:0] _RAND_3314;
  reg [31:0] _RAND_3315;
  reg [31:0] _RAND_3316;
  reg [31:0] _RAND_3317;
  reg [31:0] _RAND_3318;
  reg [31:0] _RAND_3319;
  reg [31:0] _RAND_3320;
  reg [31:0] _RAND_3321;
  reg [31:0] _RAND_3322;
  reg [31:0] _RAND_3323;
  reg [31:0] _RAND_3324;
  reg [31:0] _RAND_3325;
  reg [31:0] _RAND_3326;
  reg [31:0] _RAND_3327;
  reg [31:0] _RAND_3328;
  reg [31:0] _RAND_3329;
  reg [31:0] _RAND_3330;
  reg [31:0] _RAND_3331;
  reg [31:0] _RAND_3332;
  reg [63:0] _RAND_3333;
  reg [31:0] _RAND_3334;
  reg [31:0] _RAND_3335;
  reg [31:0] _RAND_3336;
  reg [31:0] _RAND_3337;
  reg [31:0] _RAND_3338;
  reg [31:0] _RAND_3339;
  reg [31:0] _RAND_3340;
  reg [31:0] _RAND_3341;
  reg [31:0] _RAND_3342;
  reg [31:0] _RAND_3343;
  reg [31:0] _RAND_3344;
  reg [31:0] _RAND_3345;
  reg [31:0] _RAND_3346;
  reg [31:0] _RAND_3347;
  reg [31:0] _RAND_3348;
  reg [31:0] _RAND_3349;
  reg [31:0] _RAND_3350;
  reg [31:0] _RAND_3351;
  reg [31:0] _RAND_3352;
  reg [31:0] _RAND_3353;
  reg [31:0] _RAND_3354;
  reg [31:0] _RAND_3355;
  reg [31:0] _RAND_3356;
  reg [63:0] _RAND_3357;
  reg [31:0] _RAND_3358;
  reg [31:0] _RAND_3359;
  reg [31:0] _RAND_3360;
  reg [31:0] _RAND_3361;
  reg [31:0] _RAND_3362;
  reg [63:0] _RAND_3363;
  reg [31:0] _RAND_3364;
  reg [31:0] _RAND_3365;
  reg [31:0] _RAND_3366;
  reg [31:0] _RAND_3367;
  reg [31:0] _RAND_3368;
  reg [31:0] _RAND_3369;
  reg [31:0] _RAND_3370;
  reg [31:0] _RAND_3371;
  reg [31:0] _RAND_3372;
  reg [31:0] _RAND_3373;
  reg [31:0] _RAND_3374;
  reg [31:0] _RAND_3375;
  reg [31:0] _RAND_3376;
  reg [31:0] _RAND_3377;
  reg [31:0] _RAND_3378;
  reg [31:0] _RAND_3379;
  reg [31:0] _RAND_3380;
  reg [31:0] _RAND_3381;
  reg [31:0] _RAND_3382;
  reg [31:0] _RAND_3383;
  reg [31:0] _RAND_3384;
  reg [31:0] _RAND_3385;
  reg [31:0] _RAND_3386;
  reg [31:0] _RAND_3387;
  reg [31:0] _RAND_3388;
  reg [31:0] _RAND_3389;
  reg [31:0] _RAND_3390;
  reg [31:0] _RAND_3391;
  reg [31:0] _RAND_3392;
  reg [31:0] _RAND_3393;
  reg [31:0] _RAND_3394;
  reg [31:0] _RAND_3395;
  reg [31:0] _RAND_3396;
  reg [31:0] _RAND_3397;
  reg [31:0] _RAND_3398;
  reg [31:0] _RAND_3399;
  reg [31:0] _RAND_3400;
  reg [31:0] _RAND_3401;
  reg [31:0] _RAND_3402;
  reg [31:0] _RAND_3403;
  reg [31:0] _RAND_3404;
  reg [31:0] _RAND_3405;
  reg [31:0] _RAND_3406;
  reg [31:0] _RAND_3407;
  reg [31:0] _RAND_3408;
  reg [31:0] _RAND_3409;
  reg [31:0] _RAND_3410;
  reg [63:0] _RAND_3411;
  reg [31:0] _RAND_3412;
  reg [31:0] _RAND_3413;
  reg [31:0] _RAND_3414;
  reg [31:0] _RAND_3415;
  reg [31:0] _RAND_3416;
  reg [31:0] _RAND_3417;
  reg [31:0] _RAND_3418;
  reg [31:0] _RAND_3419;
  reg [31:0] _RAND_3420;
  reg [31:0] _RAND_3421;
  reg [31:0] _RAND_3422;
  reg [31:0] _RAND_3423;
  reg [31:0] _RAND_3424;
  reg [31:0] _RAND_3425;
  reg [31:0] _RAND_3426;
  reg [31:0] _RAND_3427;
  reg [31:0] _RAND_3428;
  reg [31:0] _RAND_3429;
  reg [31:0] _RAND_3430;
  reg [31:0] _RAND_3431;
  reg [31:0] _RAND_3432;
  reg [31:0] _RAND_3433;
  reg [31:0] _RAND_3434;
  reg [63:0] _RAND_3435;
  reg [31:0] _RAND_3436;
  reg [31:0] _RAND_3437;
  reg [31:0] _RAND_3438;
  reg [31:0] _RAND_3439;
  reg [31:0] _RAND_3440;
  reg [63:0] _RAND_3441;
  reg [31:0] _RAND_3442;
  reg [31:0] _RAND_3443;
  reg [31:0] _RAND_3444;
  reg [31:0] _RAND_3445;
  reg [31:0] _RAND_3446;
  reg [31:0] _RAND_3447;
  reg [31:0] _RAND_3448;
  reg [31:0] _RAND_3449;
  reg [31:0] _RAND_3450;
  reg [31:0] _RAND_3451;
  reg [31:0] _RAND_3452;
  reg [31:0] _RAND_3453;
  reg [31:0] _RAND_3454;
  reg [31:0] _RAND_3455;
  reg [31:0] _RAND_3456;
  reg [31:0] _RAND_3457;
  reg [31:0] _RAND_3458;
  reg [31:0] _RAND_3459;
  reg [31:0] _RAND_3460;
  reg [31:0] _RAND_3461;
  reg [31:0] _RAND_3462;
  reg [31:0] _RAND_3463;
  reg [31:0] _RAND_3464;
  reg [31:0] _RAND_3465;
  reg [31:0] _RAND_3466;
  reg [31:0] _RAND_3467;
  reg [31:0] _RAND_3468;
  reg [31:0] _RAND_3469;
  reg [31:0] _RAND_3470;
  reg [31:0] _RAND_3471;
  reg [31:0] _RAND_3472;
  reg [31:0] _RAND_3473;
  reg [31:0] _RAND_3474;
  reg [31:0] _RAND_3475;
  reg [31:0] _RAND_3476;
  reg [31:0] _RAND_3477;
  reg [31:0] _RAND_3478;
  reg [31:0] _RAND_3479;
  reg [31:0] _RAND_3480;
  reg [31:0] _RAND_3481;
  reg [31:0] _RAND_3482;
  reg [31:0] _RAND_3483;
  reg [31:0] _RAND_3484;
  reg [31:0] _RAND_3485;
  reg [31:0] _RAND_3486;
  reg [31:0] _RAND_3487;
  reg [31:0] _RAND_3488;
  reg [63:0] _RAND_3489;
  reg [31:0] _RAND_3490;
  reg [31:0] _RAND_3491;
  reg [31:0] _RAND_3492;
  reg [31:0] _RAND_3493;
  reg [31:0] _RAND_3494;
  reg [31:0] _RAND_3495;
  reg [31:0] _RAND_3496;
  reg [31:0] _RAND_3497;
  reg [31:0] _RAND_3498;
  reg [31:0] _RAND_3499;
  reg [31:0] _RAND_3500;
  reg [31:0] _RAND_3501;
  reg [31:0] _RAND_3502;
  reg [31:0] _RAND_3503;
  reg [31:0] _RAND_3504;
  reg [31:0] _RAND_3505;
  reg [31:0] _RAND_3506;
  reg [31:0] _RAND_3507;
  reg [31:0] _RAND_3508;
  reg [31:0] _RAND_3509;
  reg [31:0] _RAND_3510;
  reg [31:0] _RAND_3511;
  reg [31:0] _RAND_3512;
  reg [63:0] _RAND_3513;
  reg [31:0] _RAND_3514;
  reg [31:0] _RAND_3515;
  reg [31:0] _RAND_3516;
  reg [31:0] _RAND_3517;
  reg [31:0] _RAND_3518;
  reg [63:0] _RAND_3519;
  reg [31:0] _RAND_3520;
  reg [31:0] _RAND_3521;
  reg [31:0] _RAND_3522;
  reg [31:0] _RAND_3523;
  reg [31:0] _RAND_3524;
  reg [31:0] _RAND_3525;
  reg [31:0] _RAND_3526;
  reg [31:0] _RAND_3527;
  reg [31:0] _RAND_3528;
  reg [31:0] _RAND_3529;
  reg [31:0] _RAND_3530;
  reg [31:0] _RAND_3531;
  reg [31:0] _RAND_3532;
  reg [31:0] _RAND_3533;
  reg [31:0] _RAND_3534;
  reg [31:0] _RAND_3535;
  reg [31:0] _RAND_3536;
  reg [31:0] _RAND_3537;
  reg [31:0] _RAND_3538;
  reg [31:0] _RAND_3539;
  reg [31:0] _RAND_3540;
  reg [31:0] _RAND_3541;
  reg [31:0] _RAND_3542;
  reg [31:0] _RAND_3543;
  reg [31:0] _RAND_3544;
  reg [31:0] _RAND_3545;
  reg [31:0] _RAND_3546;
  reg [31:0] _RAND_3547;
  reg [31:0] _RAND_3548;
  reg [31:0] _RAND_3549;
  reg [31:0] _RAND_3550;
  reg [31:0] _RAND_3551;
  reg [31:0] _RAND_3552;
  reg [31:0] _RAND_3553;
  reg [31:0] _RAND_3554;
  reg [31:0] _RAND_3555;
  reg [31:0] _RAND_3556;
  reg [31:0] _RAND_3557;
  reg [31:0] _RAND_3558;
  reg [31:0] _RAND_3559;
  reg [31:0] _RAND_3560;
  reg [31:0] _RAND_3561;
  reg [31:0] _RAND_3562;
  reg [31:0] _RAND_3563;
  reg [31:0] _RAND_3564;
  reg [31:0] _RAND_3565;
  reg [31:0] _RAND_3566;
  reg [63:0] _RAND_3567;
  reg [31:0] _RAND_3568;
  reg [31:0] _RAND_3569;
  reg [31:0] _RAND_3570;
  reg [31:0] _RAND_3571;
  reg [31:0] _RAND_3572;
  reg [31:0] _RAND_3573;
  reg [31:0] _RAND_3574;
  reg [31:0] _RAND_3575;
  reg [31:0] _RAND_3576;
  reg [31:0] _RAND_3577;
  reg [31:0] _RAND_3578;
  reg [31:0] _RAND_3579;
  reg [31:0] _RAND_3580;
  reg [31:0] _RAND_3581;
  reg [31:0] _RAND_3582;
  reg [31:0] _RAND_3583;
  reg [31:0] _RAND_3584;
  reg [31:0] _RAND_3585;
  reg [31:0] _RAND_3586;
  reg [31:0] _RAND_3587;
  reg [31:0] _RAND_3588;
  reg [31:0] _RAND_3589;
  reg [31:0] _RAND_3590;
  reg [63:0] _RAND_3591;
  reg [31:0] _RAND_3592;
  reg [31:0] _RAND_3593;
  reg [31:0] _RAND_3594;
  reg [31:0] _RAND_3595;
  reg [31:0] _RAND_3596;
  reg [63:0] _RAND_3597;
  reg [31:0] _RAND_3598;
  reg [31:0] _RAND_3599;
  reg [31:0] _RAND_3600;
  reg [31:0] _RAND_3601;
  reg [31:0] _RAND_3602;
  reg [31:0] _RAND_3603;
  reg [31:0] _RAND_3604;
  reg [31:0] _RAND_3605;
  reg [31:0] _RAND_3606;
  reg [31:0] _RAND_3607;
  reg [31:0] _RAND_3608;
  reg [31:0] _RAND_3609;
  reg [31:0] _RAND_3610;
  reg [31:0] _RAND_3611;
  reg [31:0] _RAND_3612;
  reg [31:0] _RAND_3613;
  reg [31:0] _RAND_3614;
  reg [31:0] _RAND_3615;
  reg [31:0] _RAND_3616;
  reg [31:0] _RAND_3617;
  reg [31:0] _RAND_3618;
  reg [31:0] _RAND_3619;
  reg [31:0] _RAND_3620;
  reg [31:0] _RAND_3621;
  reg [31:0] _RAND_3622;
  reg [31:0] _RAND_3623;
  reg [31:0] _RAND_3624;
  reg [31:0] _RAND_3625;
  reg [31:0] _RAND_3626;
  reg [31:0] _RAND_3627;
  reg [31:0] _RAND_3628;
  reg [31:0] _RAND_3629;
  reg [31:0] _RAND_3630;
  reg [31:0] _RAND_3631;
  reg [31:0] _RAND_3632;
  reg [31:0] _RAND_3633;
  reg [31:0] _RAND_3634;
  reg [31:0] _RAND_3635;
  reg [31:0] _RAND_3636;
  reg [31:0] _RAND_3637;
  reg [31:0] _RAND_3638;
  reg [31:0] _RAND_3639;
  reg [31:0] _RAND_3640;
  reg [31:0] _RAND_3641;
  reg [31:0] _RAND_3642;
  reg [31:0] _RAND_3643;
  reg [31:0] _RAND_3644;
  reg [63:0] _RAND_3645;
  reg [31:0] _RAND_3646;
  reg [31:0] _RAND_3647;
  reg [31:0] _RAND_3648;
  reg [31:0] _RAND_3649;
  reg [31:0] _RAND_3650;
  reg [31:0] _RAND_3651;
  reg [31:0] _RAND_3652;
  reg [31:0] _RAND_3653;
  reg [31:0] _RAND_3654;
  reg [31:0] _RAND_3655;
  reg [31:0] _RAND_3656;
  reg [31:0] _RAND_3657;
  reg [31:0] _RAND_3658;
  reg [31:0] _RAND_3659;
  reg [31:0] _RAND_3660;
  reg [31:0] _RAND_3661;
  reg [31:0] _RAND_3662;
  reg [31:0] _RAND_3663;
  reg [31:0] _RAND_3664;
  reg [31:0] _RAND_3665;
  reg [31:0] _RAND_3666;
  reg [31:0] _RAND_3667;
  reg [31:0] _RAND_3668;
  reg [63:0] _RAND_3669;
  reg [31:0] _RAND_3670;
  reg [31:0] _RAND_3671;
  reg [31:0] _RAND_3672;
  reg [31:0] _RAND_3673;
  reg [31:0] _RAND_3674;
  reg [63:0] _RAND_3675;
  reg [31:0] _RAND_3676;
  reg [31:0] _RAND_3677;
  reg [31:0] _RAND_3678;
  reg [31:0] _RAND_3679;
  reg [31:0] _RAND_3680;
  reg [31:0] _RAND_3681;
  reg [31:0] _RAND_3682;
  reg [31:0] _RAND_3683;
  reg [31:0] _RAND_3684;
  reg [31:0] _RAND_3685;
  reg [31:0] _RAND_3686;
  reg [31:0] _RAND_3687;
  reg [31:0] _RAND_3688;
  reg [31:0] _RAND_3689;
  reg [31:0] _RAND_3690;
  reg [31:0] _RAND_3691;
  reg [31:0] _RAND_3692;
  reg [31:0] _RAND_3693;
  reg [31:0] _RAND_3694;
  reg [31:0] _RAND_3695;
  reg [31:0] _RAND_3696;
  reg [31:0] _RAND_3697;
  reg [31:0] _RAND_3698;
  reg [31:0] _RAND_3699;
  reg [31:0] _RAND_3700;
  reg [31:0] _RAND_3701;
  reg [31:0] _RAND_3702;
  reg [31:0] _RAND_3703;
  reg [31:0] _RAND_3704;
  reg [31:0] _RAND_3705;
  reg [31:0] _RAND_3706;
  reg [31:0] _RAND_3707;
  reg [31:0] _RAND_3708;
  reg [31:0] _RAND_3709;
  reg [31:0] _RAND_3710;
  reg [31:0] _RAND_3711;
  reg [31:0] _RAND_3712;
  reg [31:0] _RAND_3713;
  reg [31:0] _RAND_3714;
  reg [31:0] _RAND_3715;
  reg [31:0] _RAND_3716;
  reg [31:0] _RAND_3717;
  reg [31:0] _RAND_3718;
  reg [31:0] _RAND_3719;
  reg [31:0] _RAND_3720;
  reg [31:0] _RAND_3721;
  reg [31:0] _RAND_3722;
  reg [63:0] _RAND_3723;
  reg [31:0] _RAND_3724;
  reg [31:0] _RAND_3725;
  reg [31:0] _RAND_3726;
  reg [31:0] _RAND_3727;
  reg [31:0] _RAND_3728;
  reg [31:0] _RAND_3729;
  reg [31:0] _RAND_3730;
  reg [31:0] _RAND_3731;
  reg [31:0] _RAND_3732;
  reg [31:0] _RAND_3733;
  reg [31:0] _RAND_3734;
  reg [31:0] _RAND_3735;
  reg [31:0] _RAND_3736;
  reg [31:0] _RAND_3737;
  reg [31:0] _RAND_3738;
  reg [31:0] _RAND_3739;
  reg [31:0] _RAND_3740;
  reg [31:0] _RAND_3741;
  reg [31:0] _RAND_3742;
  reg [31:0] _RAND_3743;
  reg [31:0] _RAND_3744;
  reg [31:0] _RAND_3745;
  reg [31:0] _RAND_3746;
  reg [63:0] _RAND_3747;
  reg [31:0] _RAND_3748;
  reg [31:0] _RAND_3749;
  reg [31:0] _RAND_3750;
  reg [31:0] _RAND_3751;
  reg [31:0] _RAND_3752;
  reg [63:0] _RAND_3753;
  reg [31:0] _RAND_3754;
  reg [31:0] _RAND_3755;
  reg [31:0] _RAND_3756;
  reg [31:0] _RAND_3757;
  reg [31:0] _RAND_3758;
  reg [31:0] _RAND_3759;
  reg [31:0] _RAND_3760;
  reg [31:0] _RAND_3761;
  reg [31:0] _RAND_3762;
  reg [31:0] _RAND_3763;
  reg [31:0] _RAND_3764;
  reg [31:0] _RAND_3765;
  reg [31:0] _RAND_3766;
  reg [31:0] _RAND_3767;
  reg [31:0] _RAND_3768;
  reg [31:0] _RAND_3769;
  reg [31:0] _RAND_3770;
  reg [31:0] _RAND_3771;
  reg [31:0] _RAND_3772;
  reg [31:0] _RAND_3773;
  reg [31:0] _RAND_3774;
  reg [31:0] _RAND_3775;
  reg [31:0] _RAND_3776;
  reg [31:0] _RAND_3777;
  reg [31:0] _RAND_3778;
  reg [31:0] _RAND_3779;
  reg [31:0] _RAND_3780;
  reg [31:0] _RAND_3781;
  reg [31:0] _RAND_3782;
  reg [31:0] _RAND_3783;
  reg [31:0] _RAND_3784;
  reg [31:0] _RAND_3785;
  reg [31:0] _RAND_3786;
  reg [31:0] _RAND_3787;
  reg [31:0] _RAND_3788;
  reg [31:0] _RAND_3789;
  reg [31:0] _RAND_3790;
  reg [31:0] _RAND_3791;
  reg [31:0] _RAND_3792;
  reg [31:0] _RAND_3793;
  reg [31:0] _RAND_3794;
  reg [31:0] _RAND_3795;
  reg [31:0] _RAND_3796;
  reg [31:0] _RAND_3797;
  reg [31:0] _RAND_3798;
  reg [31:0] _RAND_3799;
  reg [31:0] _RAND_3800;
  reg [63:0] _RAND_3801;
  reg [31:0] _RAND_3802;
  reg [31:0] _RAND_3803;
  reg [31:0] _RAND_3804;
  reg [31:0] _RAND_3805;
  reg [31:0] _RAND_3806;
  reg [31:0] _RAND_3807;
  reg [31:0] _RAND_3808;
  reg [31:0] _RAND_3809;
  reg [31:0] _RAND_3810;
  reg [31:0] _RAND_3811;
  reg [31:0] _RAND_3812;
  reg [31:0] _RAND_3813;
  reg [31:0] _RAND_3814;
  reg [31:0] _RAND_3815;
  reg [31:0] _RAND_3816;
  reg [31:0] _RAND_3817;
  reg [31:0] _RAND_3818;
  reg [31:0] _RAND_3819;
  reg [31:0] _RAND_3820;
  reg [31:0] _RAND_3821;
  reg [31:0] _RAND_3822;
  reg [31:0] _RAND_3823;
  reg [31:0] _RAND_3824;
  reg [63:0] _RAND_3825;
  reg [31:0] _RAND_3826;
  reg [31:0] _RAND_3827;
  reg [31:0] _RAND_3828;
  reg [31:0] _RAND_3829;
  reg [31:0] _RAND_3830;
  reg [63:0] _RAND_3831;
  reg [31:0] _RAND_3832;
  reg [31:0] _RAND_3833;
  reg [31:0] _RAND_3834;
  reg [31:0] _RAND_3835;
  reg [31:0] _RAND_3836;
  reg [31:0] _RAND_3837;
  reg [31:0] _RAND_3838;
  reg [31:0] _RAND_3839;
  reg [31:0] _RAND_3840;
  reg [31:0] _RAND_3841;
  reg [31:0] _RAND_3842;
  reg [31:0] _RAND_3843;
  reg [31:0] _RAND_3844;
  reg [31:0] _RAND_3845;
  reg [31:0] _RAND_3846;
  reg [31:0] _RAND_3847;
  reg [31:0] _RAND_3848;
  reg [31:0] _RAND_3849;
  reg [31:0] _RAND_3850;
  reg [31:0] _RAND_3851;
  reg [31:0] _RAND_3852;
  reg [31:0] _RAND_3853;
  reg [31:0] _RAND_3854;
  reg [31:0] _RAND_3855;
  reg [31:0] _RAND_3856;
  reg [31:0] _RAND_3857;
  reg [31:0] _RAND_3858;
  reg [31:0] _RAND_3859;
  reg [31:0] _RAND_3860;
  reg [31:0] _RAND_3861;
  reg [31:0] _RAND_3862;
  reg [31:0] _RAND_3863;
  reg [31:0] _RAND_3864;
  reg [31:0] _RAND_3865;
  reg [31:0] _RAND_3866;
  reg [31:0] _RAND_3867;
  reg [31:0] _RAND_3868;
  reg [31:0] _RAND_3869;
  reg [31:0] _RAND_3870;
  reg [31:0] _RAND_3871;
  reg [31:0] _RAND_3872;
  reg [31:0] _RAND_3873;
  reg [31:0] _RAND_3874;
  reg [31:0] _RAND_3875;
  reg [31:0] _RAND_3876;
  reg [31:0] _RAND_3877;
  reg [31:0] _RAND_3878;
  reg [63:0] _RAND_3879;
  reg [31:0] _RAND_3880;
  reg [31:0] _RAND_3881;
  reg [31:0] _RAND_3882;
  reg [31:0] _RAND_3883;
  reg [31:0] _RAND_3884;
  reg [31:0] _RAND_3885;
  reg [31:0] _RAND_3886;
  reg [31:0] _RAND_3887;
  reg [31:0] _RAND_3888;
  reg [31:0] _RAND_3889;
  reg [31:0] _RAND_3890;
  reg [31:0] _RAND_3891;
  reg [31:0] _RAND_3892;
  reg [31:0] _RAND_3893;
  reg [31:0] _RAND_3894;
  reg [31:0] _RAND_3895;
  reg [31:0] _RAND_3896;
  reg [31:0] _RAND_3897;
  reg [31:0] _RAND_3898;
  reg [31:0] _RAND_3899;
  reg [31:0] _RAND_3900;
  reg [31:0] _RAND_3901;
  reg [31:0] _RAND_3902;
  reg [63:0] _RAND_3903;
  reg [31:0] _RAND_3904;
  reg [31:0] _RAND_3905;
  reg [31:0] _RAND_3906;
  reg [31:0] _RAND_3907;
  reg [31:0] _RAND_3908;
  reg [63:0] _RAND_3909;
  reg [31:0] _RAND_3910;
  reg [31:0] _RAND_3911;
  reg [31:0] _RAND_3912;
  reg [31:0] _RAND_3913;
  reg [31:0] _RAND_3914;
  reg [31:0] _RAND_3915;
  reg [31:0] _RAND_3916;
  reg [31:0] _RAND_3917;
  reg [31:0] _RAND_3918;
  reg [31:0] _RAND_3919;
  reg [31:0] _RAND_3920;
  reg [31:0] _RAND_3921;
  reg [31:0] _RAND_3922;
  reg [31:0] _RAND_3923;
  reg [31:0] _RAND_3924;
  reg [31:0] _RAND_3925;
  reg [31:0] _RAND_3926;
  reg [31:0] _RAND_3927;
  reg [31:0] _RAND_3928;
  reg [31:0] _RAND_3929;
  reg [31:0] _RAND_3930;
  reg [31:0] _RAND_3931;
  reg [31:0] _RAND_3932;
  reg [31:0] _RAND_3933;
  reg [31:0] _RAND_3934;
  reg [31:0] _RAND_3935;
  reg [31:0] _RAND_3936;
  reg [31:0] _RAND_3937;
  reg [31:0] _RAND_3938;
  reg [31:0] _RAND_3939;
  reg [31:0] _RAND_3940;
  reg [31:0] _RAND_3941;
  reg [31:0] _RAND_3942;
  reg [31:0] _RAND_3943;
  reg [31:0] _RAND_3944;
  reg [31:0] _RAND_3945;
  reg [31:0] _RAND_3946;
  reg [31:0] _RAND_3947;
  reg [31:0] _RAND_3948;
  reg [31:0] _RAND_3949;
  reg [31:0] _RAND_3950;
  reg [31:0] _RAND_3951;
  reg [31:0] _RAND_3952;
  reg [31:0] _RAND_3953;
  reg [31:0] _RAND_3954;
  reg [31:0] _RAND_3955;
  reg [31:0] _RAND_3956;
  reg [63:0] _RAND_3957;
  reg [31:0] _RAND_3958;
  reg [31:0] _RAND_3959;
  reg [31:0] _RAND_3960;
  reg [31:0] _RAND_3961;
  reg [31:0] _RAND_3962;
  reg [31:0] _RAND_3963;
  reg [31:0] _RAND_3964;
  reg [31:0] _RAND_3965;
  reg [31:0] _RAND_3966;
  reg [31:0] _RAND_3967;
  reg [31:0] _RAND_3968;
  reg [31:0] _RAND_3969;
  reg [31:0] _RAND_3970;
  reg [31:0] _RAND_3971;
  reg [31:0] _RAND_3972;
  reg [31:0] _RAND_3973;
  reg [31:0] _RAND_3974;
  reg [31:0] _RAND_3975;
  reg [31:0] _RAND_3976;
  reg [31:0] _RAND_3977;
  reg [31:0] _RAND_3978;
  reg [31:0] _RAND_3979;
  reg [31:0] _RAND_3980;
  reg [63:0] _RAND_3981;
  reg [31:0] _RAND_3982;
  reg [31:0] _RAND_3983;
  reg [31:0] _RAND_3984;
  reg [31:0] _RAND_3985;
  reg [31:0] _RAND_3986;
  reg [63:0] _RAND_3987;
  reg [31:0] _RAND_3988;
  reg [31:0] _RAND_3989;
  reg [31:0] _RAND_3990;
  reg [31:0] _RAND_3991;
  reg [31:0] _RAND_3992;
  reg [31:0] _RAND_3993;
  reg [31:0] _RAND_3994;
  reg [31:0] _RAND_3995;
  reg [31:0] _RAND_3996;
  reg [31:0] _RAND_3997;
  reg [31:0] _RAND_3998;
  reg [31:0] _RAND_3999;
  reg [31:0] _RAND_4000;
  reg [31:0] _RAND_4001;
  reg [31:0] _RAND_4002;
  reg [31:0] _RAND_4003;
  reg [31:0] _RAND_4004;
  reg [31:0] _RAND_4005;
  reg [31:0] _RAND_4006;
  reg [31:0] _RAND_4007;
  reg [31:0] _RAND_4008;
  reg [31:0] _RAND_4009;
  reg [31:0] _RAND_4010;
  reg [31:0] _RAND_4011;
  reg [31:0] _RAND_4012;
  reg [31:0] _RAND_4013;
  reg [31:0] _RAND_4014;
  reg [31:0] _RAND_4015;
  reg [31:0] _RAND_4016;
  reg [31:0] _RAND_4017;
  reg [31:0] _RAND_4018;
  reg [31:0] _RAND_4019;
  reg [31:0] _RAND_4020;
  reg [31:0] _RAND_4021;
  reg [31:0] _RAND_4022;
  reg [31:0] _RAND_4023;
  reg [31:0] _RAND_4024;
  reg [31:0] _RAND_4025;
  reg [31:0] _RAND_4026;
  reg [31:0] _RAND_4027;
  reg [31:0] _RAND_4028;
  reg [31:0] _RAND_4029;
  reg [31:0] _RAND_4030;
  reg [31:0] _RAND_4031;
  reg [31:0] _RAND_4032;
  reg [31:0] _RAND_4033;
  reg [31:0] _RAND_4034;
  reg [63:0] _RAND_4035;
  reg [31:0] _RAND_4036;
  reg [31:0] _RAND_4037;
  reg [31:0] _RAND_4038;
  reg [31:0] _RAND_4039;
  reg [31:0] _RAND_4040;
  reg [31:0] _RAND_4041;
  reg [31:0] _RAND_4042;
  reg [31:0] _RAND_4043;
  reg [31:0] _RAND_4044;
  reg [31:0] _RAND_4045;
  reg [31:0] _RAND_4046;
  reg [31:0] _RAND_4047;
  reg [31:0] _RAND_4048;
  reg [31:0] _RAND_4049;
  reg [31:0] _RAND_4050;
  reg [31:0] _RAND_4051;
  reg [31:0] _RAND_4052;
  reg [31:0] _RAND_4053;
  reg [31:0] _RAND_4054;
  reg [31:0] _RAND_4055;
  reg [31:0] _RAND_4056;
  reg [31:0] _RAND_4057;
  reg [31:0] _RAND_4058;
  reg [63:0] _RAND_4059;
  reg [31:0] _RAND_4060;
  reg [31:0] _RAND_4061;
  reg [31:0] _RAND_4062;
  reg [31:0] _RAND_4063;
  reg [31:0] _RAND_4064;
  reg [63:0] _RAND_4065;
  reg [31:0] _RAND_4066;
  reg [31:0] _RAND_4067;
  reg [31:0] _RAND_4068;
  reg [31:0] _RAND_4069;
  reg [31:0] _RAND_4070;
  reg [31:0] _RAND_4071;
  reg [31:0] _RAND_4072;
  reg [31:0] _RAND_4073;
  reg [31:0] _RAND_4074;
  reg [31:0] _RAND_4075;
  reg [31:0] _RAND_4076;
  reg [31:0] _RAND_4077;
  reg [31:0] _RAND_4078;
  reg [31:0] _RAND_4079;
  reg [31:0] _RAND_4080;
  reg [31:0] _RAND_4081;
  reg [31:0] _RAND_4082;
  reg [31:0] _RAND_4083;
  reg [31:0] _RAND_4084;
  reg [31:0] _RAND_4085;
  reg [31:0] _RAND_4086;
  reg [31:0] _RAND_4087;
  reg [31:0] _RAND_4088;
  reg [31:0] _RAND_4089;
  reg [31:0] _RAND_4090;
  reg [31:0] _RAND_4091;
  reg [31:0] _RAND_4092;
  reg [31:0] _RAND_4093;
  reg [31:0] _RAND_4094;
  reg [31:0] _RAND_4095;
  reg [31:0] _RAND_4096;
  reg [31:0] _RAND_4097;
  reg [31:0] _RAND_4098;
  reg [31:0] _RAND_4099;
  reg [31:0] _RAND_4100;
  reg [31:0] _RAND_4101;
  reg [31:0] _RAND_4102;
  reg [31:0] _RAND_4103;
  reg [31:0] _RAND_4104;
  reg [31:0] _RAND_4105;
  reg [31:0] _RAND_4106;
  reg [31:0] _RAND_4107;
  reg [31:0] _RAND_4108;
  reg [31:0] _RAND_4109;
  reg [31:0] _RAND_4110;
  reg [31:0] _RAND_4111;
  reg [31:0] _RAND_4112;
  reg [63:0] _RAND_4113;
  reg [31:0] _RAND_4114;
  reg [31:0] _RAND_4115;
  reg [31:0] _RAND_4116;
  reg [31:0] _RAND_4117;
  reg [31:0] _RAND_4118;
  reg [31:0] _RAND_4119;
  reg [31:0] _RAND_4120;
  reg [31:0] _RAND_4121;
  reg [31:0] _RAND_4122;
  reg [31:0] _RAND_4123;
  reg [31:0] _RAND_4124;
  reg [31:0] _RAND_4125;
  reg [31:0] _RAND_4126;
  reg [31:0] _RAND_4127;
  reg [31:0] _RAND_4128;
  reg [31:0] _RAND_4129;
  reg [31:0] _RAND_4130;
  reg [31:0] _RAND_4131;
  reg [31:0] _RAND_4132;
  reg [31:0] _RAND_4133;
  reg [31:0] _RAND_4134;
  reg [31:0] _RAND_4135;
  reg [31:0] _RAND_4136;
  reg [63:0] _RAND_4137;
  reg [31:0] _RAND_4138;
  reg [31:0] _RAND_4139;
  reg [31:0] _RAND_4140;
`endif // RANDOMIZE_REG_INIT
  reg [36:0] T_23555 [0:11]; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_23587_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_23587_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_32958_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_32958_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33072_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33072_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33186_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33186_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33300_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33300_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33414_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33414_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33528_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33528_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33642_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33642_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33756_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33756_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33870_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33870_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_33984_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_33984_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34098_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34098_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34212_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34212_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34326_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34326_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34440_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34440_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34554_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34554_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34668_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34668_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34782_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34782_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_34896_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_34896_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_35010_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_35010_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_35124_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_35124_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_35238_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_35238_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_35352_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_35352_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_35466_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_35466_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_35580_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_35580_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_44886_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_44886_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45000_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45000_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45114_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45114_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45228_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45228_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45342_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45342_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45456_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45456_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45570_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45570_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45684_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45684_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45798_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45798_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_45912_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_45912_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46026_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46026_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46140_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46140_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46254_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46254_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46368_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46368_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46482_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46482_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46596_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46596_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46710_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46710_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46824_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46824_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_46938_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_46938_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_47052_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_47052_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_47166_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_47166_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_47280_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_47280_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_47394_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_47394_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_47508_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_47508_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_47587_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_47587_addr; // @[rob.scala 893:22]
  wire [36:0] T_23555_T_23571_data; // @[rob.scala 893:22]
  wire [3:0] T_23555_T_23571_addr; // @[rob.scala 893:22]
  wire  T_23555_T_23571_mask; // @[rob.scala 893:22]
  wire  T_23555_T_23571_en; // @[rob.scala 893:22]
  reg [36:0] T_23558 [0:11]; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_23592_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_23592_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_32964_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_32964_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33078_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33078_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33192_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33192_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33306_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33306_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33420_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33420_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33534_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33534_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33648_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33648_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33762_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33762_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33876_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33876_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_33990_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_33990_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34104_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34104_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34218_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34218_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34332_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34332_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34446_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34446_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34560_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34560_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34674_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34674_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34788_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34788_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_34902_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_34902_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_35016_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_35016_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_35130_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_35130_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_35244_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_35244_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_35358_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_35358_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_35472_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_35472_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_35586_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_35586_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_44892_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_44892_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45006_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45006_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45120_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45120_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45234_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45234_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45348_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45348_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45462_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45462_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45576_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45576_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45690_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45690_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45804_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45804_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_45918_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_45918_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46032_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46032_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46146_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46146_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46260_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46260_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46374_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46374_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46488_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46488_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46602_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46602_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46716_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46716_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46830_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46830_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_46944_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_46944_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_47058_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_47058_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_47172_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_47172_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_47286_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_47286_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_47400_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_47400_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_47514_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_47514_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_47593_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_47593_addr; // @[rob.scala 894:22]
  wire [36:0] T_23558_T_23566_data; // @[rob.scala 894:22]
  wire [3:0] T_23558_T_23566_addr; // @[rob.scala 894:22]
  wire  T_23558_T_23566_mask; // @[rob.scala 894:22]
  wire  T_23558_T_23566_en; // @[rob.scala 894:22]
  reg [4:0] row_metadata_brob_idx [0:23]; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_23666_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_23666_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_23669_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_23669_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48247_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48247_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48333_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48333_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48419_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48419_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48505_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48505_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48591_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48591_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48677_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48677_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48763_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48763_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48849_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48849_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48935_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_48935_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49021_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49021_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49107_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49107_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49193_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49193_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49279_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49279_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49365_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49365_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49451_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49451_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49537_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49537_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49623_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49623_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49709_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49709_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49795_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49795_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49881_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49881_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49967_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_49967_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_50053_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_50053_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_50139_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_50139_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_50225_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_50225_addr; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_23653_data; // @[rob.scala 295:35]
  wire [4:0] row_metadata_brob_idx_T_23653_addr; // @[rob.scala 295:35]
  wire  row_metadata_brob_idx_T_23653_mask; // @[rob.scala 295:35]
  wire  row_metadata_brob_idx_T_23653_en; // @[rob.scala 295:35]
  reg  row_metadata_has_brorjalr [0:23]; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23664_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_23664_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48249_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48249_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48335_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48335_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48421_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48421_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48507_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48507_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48593_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48593_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48679_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48679_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48765_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48765_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48851_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48851_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_48937_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_48937_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49023_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49023_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49109_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49109_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49195_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49195_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49281_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49281_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49367_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49367_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49453_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49453_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49539_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49539_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49625_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49625_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49711_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49711_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49797_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49797_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49883_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49883_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_49969_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_49969_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_50055_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_50055_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_50141_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_50141_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_50227_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_50227_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23654_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_23654_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23654_mask; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23654_en; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23662_data; // @[rob.scala 296:38]
  wire [4:0] row_metadata_has_brorjalr_T_23662_addr; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23662_mask; // @[rob.scala 296:38]
  wire  row_metadata_has_brorjalr_T_23662_en; // @[rob.scala 296:38]
  reg  T_23710 [0:23]; // @[rob.scala 335:30]
  wire  T_23710_T_29091_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_29091_addr; // @[rob.scala 335:30]
  wire  T_23710_T_32866_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_32866_addr; // @[rob.scala 335:30]
  wire  T_23710_T_32980_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_32980_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33094_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33094_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33208_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33208_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33322_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33322_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33436_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33436_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33550_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33550_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33664_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33664_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33778_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33778_addr; // @[rob.scala 335:30]
  wire  T_23710_T_33892_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_33892_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34006_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34006_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34120_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34120_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34234_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34234_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34348_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34348_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34462_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34462_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34576_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34576_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34690_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34690_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34804_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34804_addr; // @[rob.scala 335:30]
  wire  T_23710_T_34918_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_34918_addr; // @[rob.scala 335:30]
  wire  T_23710_T_35032_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_35032_addr; // @[rob.scala 335:30]
  wire  T_23710_T_35146_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_35146_addr; // @[rob.scala 335:30]
  wire  T_23710_T_35260_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_35260_addr; // @[rob.scala 335:30]
  wire  T_23710_T_35374_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_35374_addr; // @[rob.scala 335:30]
  wire  T_23710_T_35488_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_35488_addr; // @[rob.scala 335:30]
  wire  T_23710_T_28316_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_28316_addr; // @[rob.scala 335:30]
  wire  T_23710_T_28316_mask; // @[rob.scala 335:30]
  wire  T_23710_T_28316_en; // @[rob.scala 335:30]
  wire  T_23710_T_28594_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_28594_addr; // @[rob.scala 335:30]
  wire  T_23710_T_28594_mask; // @[rob.scala 335:30]
  wire  T_23710_T_28594_en; // @[rob.scala 335:30]
  wire  T_23710_T_28602_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_28602_addr; // @[rob.scala 335:30]
  wire  T_23710_T_28602_mask; // @[rob.scala 335:30]
  wire  T_23710_T_28602_en; // @[rob.scala 335:30]
  wire  T_23710_T_28610_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_28610_addr; // @[rob.scala 335:30]
  wire  T_23710_T_28610_mask; // @[rob.scala 335:30]
  wire  T_23710_T_28610_en; // @[rob.scala 335:30]
  wire  T_23710_T_28618_data; // @[rob.scala 335:30]
  wire [4:0] T_23710_T_28618_addr; // @[rob.scala 335:30]
  wire  T_23710_T_28618_mask; // @[rob.scala 335:30]
  wire  T_23710_T_28618_en; // @[rob.scala 335:30]
  reg  T_28311 [0:23]; // @[rob.scala 339:30]
  wire  T_28311_T_29089_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_29089_addr; // @[rob.scala 339:30]
  wire  T_28311_T_32978_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_32978_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33092_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33092_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33206_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33206_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33320_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33320_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33434_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33434_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33548_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33548_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33662_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33662_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33776_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33776_addr; // @[rob.scala 339:30]
  wire  T_28311_T_33890_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_33890_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34004_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34004_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34118_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34118_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34232_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34232_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34346_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34346_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34460_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34460_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34574_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34574_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34688_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34688_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34802_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34802_addr; // @[rob.scala 339:30]
  wire  T_28311_T_34916_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_34916_addr; // @[rob.scala 339:30]
  wire  T_28311_T_35030_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_35030_addr; // @[rob.scala 339:30]
  wire  T_28311_T_35144_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_35144_addr; // @[rob.scala 339:30]
  wire  T_28311_T_35258_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_35258_addr; // @[rob.scala 339:30]
  wire  T_28311_T_35372_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_35372_addr; // @[rob.scala 339:30]
  wire  T_28311_T_35486_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_35486_addr; // @[rob.scala 339:30]
  wire  T_28311_T_35600_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_35600_addr; // @[rob.scala 339:30]
  wire  T_28311_T_28407_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_28407_addr; // @[rob.scala 339:30]
  wire  T_28311_T_28407_mask; // @[rob.scala 339:30]
  wire  T_28311_T_28407_en; // @[rob.scala 339:30]
  wire  T_28311_T_29079_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_29079_addr; // @[rob.scala 339:30]
  wire  T_28311_T_29079_mask; // @[rob.scala 339:30]
  wire  T_28311_T_29079_en; // @[rob.scala 339:30]
  wire  T_28311_T_29087_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_29087_addr; // @[rob.scala 339:30]
  wire  T_28311_T_29087_mask; // @[rob.scala 339:30]
  wire  T_28311_T_29087_en; // @[rob.scala 339:30]
  wire  T_28311_T_29363_data; // @[rob.scala 339:30]
  wire [4:0] T_28311_T_29363_addr; // @[rob.scala 339:30]
  wire  T_28311_T_29363_mask; // @[rob.scala 339:30]
  wire  T_28311_T_29363_en; // @[rob.scala 339:30]
  reg [4:0] T_28314 [0:23]; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_31814_data; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_31814_addr; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_28408_data; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_28408_addr; // @[rob.scala 340:30]
  wire  T_28314_T_28408_mask; // @[rob.scala 340:30]
  wire  T_28314_T_28408_en; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_29065_data; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_29065_addr; // @[rob.scala 340:30]
  wire  T_28314_T_29065_mask; // @[rob.scala 340:30]
  wire  T_28314_T_29065_en; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_29072_data; // @[rob.scala 340:30]
  wire [4:0] T_28314_T_29072_addr; // @[rob.scala 340:30]
  wire  T_28314_T_29072_mask; // @[rob.scala 340:30]
  wire  T_28314_T_29072_en; // @[rob.scala 340:30]
  reg  T_35638 [0:23]; // @[rob.scala 335:30]
  wire  T_35638_T_41019_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_41019_addr; // @[rob.scala 335:30]
  wire  T_35638_T_44794_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_44794_addr; // @[rob.scala 335:30]
  wire  T_35638_T_44908_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_44908_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45022_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45022_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45136_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45136_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45250_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45250_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45364_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45364_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45478_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45478_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45592_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45592_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45706_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45706_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45820_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45820_addr; // @[rob.scala 335:30]
  wire  T_35638_T_45934_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_45934_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46048_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46048_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46162_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46162_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46276_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46276_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46390_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46390_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46504_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46504_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46618_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46618_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46732_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46732_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46846_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46846_addr; // @[rob.scala 335:30]
  wire  T_35638_T_46960_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_46960_addr; // @[rob.scala 335:30]
  wire  T_35638_T_47074_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_47074_addr; // @[rob.scala 335:30]
  wire  T_35638_T_47188_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_47188_addr; // @[rob.scala 335:30]
  wire  T_35638_T_47302_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_47302_addr; // @[rob.scala 335:30]
  wire  T_35638_T_47416_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_47416_addr; // @[rob.scala 335:30]
  wire  T_35638_T_40244_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_40244_addr; // @[rob.scala 335:30]
  wire  T_35638_T_40244_mask; // @[rob.scala 335:30]
  wire  T_35638_T_40244_en; // @[rob.scala 335:30]
  wire  T_35638_T_40522_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_40522_addr; // @[rob.scala 335:30]
  wire  T_35638_T_40522_mask; // @[rob.scala 335:30]
  wire  T_35638_T_40522_en; // @[rob.scala 335:30]
  wire  T_35638_T_40530_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_40530_addr; // @[rob.scala 335:30]
  wire  T_35638_T_40530_mask; // @[rob.scala 335:30]
  wire  T_35638_T_40530_en; // @[rob.scala 335:30]
  wire  T_35638_T_40538_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_40538_addr; // @[rob.scala 335:30]
  wire  T_35638_T_40538_mask; // @[rob.scala 335:30]
  wire  T_35638_T_40538_en; // @[rob.scala 335:30]
  wire  T_35638_T_40546_data; // @[rob.scala 335:30]
  wire [4:0] T_35638_T_40546_addr; // @[rob.scala 335:30]
  wire  T_35638_T_40546_mask; // @[rob.scala 335:30]
  wire  T_35638_T_40546_en; // @[rob.scala 335:30]
  reg  T_40239 [0:23]; // @[rob.scala 339:30]
  wire  T_40239_T_41017_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_41017_addr; // @[rob.scala 339:30]
  wire  T_40239_T_44906_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_44906_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45020_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45020_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45134_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45134_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45248_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45248_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45362_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45362_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45476_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45476_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45590_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45590_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45704_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45704_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45818_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45818_addr; // @[rob.scala 339:30]
  wire  T_40239_T_45932_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_45932_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46046_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46046_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46160_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46160_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46274_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46274_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46388_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46388_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46502_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46502_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46616_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46616_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46730_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46730_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46844_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46844_addr; // @[rob.scala 339:30]
  wire  T_40239_T_46958_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_46958_addr; // @[rob.scala 339:30]
  wire  T_40239_T_47072_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_47072_addr; // @[rob.scala 339:30]
  wire  T_40239_T_47186_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_47186_addr; // @[rob.scala 339:30]
  wire  T_40239_T_47300_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_47300_addr; // @[rob.scala 339:30]
  wire  T_40239_T_47414_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_47414_addr; // @[rob.scala 339:30]
  wire  T_40239_T_47528_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_47528_addr; // @[rob.scala 339:30]
  wire  T_40239_T_40335_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_40335_addr; // @[rob.scala 339:30]
  wire  T_40239_T_40335_mask; // @[rob.scala 339:30]
  wire  T_40239_T_40335_en; // @[rob.scala 339:30]
  wire  T_40239_T_41007_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_41007_addr; // @[rob.scala 339:30]
  wire  T_40239_T_41007_mask; // @[rob.scala 339:30]
  wire  T_40239_T_41007_en; // @[rob.scala 339:30]
  wire  T_40239_T_41015_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_41015_addr; // @[rob.scala 339:30]
  wire  T_40239_T_41015_mask; // @[rob.scala 339:30]
  wire  T_40239_T_41015_en; // @[rob.scala 339:30]
  wire  T_40239_T_41291_data; // @[rob.scala 339:30]
  wire [4:0] T_40239_T_41291_addr; // @[rob.scala 339:30]
  wire  T_40239_T_41291_mask; // @[rob.scala 339:30]
  wire  T_40239_T_41291_en; // @[rob.scala 339:30]
  reg [4:0] T_40242 [0:23]; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_43742_data; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_43742_addr; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_40336_data; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_40336_addr; // @[rob.scala 340:30]
  wire  T_40242_T_40336_mask; // @[rob.scala 340:30]
  wire  T_40242_T_40336_en; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_40993_data; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_40993_addr; // @[rob.scala 340:30]
  wire  T_40242_T_40993_mask; // @[rob.scala 340:30]
  wire  T_40242_T_40993_en; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_41000_data; // @[rob.scala 340:30]
  wire [4:0] T_40242_T_41000_addr; // @[rob.scala 340:30]
  wire  T_40242_T_41000_mask; // @[rob.scala 340:30]
  wire  T_40242_T_41000_en; // @[rob.scala 340:30]
  reg [1:0] rob_state;
  reg [4:0] rob_head;
  reg [4:0] rob_tail;
  wire [5:0] rob_tail_idx = {rob_tail, 1'h0}; // @[rob.scala 192:32]
  reg  r_xcpt_val;
  reg  r_xcpt_uop_valid;
  reg [1:0] r_xcpt_uop_iw_state;
  reg [8:0] r_xcpt_uop_uopc;
  reg [31:0] r_xcpt_uop_inst;
  reg [39:0] r_xcpt_uop_pc;
  reg [7:0] r_xcpt_uop_fu_code;
  reg [3:0] r_xcpt_uop_ctrl_br_type;
  reg [1:0] r_xcpt_uop_ctrl_op1_sel;
  reg [2:0] r_xcpt_uop_ctrl_op2_sel;
  reg [2:0] r_xcpt_uop_ctrl_imm_sel;
  reg [3:0] r_xcpt_uop_ctrl_op_fcn;
  reg  r_xcpt_uop_ctrl_fcn_dw;
  reg  r_xcpt_uop_ctrl_rf_wen;
  reg [2:0] r_xcpt_uop_ctrl_csr_cmd;
  reg  r_xcpt_uop_ctrl_is_load;
  reg  r_xcpt_uop_ctrl_is_sta;
  reg  r_xcpt_uop_ctrl_is_std;
  reg [1:0] r_xcpt_uop_wakeup_delay;
  reg  r_xcpt_uop_allocate_brtag;
  reg  r_xcpt_uop_is_br_or_jmp;
  reg  r_xcpt_uop_is_jump;
  reg  r_xcpt_uop_is_jal;
  reg  r_xcpt_uop_is_ret;
  reg  r_xcpt_uop_is_call;
  reg [7:0] r_xcpt_uop_br_mask;
  reg [2:0] r_xcpt_uop_br_tag;
  reg  r_xcpt_uop_br_prediction_bpd_predict_val;
  reg  r_xcpt_uop_br_prediction_bpd_predict_taken;
  reg  r_xcpt_uop_br_prediction_btb_hit;
  reg  r_xcpt_uop_br_prediction_btb_predicted;
  reg  r_xcpt_uop_br_prediction_is_br_or_jalr;
  reg  r_xcpt_uop_stat_brjmp_mispredicted;
  reg  r_xcpt_uop_stat_btb_made_pred;
  reg  r_xcpt_uop_stat_btb_mispredicted;
  reg  r_xcpt_uop_stat_bpd_made_pred;
  reg  r_xcpt_uop_stat_bpd_mispredicted;
  reg [2:0] r_xcpt_uop_fetch_pc_lob;
  reg [19:0] r_xcpt_uop_imm_packed;
  reg [11:0] r_xcpt_uop_csr_addr;
  reg [5:0] r_xcpt_uop_rob_idx;
  reg [3:0] r_xcpt_uop_ldq_idx;
  reg [3:0] r_xcpt_uop_stq_idx;
  reg [4:0] r_xcpt_uop_brob_idx;
  reg [6:0] r_xcpt_uop_pdst;
  reg [6:0] r_xcpt_uop_pop1;
  reg [6:0] r_xcpt_uop_pop2;
  reg [6:0] r_xcpt_uop_pop3;
  reg  r_xcpt_uop_prs1_busy;
  reg  r_xcpt_uop_prs2_busy;
  reg  r_xcpt_uop_prs3_busy;
  reg [6:0] r_xcpt_uop_stale_pdst;
  reg  r_xcpt_uop_exception;
  reg [63:0] r_xcpt_uop_exc_cause;
  reg  r_xcpt_uop_bypassable;
  reg [3:0] r_xcpt_uop_mem_cmd;
  reg [2:0] r_xcpt_uop_mem_typ;
  reg  r_xcpt_uop_is_fence;
  reg  r_xcpt_uop_is_fencei;
  reg  r_xcpt_uop_is_store;
  reg  r_xcpt_uop_is_amo;
  reg  r_xcpt_uop_is_load;
  reg  r_xcpt_uop_is_unique;
  reg  r_xcpt_uop_flush_on_commit;
  reg [5:0] r_xcpt_uop_ldst;
  reg [5:0] r_xcpt_uop_lrs1;
  reg [5:0] r_xcpt_uop_lrs2;
  reg [5:0] r_xcpt_uop_lrs3;
  reg  r_xcpt_uop_ldst_val;
  reg [1:0] r_xcpt_uop_dst_rtype;
  reg [1:0] r_xcpt_uop_lrs1_rtype;
  reg [1:0] r_xcpt_uop_lrs2_rtype;
  reg  r_xcpt_uop_frs3_en;
  reg  r_xcpt_uop_fp_val;
  reg  r_xcpt_uop_fp_single;
  reg  r_xcpt_uop_xcpt_if;
  reg  r_xcpt_uop_replay_if;
  reg [63:0] r_xcpt_uop_debug_wdata;
  reg [31:0] r_xcpt_uop_debug_events_fetch_seq;
  reg [39:0] r_xcpt_badvaddr;
  wire  T_23559 = io_dis_valids_0 | io_dis_valids_1; // @[rob.scala 260:32]
  wire [39:0] T_23562 = {{3'd0}, io_dis_uops_0_pc[39:3]}; // @[rob.scala 931:42]
  wire  T_23563 = rob_tail[0]; // @[rob.scala 932:25]
  wire [4:0] T_23565 = {{1'd0}, rob_tail[4:1]}; // @[rob.scala 934:29]
  wire  T_23568 = ~T_23563; // @[rob.scala 933:10]
  wire [5:0] T_23573 = {{1'd0}, io_get_pc_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_23574 = T_23573[0]; // @[rob.scala 913:37]
  wire [5:0] T_23576 = {{1'd0}, T_23573[5:1]}; // @[rob.scala 913:58]
  wire  T_23578 = T_23576 == 6'hb; // @[util.scala 75:28]
  wire [5:0] T_23582 = T_23576 + 6'h1; // @[util.scala 76:35]
  wire [5:0] T_23583 = T_23578 ? 6'h0 : T_23582; // @[util.scala 76:13]
  wire [5:0] T_23586 = T_23574 ? T_23583 : T_23576; // @[rob.scala 913:29]
  wire [39:0] T_23589 = {T_23555_T_23587_data, 3'h0}; // @[rob.scala 915:39]
  wire [39:0] T_23594 = {T_23558_T_23592_data, 3'h0}; // @[rob.scala 916:48]
  wire [39:0] T_23600 = T_23574 ? T_23594 : T_23589; // @[rob.scala 920:24]
  wire [39:0] T_23602 = T_23574 ? T_23589 : T_23594; // @[rob.scala 921:24]
  wire [63:0] T_23596 = {{24'd0}, T_23600}; // @[rob.scala 918:28 rob.scala 920:18]
  wire [39:0] T_23603 = T_23596[39:0]; // @[rob.scala 922:40]
  wire  T_23604 = T_23603[39]; // @[util.scala 114:43]
  wire [23:0] T_23608 = T_23604 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] curr_row_pc = {T_23608,T_23603}; // @[Cat.scala 20:58]
  wire [63:0] T_23598 = {{24'd0}, T_23602}; // @[rob.scala 919:28 rob.scala 921:18]
  wire [39:0] T_23609 = T_23598[39:0]; // @[rob.scala 923:40]
  wire  T_23610 = T_23609[39]; // @[util.scala 114:43]
  wire [23:0] T_23614 = T_23610 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] next_row_pc = {T_23614,T_23609}; // @[Cat.scala 20:58]
  wire  T_23615 = io_get_pc_rob_idx[0]; // @[rob.scala 227:38]
  wire [2:0] T_23617 = {T_23615,2'h0}; // @[Cat.scala 20:58]
  wire [63:0] _GEN_28820 = {{61'd0}, T_23617}; // @[rob.scala 268:37]
  wire [63:0] T_23619 = curr_row_pc + _GEN_28820; // @[rob.scala 268:37]
  wire  T_43916 = T_23573 == 6'h17; // @[util.scala 75:28]
  wire [5:0] T_43920 = T_23573 + 6'h1; // @[util.scala 76:35]
  wire [5:0] T_43921 = T_43916 ? 6'h0 : T_43920; // @[util.scala 76:13]
  reg  T_35634_23;
  reg  T_35634_22;
  reg  T_35634_21;
  reg  T_35634_20;
  reg  T_35634_19;
  reg  T_35634_18;
  reg  T_35634_17;
  reg  T_35634_16;
  reg  T_35634_15;
  reg  T_35634_14;
  reg  T_35634_13;
  reg  T_35634_12;
  reg  T_35634_11;
  reg  T_35634_10;
  reg  T_35634_9;
  reg  T_35634_8;
  reg  T_35634_7;
  reg  T_35634_6;
  reg  T_35634_5;
  reg  T_35634_4;
  reg  T_35634_3;
  reg  T_35634_2;
  reg  T_35634_1;
  reg  T_35634_0;
  wire  _GEN_22316 = 6'h1 == T_43921 ? T_35634_1 : T_35634_0; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22317 = 6'h2 == T_43921 ? T_35634_2 : _GEN_22316; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22318 = 6'h3 == T_43921 ? T_35634_3 : _GEN_22317; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22319 = 6'h4 == T_43921 ? T_35634_4 : _GEN_22318; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22320 = 6'h5 == T_43921 ? T_35634_5 : _GEN_22319; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22321 = 6'h6 == T_43921 ? T_35634_6 : _GEN_22320; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22322 = 6'h7 == T_43921 ? T_35634_7 : _GEN_22321; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22323 = 6'h8 == T_43921 ? T_35634_8 : _GEN_22322; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22324 = 6'h9 == T_43921 ? T_35634_9 : _GEN_22323; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22325 = 6'ha == T_43921 ? T_35634_10 : _GEN_22324; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22326 = 6'hb == T_43921 ? T_35634_11 : _GEN_22325; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22327 = 6'hc == T_43921 ? T_35634_12 : _GEN_22326; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22328 = 6'hd == T_43921 ? T_35634_13 : _GEN_22327; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22329 = 6'he == T_43921 ? T_35634_14 : _GEN_22328; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22330 = 6'hf == T_43921 ? T_35634_15 : _GEN_22329; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22331 = 6'h10 == T_43921 ? T_35634_16 : _GEN_22330; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22332 = 6'h11 == T_43921 ? T_35634_17 : _GEN_22331; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22333 = 6'h12 == T_43921 ? T_35634_18 : _GEN_22332; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22334 = 6'h13 == T_43921 ? T_35634_19 : _GEN_22333; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22335 = 6'h14 == T_43921 ? T_35634_20 : _GEN_22334; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22336 = 6'h15 == T_43921 ? T_35634_21 : _GEN_22335; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_22337 = 6'h16 == T_43921 ? T_35634_22 : _GEN_22336; // @[rob.scala 509:28 rob.scala 509:28]
  wire  rob_brt_vals_1 = 6'h17 == T_43921 ? T_35634_23 : _GEN_22337; // @[rob.scala 509:28 rob.scala 509:28]
  reg  T_23706_23;
  reg  T_23706_22;
  reg  T_23706_21;
  reg  T_23706_20;
  reg  T_23706_19;
  reg  T_23706_18;
  reg  T_23706_17;
  reg  T_23706_16;
  reg  T_23706_15;
  reg  T_23706_14;
  reg  T_23706_13;
  reg  T_23706_12;
  reg  T_23706_11;
  reg  T_23706_10;
  reg  T_23706_9;
  reg  T_23706_8;
  reg  T_23706_7;
  reg  T_23706_6;
  reg  T_23706_5;
  reg  T_23706_4;
  reg  T_23706_3;
  reg  T_23706_2;
  reg  T_23706_1;
  reg  T_23706_0;
  wire  _GEN_8173 = 6'h1 == T_43921 ? T_23706_1 : T_23706_0; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8174 = 6'h2 == T_43921 ? T_23706_2 : _GEN_8173; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8175 = 6'h3 == T_43921 ? T_23706_3 : _GEN_8174; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8176 = 6'h4 == T_43921 ? T_23706_4 : _GEN_8175; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8177 = 6'h5 == T_43921 ? T_23706_5 : _GEN_8176; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8178 = 6'h6 == T_43921 ? T_23706_6 : _GEN_8177; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8179 = 6'h7 == T_43921 ? T_23706_7 : _GEN_8178; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8180 = 6'h8 == T_43921 ? T_23706_8 : _GEN_8179; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8181 = 6'h9 == T_43921 ? T_23706_9 : _GEN_8180; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8182 = 6'ha == T_43921 ? T_23706_10 : _GEN_8181; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8183 = 6'hb == T_43921 ? T_23706_11 : _GEN_8182; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8184 = 6'hc == T_43921 ? T_23706_12 : _GEN_8183; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8185 = 6'hd == T_43921 ? T_23706_13 : _GEN_8184; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8186 = 6'he == T_43921 ? T_23706_14 : _GEN_8185; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8187 = 6'hf == T_43921 ? T_23706_15 : _GEN_8186; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8188 = 6'h10 == T_43921 ? T_23706_16 : _GEN_8187; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8189 = 6'h11 == T_43921 ? T_23706_17 : _GEN_8188; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8190 = 6'h12 == T_43921 ? T_23706_18 : _GEN_8189; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8191 = 6'h13 == T_43921 ? T_23706_19 : _GEN_8190; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8192 = 6'h14 == T_43921 ? T_23706_20 : _GEN_8191; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8193 = 6'h15 == T_43921 ? T_23706_21 : _GEN_8192; // @[rob.scala 509:28 rob.scala 509:28]
  wire  _GEN_8194 = 6'h16 == T_43921 ? T_23706_22 : _GEN_8193; // @[rob.scala 509:28 rob.scala 509:28]
  wire  rob_brt_vals_0 = 6'h17 == T_43921 ? T_23706_23 : _GEN_8194; // @[rob.scala 509:28 rob.scala 509:28]
  wire [1:0] T_23620 = {rob_brt_vals_1,rob_brt_vals_0};
  wire  T_23621 = T_23620[0]; // @[OneHot.scala 35:40]
  wire  next_bank_idx = T_23621 ? 1'h0 : 1'h1; // @[Mux.scala 31:69]
  wire  rob_pc_hob_next_val = rob_brt_vals_0 | rob_brt_vals_1; // @[rob.scala 273:51]
  wire [1:0] T_23625 = {io_dis_valids_1,io_dis_valids_0};
  wire  T_23626 = T_23625[0]; // @[OneHot.scala 35:40]
  wire  bypass_next_bank_idx = T_23626 ? 1'h0 : 1'h1; // @[Mux.scala 31:69]
  wire [39:0] T_23634 = $signed(io_dis_uops_0_pc) & -40'sh8;
  wire [2:0] T_23636 = {bypass_next_bank_idx,2'h0}; // @[Cat.scala 20:58]
  wire [39:0] _GEN_28823 = {{37'd0}, T_23636}; // @[rob.scala 276:97]
  wire [39:0] bypass_next_pc = T_23634 + _GEN_28823; // @[rob.scala 276:97]
  wire [2:0] T_23641 = {next_bank_idx,2'h0}; // @[Cat.scala 20:58]
  wire [63:0] _GEN_28824 = {{61'd0}, T_23641}; // @[rob.scala 281:40]
  wire [63:0] T_23643 = next_row_pc + _GEN_28824; // @[rob.scala 281:40]
  wire [63:0] T_23644 = rob_pc_hob_next_val ? T_23643 : {{24'd0}, bypass_next_pc}; // @[rob.scala 280:28]
  reg  r_partial_row;
  wire  T_23652 = T_23559 & io_dis_new_packet; // @[rob.scala 297:36]
  wire  T_23657 = ~io_dis_new_packet; // @[rob.scala 303:44]
  wire  T_23658 = T_23559 & T_23657; // @[rob.scala 303:41]
  wire  T_23660 = ~T_23652; // @[rob.scala 298:4]
  wire  T_23661 = T_23660 & T_23658; // @[rob.scala 304:4]
  wire [1:0] T_48121 = {io_com_valids_1,io_com_valids_0};
  wire  T_48123 = T_48121 != 2'h0; // @[rob.scala 715:53]
  wire  _GEN_18350 = 5'h1 == rob_head ? T_35634_1 : T_35634_0; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18351 = 5'h2 == rob_head ? T_35634_2 : _GEN_18350; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18352 = 5'h3 == rob_head ? T_35634_3 : _GEN_18351; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18353 = 5'h4 == rob_head ? T_35634_4 : _GEN_18352; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18354 = 5'h5 == rob_head ? T_35634_5 : _GEN_18353; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18355 = 5'h6 == rob_head ? T_35634_6 : _GEN_18354; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18356 = 5'h7 == rob_head ? T_35634_7 : _GEN_18355; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18357 = 5'h8 == rob_head ? T_35634_8 : _GEN_18356; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18358 = 5'h9 == rob_head ? T_35634_9 : _GEN_18357; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18359 = 5'ha == rob_head ? T_35634_10 : _GEN_18358; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18360 = 5'hb == rob_head ? T_35634_11 : _GEN_18359; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18361 = 5'hc == rob_head ? T_35634_12 : _GEN_18360; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18362 = 5'hd == rob_head ? T_35634_13 : _GEN_18361; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18363 = 5'he == rob_head ? T_35634_14 : _GEN_18362; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18364 = 5'hf == rob_head ? T_35634_15 : _GEN_18363; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18365 = 5'h10 == rob_head ? T_35634_16 : _GEN_18364; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18366 = 5'h11 == rob_head ? T_35634_17 : _GEN_18365; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18367 = 5'h12 == rob_head ? T_35634_18 : _GEN_18366; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18368 = 5'h13 == rob_head ? T_35634_19 : _GEN_18367; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18369 = 5'h14 == rob_head ? T_35634_20 : _GEN_18368; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18370 = 5'h15 == rob_head ? T_35634_21 : _GEN_18369; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_18371 = 5'h16 == rob_head ? T_35634_22 : _GEN_18370; // @[rob.scala 433:51 rob.scala 433:51]
  wire  rob_head_vals_1 = 5'h17 == rob_head ? T_35634_23 : _GEN_18371; // @[rob.scala 433:51 rob.scala 433:51]
  wire  T_41021 = ~T_35638_T_41019_data; // @[rob.scala 439:45]
  wire  T_41022 = rob_head_vals_1 & T_41021; // @[rob.scala 439:42]
  wire  T_41018 = rob_head_vals_1 & T_40239_T_41017_data; // @[rob.scala 433:51]
  wire  T_47559 = ~T_41018; // @[rob.scala 585:48]
  wire  T_47560 = T_41022 & T_47559; // @[rob.scala 585:45]
  wire  _GEN_4207 = 5'h1 == rob_head ? T_23706_1 : T_23706_0; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4208 = 5'h2 == rob_head ? T_23706_2 : _GEN_4207; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4209 = 5'h3 == rob_head ? T_23706_3 : _GEN_4208; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4210 = 5'h4 == rob_head ? T_23706_4 : _GEN_4209; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4211 = 5'h5 == rob_head ? T_23706_5 : _GEN_4210; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4212 = 5'h6 == rob_head ? T_23706_6 : _GEN_4211; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4213 = 5'h7 == rob_head ? T_23706_7 : _GEN_4212; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4214 = 5'h8 == rob_head ? T_23706_8 : _GEN_4213; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4215 = 5'h9 == rob_head ? T_23706_9 : _GEN_4214; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4216 = 5'ha == rob_head ? T_23706_10 : _GEN_4215; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4217 = 5'hb == rob_head ? T_23706_11 : _GEN_4216; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4218 = 5'hc == rob_head ? T_23706_12 : _GEN_4217; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4219 = 5'hd == rob_head ? T_23706_13 : _GEN_4218; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4220 = 5'he == rob_head ? T_23706_14 : _GEN_4219; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4221 = 5'hf == rob_head ? T_23706_15 : _GEN_4220; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4222 = 5'h10 == rob_head ? T_23706_16 : _GEN_4221; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4223 = 5'h11 == rob_head ? T_23706_17 : _GEN_4222; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4224 = 5'h12 == rob_head ? T_23706_18 : _GEN_4223; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4225 = 5'h13 == rob_head ? T_23706_19 : _GEN_4224; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4226 = 5'h14 == rob_head ? T_23706_20 : _GEN_4225; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4227 = 5'h15 == rob_head ? T_23706_21 : _GEN_4226; // @[rob.scala 433:51 rob.scala 433:51]
  wire  _GEN_4228 = 5'h16 == rob_head ? T_23706_22 : _GEN_4227; // @[rob.scala 433:51 rob.scala 433:51]
  wire  rob_head_vals_0 = 5'h17 == rob_head ? T_23706_23 : _GEN_4228; // @[rob.scala 433:51 rob.scala 433:51]
  wire  T_29093 = ~T_23710_T_29091_data; // @[rob.scala 439:45]
  wire  T_29094 = rob_head_vals_0 & T_29093; // @[rob.scala 439:42]
  wire  T_47548 = ~T_29094; // @[rob.scala 587:31]
  wire  T_29090 = rob_head_vals_0 & T_28311_T_29089_data; // @[rob.scala 433:51]
  wire  T_47549 = T_47548 | T_29090; // @[rob.scala 587:46]
  wire  T_47550 = rob_head_vals_0 & T_47549; // @[rob.scala 586:48]
  wire  T_47529 = rob_state != 2'h1; // @[rob.scala 574:34]
  wire  T_47530 = rob_state != 2'h3; // @[rob.scala 574:62]
  wire  T_47531 = T_47529 & T_47530; // @[rob.scala 574:48]
  wire  T_47551 = T_47550 | T_47531; // @[rob.scala 587:74]
  wire  T_47562 = ~T_47551; // @[rob.scala 585:75]
  wire  T_47563 = T_47560 & T_47562; // @[rob.scala 585:72]
  wire  T_47542 = ~T_29090; // @[rob.scala 585:48]
  wire  T_47543 = T_29094 & T_47542; // @[rob.scala 585:45]
  wire  T_47545 = ~T_47531; // @[rob.scala 585:75]
  wire  T_47546 = T_47543 & T_47545; // @[rob.scala 585:72]
  wire [1:0] T_48124 = {T_47563,T_47546};
  wire [1:0] T_48125 = {rob_head_vals_1,rob_head_vals_0};
  wire [1:0] T_48126 = T_48124 ^ T_48125; // @[rob.scala 716:52]
  wire  T_48128 = T_48126 == 2'h0; // @[rob.scala 716:76]
  wire  T_48129 = T_48123 & T_48128; // @[rob.scala 715:66]
  wire  T_48130 = rob_head == rob_tail; // @[rob.scala 717:59]
  wire  T_48131 = r_partial_row & T_48130; // @[rob.scala 717:47]
  wire  T_48133 = ~T_48131; // @[rob.scala 717:31]
  wire  T_48134 = T_48129 & T_48133; // @[rob.scala 716:89]
  wire  T_23670 = io_dis_valids_0 & io_dis_uops_0_is_unique; // @[rob.scala 322:24]
  wire  T_23671 = io_dis_valids_1 & io_dis_uops_1_is_unique; // @[rob.scala 322:24]
  reg  T_26182_0_valid;
  reg [1:0] T_26182_0_iw_state;
  reg [8:0] T_26182_0_uopc;
  reg [31:0] T_26182_0_inst;
  reg [39:0] T_26182_0_pc;
  reg [7:0] T_26182_0_fu_code;
  reg [3:0] T_26182_0_ctrl_br_type;
  reg [1:0] T_26182_0_ctrl_op1_sel;
  reg [2:0] T_26182_0_ctrl_op2_sel;
  reg [2:0] T_26182_0_ctrl_imm_sel;
  reg [3:0] T_26182_0_ctrl_op_fcn;
  reg  T_26182_0_ctrl_fcn_dw;
  reg  T_26182_0_ctrl_rf_wen;
  reg [2:0] T_26182_0_ctrl_csr_cmd;
  reg  T_26182_0_ctrl_is_load;
  reg  T_26182_0_ctrl_is_sta;
  reg  T_26182_0_ctrl_is_std;
  reg [1:0] T_26182_0_wakeup_delay;
  reg  T_26182_0_allocate_brtag;
  reg  T_26182_0_is_br_or_jmp;
  reg  T_26182_0_is_jump;
  reg  T_26182_0_is_jal;
  reg  T_26182_0_is_ret;
  reg  T_26182_0_is_call;
  reg [7:0] T_26182_0_br_mask;
  reg [2:0] T_26182_0_br_tag;
  reg  T_26182_0_br_prediction_bpd_predict_val;
  reg  T_26182_0_br_prediction_bpd_predict_taken;
  reg  T_26182_0_br_prediction_btb_hit;
  reg  T_26182_0_br_prediction_btb_predicted;
  reg  T_26182_0_br_prediction_is_br_or_jalr;
  reg  T_26182_0_stat_brjmp_mispredicted;
  reg  T_26182_0_stat_btb_made_pred;
  reg  T_26182_0_stat_btb_mispredicted;
  reg  T_26182_0_stat_bpd_made_pred;
  reg  T_26182_0_stat_bpd_mispredicted;
  reg [2:0] T_26182_0_fetch_pc_lob;
  reg [19:0] T_26182_0_imm_packed;
  reg [11:0] T_26182_0_csr_addr;
  reg [5:0] T_26182_0_rob_idx;
  reg [3:0] T_26182_0_ldq_idx;
  reg [3:0] T_26182_0_stq_idx;
  reg [4:0] T_26182_0_brob_idx;
  reg [6:0] T_26182_0_pdst;
  reg [6:0] T_26182_0_pop1;
  reg [6:0] T_26182_0_pop2;
  reg [6:0] T_26182_0_pop3;
  reg  T_26182_0_prs1_busy;
  reg  T_26182_0_prs2_busy;
  reg  T_26182_0_prs3_busy;
  reg [6:0] T_26182_0_stale_pdst;
  reg  T_26182_0_exception;
  reg [63:0] T_26182_0_exc_cause;
  reg  T_26182_0_bypassable;
  reg [3:0] T_26182_0_mem_cmd;
  reg [2:0] T_26182_0_mem_typ;
  reg  T_26182_0_is_fence;
  reg  T_26182_0_is_fencei;
  reg  T_26182_0_is_store;
  reg  T_26182_0_is_amo;
  reg  T_26182_0_is_load;
  reg  T_26182_0_is_unique;
  reg  T_26182_0_flush_on_commit;
  reg [5:0] T_26182_0_ldst;
  reg [5:0] T_26182_0_lrs1;
  reg [5:0] T_26182_0_lrs2;
  reg [5:0] T_26182_0_lrs3;
  reg  T_26182_0_ldst_val;
  reg [1:0] T_26182_0_dst_rtype;
  reg [1:0] T_26182_0_lrs1_rtype;
  reg [1:0] T_26182_0_lrs2_rtype;
  reg  T_26182_0_frs3_en;
  reg  T_26182_0_fp_val;
  reg  T_26182_0_fp_single;
  reg  T_26182_0_xcpt_if;
  reg  T_26182_0_replay_if;
  reg [63:0] T_26182_0_debug_wdata;
  reg [31:0] T_26182_0_debug_events_fetch_seq;
  reg  T_26182_1_valid;
  reg [1:0] T_26182_1_iw_state;
  reg [8:0] T_26182_1_uopc;
  reg [31:0] T_26182_1_inst;
  reg [39:0] T_26182_1_pc;
  reg [7:0] T_26182_1_fu_code;
  reg [3:0] T_26182_1_ctrl_br_type;
  reg [1:0] T_26182_1_ctrl_op1_sel;
  reg [2:0] T_26182_1_ctrl_op2_sel;
  reg [2:0] T_26182_1_ctrl_imm_sel;
  reg [3:0] T_26182_1_ctrl_op_fcn;
  reg  T_26182_1_ctrl_fcn_dw;
  reg  T_26182_1_ctrl_rf_wen;
  reg [2:0] T_26182_1_ctrl_csr_cmd;
  reg  T_26182_1_ctrl_is_load;
  reg  T_26182_1_ctrl_is_sta;
  reg  T_26182_1_ctrl_is_std;
  reg [1:0] T_26182_1_wakeup_delay;
  reg  T_26182_1_allocate_brtag;
  reg  T_26182_1_is_br_or_jmp;
  reg  T_26182_1_is_jump;
  reg  T_26182_1_is_jal;
  reg  T_26182_1_is_ret;
  reg  T_26182_1_is_call;
  reg [7:0] T_26182_1_br_mask;
  reg [2:0] T_26182_1_br_tag;
  reg  T_26182_1_br_prediction_bpd_predict_val;
  reg  T_26182_1_br_prediction_bpd_predict_taken;
  reg  T_26182_1_br_prediction_btb_hit;
  reg  T_26182_1_br_prediction_btb_predicted;
  reg  T_26182_1_br_prediction_is_br_or_jalr;
  reg  T_26182_1_stat_brjmp_mispredicted;
  reg  T_26182_1_stat_btb_made_pred;
  reg  T_26182_1_stat_btb_mispredicted;
  reg  T_26182_1_stat_bpd_made_pred;
  reg  T_26182_1_stat_bpd_mispredicted;
  reg [2:0] T_26182_1_fetch_pc_lob;
  reg [19:0] T_26182_1_imm_packed;
  reg [11:0] T_26182_1_csr_addr;
  reg [5:0] T_26182_1_rob_idx;
  reg [3:0] T_26182_1_ldq_idx;
  reg [3:0] T_26182_1_stq_idx;
  reg [4:0] T_26182_1_brob_idx;
  reg [6:0] T_26182_1_pdst;
  reg [6:0] T_26182_1_pop1;
  reg [6:0] T_26182_1_pop2;
  reg [6:0] T_26182_1_pop3;
  reg  T_26182_1_prs1_busy;
  reg  T_26182_1_prs2_busy;
  reg  T_26182_1_prs3_busy;
  reg [6:0] T_26182_1_stale_pdst;
  reg  T_26182_1_exception;
  reg [63:0] T_26182_1_exc_cause;
  reg  T_26182_1_bypassable;
  reg [3:0] T_26182_1_mem_cmd;
  reg [2:0] T_26182_1_mem_typ;
  reg  T_26182_1_is_fence;
  reg  T_26182_1_is_fencei;
  reg  T_26182_1_is_store;
  reg  T_26182_1_is_amo;
  reg  T_26182_1_is_load;
  reg  T_26182_1_is_unique;
  reg  T_26182_1_flush_on_commit;
  reg [5:0] T_26182_1_ldst;
  reg [5:0] T_26182_1_lrs1;
  reg [5:0] T_26182_1_lrs2;
  reg [5:0] T_26182_1_lrs3;
  reg  T_26182_1_ldst_val;
  reg [1:0] T_26182_1_dst_rtype;
  reg [1:0] T_26182_1_lrs1_rtype;
  reg [1:0] T_26182_1_lrs2_rtype;
  reg  T_26182_1_frs3_en;
  reg  T_26182_1_fp_val;
  reg  T_26182_1_fp_single;
  reg  T_26182_1_xcpt_if;
  reg  T_26182_1_replay_if;
  reg [63:0] T_26182_1_debug_wdata;
  reg [31:0] T_26182_1_debug_events_fetch_seq;
  reg  T_26182_2_valid;
  reg [1:0] T_26182_2_iw_state;
  reg [8:0] T_26182_2_uopc;
  reg [31:0] T_26182_2_inst;
  reg [39:0] T_26182_2_pc;
  reg [7:0] T_26182_2_fu_code;
  reg [3:0] T_26182_2_ctrl_br_type;
  reg [1:0] T_26182_2_ctrl_op1_sel;
  reg [2:0] T_26182_2_ctrl_op2_sel;
  reg [2:0] T_26182_2_ctrl_imm_sel;
  reg [3:0] T_26182_2_ctrl_op_fcn;
  reg  T_26182_2_ctrl_fcn_dw;
  reg  T_26182_2_ctrl_rf_wen;
  reg [2:0] T_26182_2_ctrl_csr_cmd;
  reg  T_26182_2_ctrl_is_load;
  reg  T_26182_2_ctrl_is_sta;
  reg  T_26182_2_ctrl_is_std;
  reg [1:0] T_26182_2_wakeup_delay;
  reg  T_26182_2_allocate_brtag;
  reg  T_26182_2_is_br_or_jmp;
  reg  T_26182_2_is_jump;
  reg  T_26182_2_is_jal;
  reg  T_26182_2_is_ret;
  reg  T_26182_2_is_call;
  reg [7:0] T_26182_2_br_mask;
  reg [2:0] T_26182_2_br_tag;
  reg  T_26182_2_br_prediction_bpd_predict_val;
  reg  T_26182_2_br_prediction_bpd_predict_taken;
  reg  T_26182_2_br_prediction_btb_hit;
  reg  T_26182_2_br_prediction_btb_predicted;
  reg  T_26182_2_br_prediction_is_br_or_jalr;
  reg  T_26182_2_stat_brjmp_mispredicted;
  reg  T_26182_2_stat_btb_made_pred;
  reg  T_26182_2_stat_btb_mispredicted;
  reg  T_26182_2_stat_bpd_made_pred;
  reg  T_26182_2_stat_bpd_mispredicted;
  reg [2:0] T_26182_2_fetch_pc_lob;
  reg [19:0] T_26182_2_imm_packed;
  reg [11:0] T_26182_2_csr_addr;
  reg [5:0] T_26182_2_rob_idx;
  reg [3:0] T_26182_2_ldq_idx;
  reg [3:0] T_26182_2_stq_idx;
  reg [4:0] T_26182_2_brob_idx;
  reg [6:0] T_26182_2_pdst;
  reg [6:0] T_26182_2_pop1;
  reg [6:0] T_26182_2_pop2;
  reg [6:0] T_26182_2_pop3;
  reg  T_26182_2_prs1_busy;
  reg  T_26182_2_prs2_busy;
  reg  T_26182_2_prs3_busy;
  reg [6:0] T_26182_2_stale_pdst;
  reg  T_26182_2_exception;
  reg [63:0] T_26182_2_exc_cause;
  reg  T_26182_2_bypassable;
  reg [3:0] T_26182_2_mem_cmd;
  reg [2:0] T_26182_2_mem_typ;
  reg  T_26182_2_is_fence;
  reg  T_26182_2_is_fencei;
  reg  T_26182_2_is_store;
  reg  T_26182_2_is_amo;
  reg  T_26182_2_is_load;
  reg  T_26182_2_is_unique;
  reg  T_26182_2_flush_on_commit;
  reg [5:0] T_26182_2_ldst;
  reg [5:0] T_26182_2_lrs1;
  reg [5:0] T_26182_2_lrs2;
  reg [5:0] T_26182_2_lrs3;
  reg  T_26182_2_ldst_val;
  reg [1:0] T_26182_2_dst_rtype;
  reg [1:0] T_26182_2_lrs1_rtype;
  reg [1:0] T_26182_2_lrs2_rtype;
  reg  T_26182_2_frs3_en;
  reg  T_26182_2_fp_val;
  reg  T_26182_2_fp_single;
  reg  T_26182_2_xcpt_if;
  reg  T_26182_2_replay_if;
  reg [63:0] T_26182_2_debug_wdata;
  reg [31:0] T_26182_2_debug_events_fetch_seq;
  reg  T_26182_3_valid;
  reg [1:0] T_26182_3_iw_state;
  reg [8:0] T_26182_3_uopc;
  reg [31:0] T_26182_3_inst;
  reg [39:0] T_26182_3_pc;
  reg [7:0] T_26182_3_fu_code;
  reg [3:0] T_26182_3_ctrl_br_type;
  reg [1:0] T_26182_3_ctrl_op1_sel;
  reg [2:0] T_26182_3_ctrl_op2_sel;
  reg [2:0] T_26182_3_ctrl_imm_sel;
  reg [3:0] T_26182_3_ctrl_op_fcn;
  reg  T_26182_3_ctrl_fcn_dw;
  reg  T_26182_3_ctrl_rf_wen;
  reg [2:0] T_26182_3_ctrl_csr_cmd;
  reg  T_26182_3_ctrl_is_load;
  reg  T_26182_3_ctrl_is_sta;
  reg  T_26182_3_ctrl_is_std;
  reg [1:0] T_26182_3_wakeup_delay;
  reg  T_26182_3_allocate_brtag;
  reg  T_26182_3_is_br_or_jmp;
  reg  T_26182_3_is_jump;
  reg  T_26182_3_is_jal;
  reg  T_26182_3_is_ret;
  reg  T_26182_3_is_call;
  reg [7:0] T_26182_3_br_mask;
  reg [2:0] T_26182_3_br_tag;
  reg  T_26182_3_br_prediction_bpd_predict_val;
  reg  T_26182_3_br_prediction_bpd_predict_taken;
  reg  T_26182_3_br_prediction_btb_hit;
  reg  T_26182_3_br_prediction_btb_predicted;
  reg  T_26182_3_br_prediction_is_br_or_jalr;
  reg  T_26182_3_stat_brjmp_mispredicted;
  reg  T_26182_3_stat_btb_made_pred;
  reg  T_26182_3_stat_btb_mispredicted;
  reg  T_26182_3_stat_bpd_made_pred;
  reg  T_26182_3_stat_bpd_mispredicted;
  reg [2:0] T_26182_3_fetch_pc_lob;
  reg [19:0] T_26182_3_imm_packed;
  reg [11:0] T_26182_3_csr_addr;
  reg [5:0] T_26182_3_rob_idx;
  reg [3:0] T_26182_3_ldq_idx;
  reg [3:0] T_26182_3_stq_idx;
  reg [4:0] T_26182_3_brob_idx;
  reg [6:0] T_26182_3_pdst;
  reg [6:0] T_26182_3_pop1;
  reg [6:0] T_26182_3_pop2;
  reg [6:0] T_26182_3_pop3;
  reg  T_26182_3_prs1_busy;
  reg  T_26182_3_prs2_busy;
  reg  T_26182_3_prs3_busy;
  reg [6:0] T_26182_3_stale_pdst;
  reg  T_26182_3_exception;
  reg [63:0] T_26182_3_exc_cause;
  reg  T_26182_3_bypassable;
  reg [3:0] T_26182_3_mem_cmd;
  reg [2:0] T_26182_3_mem_typ;
  reg  T_26182_3_is_fence;
  reg  T_26182_3_is_fencei;
  reg  T_26182_3_is_store;
  reg  T_26182_3_is_amo;
  reg  T_26182_3_is_load;
  reg  T_26182_3_is_unique;
  reg  T_26182_3_flush_on_commit;
  reg [5:0] T_26182_3_ldst;
  reg [5:0] T_26182_3_lrs1;
  reg [5:0] T_26182_3_lrs2;
  reg [5:0] T_26182_3_lrs3;
  reg  T_26182_3_ldst_val;
  reg [1:0] T_26182_3_dst_rtype;
  reg [1:0] T_26182_3_lrs1_rtype;
  reg [1:0] T_26182_3_lrs2_rtype;
  reg  T_26182_3_frs3_en;
  reg  T_26182_3_fp_val;
  reg  T_26182_3_fp_single;
  reg  T_26182_3_xcpt_if;
  reg  T_26182_3_replay_if;
  reg [63:0] T_26182_3_debug_wdata;
  reg [31:0] T_26182_3_debug_events_fetch_seq;
  reg  T_26182_4_valid;
  reg [1:0] T_26182_4_iw_state;
  reg [8:0] T_26182_4_uopc;
  reg [31:0] T_26182_4_inst;
  reg [39:0] T_26182_4_pc;
  reg [7:0] T_26182_4_fu_code;
  reg [3:0] T_26182_4_ctrl_br_type;
  reg [1:0] T_26182_4_ctrl_op1_sel;
  reg [2:0] T_26182_4_ctrl_op2_sel;
  reg [2:0] T_26182_4_ctrl_imm_sel;
  reg [3:0] T_26182_4_ctrl_op_fcn;
  reg  T_26182_4_ctrl_fcn_dw;
  reg  T_26182_4_ctrl_rf_wen;
  reg [2:0] T_26182_4_ctrl_csr_cmd;
  reg  T_26182_4_ctrl_is_load;
  reg  T_26182_4_ctrl_is_sta;
  reg  T_26182_4_ctrl_is_std;
  reg [1:0] T_26182_4_wakeup_delay;
  reg  T_26182_4_allocate_brtag;
  reg  T_26182_4_is_br_or_jmp;
  reg  T_26182_4_is_jump;
  reg  T_26182_4_is_jal;
  reg  T_26182_4_is_ret;
  reg  T_26182_4_is_call;
  reg [7:0] T_26182_4_br_mask;
  reg [2:0] T_26182_4_br_tag;
  reg  T_26182_4_br_prediction_bpd_predict_val;
  reg  T_26182_4_br_prediction_bpd_predict_taken;
  reg  T_26182_4_br_prediction_btb_hit;
  reg  T_26182_4_br_prediction_btb_predicted;
  reg  T_26182_4_br_prediction_is_br_or_jalr;
  reg  T_26182_4_stat_brjmp_mispredicted;
  reg  T_26182_4_stat_btb_made_pred;
  reg  T_26182_4_stat_btb_mispredicted;
  reg  T_26182_4_stat_bpd_made_pred;
  reg  T_26182_4_stat_bpd_mispredicted;
  reg [2:0] T_26182_4_fetch_pc_lob;
  reg [19:0] T_26182_4_imm_packed;
  reg [11:0] T_26182_4_csr_addr;
  reg [5:0] T_26182_4_rob_idx;
  reg [3:0] T_26182_4_ldq_idx;
  reg [3:0] T_26182_4_stq_idx;
  reg [4:0] T_26182_4_brob_idx;
  reg [6:0] T_26182_4_pdst;
  reg [6:0] T_26182_4_pop1;
  reg [6:0] T_26182_4_pop2;
  reg [6:0] T_26182_4_pop3;
  reg  T_26182_4_prs1_busy;
  reg  T_26182_4_prs2_busy;
  reg  T_26182_4_prs3_busy;
  reg [6:0] T_26182_4_stale_pdst;
  reg  T_26182_4_exception;
  reg [63:0] T_26182_4_exc_cause;
  reg  T_26182_4_bypassable;
  reg [3:0] T_26182_4_mem_cmd;
  reg [2:0] T_26182_4_mem_typ;
  reg  T_26182_4_is_fence;
  reg  T_26182_4_is_fencei;
  reg  T_26182_4_is_store;
  reg  T_26182_4_is_amo;
  reg  T_26182_4_is_load;
  reg  T_26182_4_is_unique;
  reg  T_26182_4_flush_on_commit;
  reg [5:0] T_26182_4_ldst;
  reg [5:0] T_26182_4_lrs1;
  reg [5:0] T_26182_4_lrs2;
  reg [5:0] T_26182_4_lrs3;
  reg  T_26182_4_ldst_val;
  reg [1:0] T_26182_4_dst_rtype;
  reg [1:0] T_26182_4_lrs1_rtype;
  reg [1:0] T_26182_4_lrs2_rtype;
  reg  T_26182_4_frs3_en;
  reg  T_26182_4_fp_val;
  reg  T_26182_4_fp_single;
  reg  T_26182_4_xcpt_if;
  reg  T_26182_4_replay_if;
  reg [63:0] T_26182_4_debug_wdata;
  reg [31:0] T_26182_4_debug_events_fetch_seq;
  reg  T_26182_5_valid;
  reg [1:0] T_26182_5_iw_state;
  reg [8:0] T_26182_5_uopc;
  reg [31:0] T_26182_5_inst;
  reg [39:0] T_26182_5_pc;
  reg [7:0] T_26182_5_fu_code;
  reg [3:0] T_26182_5_ctrl_br_type;
  reg [1:0] T_26182_5_ctrl_op1_sel;
  reg [2:0] T_26182_5_ctrl_op2_sel;
  reg [2:0] T_26182_5_ctrl_imm_sel;
  reg [3:0] T_26182_5_ctrl_op_fcn;
  reg  T_26182_5_ctrl_fcn_dw;
  reg  T_26182_5_ctrl_rf_wen;
  reg [2:0] T_26182_5_ctrl_csr_cmd;
  reg  T_26182_5_ctrl_is_load;
  reg  T_26182_5_ctrl_is_sta;
  reg  T_26182_5_ctrl_is_std;
  reg [1:0] T_26182_5_wakeup_delay;
  reg  T_26182_5_allocate_brtag;
  reg  T_26182_5_is_br_or_jmp;
  reg  T_26182_5_is_jump;
  reg  T_26182_5_is_jal;
  reg  T_26182_5_is_ret;
  reg  T_26182_5_is_call;
  reg [7:0] T_26182_5_br_mask;
  reg [2:0] T_26182_5_br_tag;
  reg  T_26182_5_br_prediction_bpd_predict_val;
  reg  T_26182_5_br_prediction_bpd_predict_taken;
  reg  T_26182_5_br_prediction_btb_hit;
  reg  T_26182_5_br_prediction_btb_predicted;
  reg  T_26182_5_br_prediction_is_br_or_jalr;
  reg  T_26182_5_stat_brjmp_mispredicted;
  reg  T_26182_5_stat_btb_made_pred;
  reg  T_26182_5_stat_btb_mispredicted;
  reg  T_26182_5_stat_bpd_made_pred;
  reg  T_26182_5_stat_bpd_mispredicted;
  reg [2:0] T_26182_5_fetch_pc_lob;
  reg [19:0] T_26182_5_imm_packed;
  reg [11:0] T_26182_5_csr_addr;
  reg [5:0] T_26182_5_rob_idx;
  reg [3:0] T_26182_5_ldq_idx;
  reg [3:0] T_26182_5_stq_idx;
  reg [4:0] T_26182_5_brob_idx;
  reg [6:0] T_26182_5_pdst;
  reg [6:0] T_26182_5_pop1;
  reg [6:0] T_26182_5_pop2;
  reg [6:0] T_26182_5_pop3;
  reg  T_26182_5_prs1_busy;
  reg  T_26182_5_prs2_busy;
  reg  T_26182_5_prs3_busy;
  reg [6:0] T_26182_5_stale_pdst;
  reg  T_26182_5_exception;
  reg [63:0] T_26182_5_exc_cause;
  reg  T_26182_5_bypassable;
  reg [3:0] T_26182_5_mem_cmd;
  reg [2:0] T_26182_5_mem_typ;
  reg  T_26182_5_is_fence;
  reg  T_26182_5_is_fencei;
  reg  T_26182_5_is_store;
  reg  T_26182_5_is_amo;
  reg  T_26182_5_is_load;
  reg  T_26182_5_is_unique;
  reg  T_26182_5_flush_on_commit;
  reg [5:0] T_26182_5_ldst;
  reg [5:0] T_26182_5_lrs1;
  reg [5:0] T_26182_5_lrs2;
  reg [5:0] T_26182_5_lrs3;
  reg  T_26182_5_ldst_val;
  reg [1:0] T_26182_5_dst_rtype;
  reg [1:0] T_26182_5_lrs1_rtype;
  reg [1:0] T_26182_5_lrs2_rtype;
  reg  T_26182_5_frs3_en;
  reg  T_26182_5_fp_val;
  reg  T_26182_5_fp_single;
  reg  T_26182_5_xcpt_if;
  reg  T_26182_5_replay_if;
  reg [63:0] T_26182_5_debug_wdata;
  reg [31:0] T_26182_5_debug_events_fetch_seq;
  reg  T_26182_6_valid;
  reg [1:0] T_26182_6_iw_state;
  reg [8:0] T_26182_6_uopc;
  reg [31:0] T_26182_6_inst;
  reg [39:0] T_26182_6_pc;
  reg [7:0] T_26182_6_fu_code;
  reg [3:0] T_26182_6_ctrl_br_type;
  reg [1:0] T_26182_6_ctrl_op1_sel;
  reg [2:0] T_26182_6_ctrl_op2_sel;
  reg [2:0] T_26182_6_ctrl_imm_sel;
  reg [3:0] T_26182_6_ctrl_op_fcn;
  reg  T_26182_6_ctrl_fcn_dw;
  reg  T_26182_6_ctrl_rf_wen;
  reg [2:0] T_26182_6_ctrl_csr_cmd;
  reg  T_26182_6_ctrl_is_load;
  reg  T_26182_6_ctrl_is_sta;
  reg  T_26182_6_ctrl_is_std;
  reg [1:0] T_26182_6_wakeup_delay;
  reg  T_26182_6_allocate_brtag;
  reg  T_26182_6_is_br_or_jmp;
  reg  T_26182_6_is_jump;
  reg  T_26182_6_is_jal;
  reg  T_26182_6_is_ret;
  reg  T_26182_6_is_call;
  reg [7:0] T_26182_6_br_mask;
  reg [2:0] T_26182_6_br_tag;
  reg  T_26182_6_br_prediction_bpd_predict_val;
  reg  T_26182_6_br_prediction_bpd_predict_taken;
  reg  T_26182_6_br_prediction_btb_hit;
  reg  T_26182_6_br_prediction_btb_predicted;
  reg  T_26182_6_br_prediction_is_br_or_jalr;
  reg  T_26182_6_stat_brjmp_mispredicted;
  reg  T_26182_6_stat_btb_made_pred;
  reg  T_26182_6_stat_btb_mispredicted;
  reg  T_26182_6_stat_bpd_made_pred;
  reg  T_26182_6_stat_bpd_mispredicted;
  reg [2:0] T_26182_6_fetch_pc_lob;
  reg [19:0] T_26182_6_imm_packed;
  reg [11:0] T_26182_6_csr_addr;
  reg [5:0] T_26182_6_rob_idx;
  reg [3:0] T_26182_6_ldq_idx;
  reg [3:0] T_26182_6_stq_idx;
  reg [4:0] T_26182_6_brob_idx;
  reg [6:0] T_26182_6_pdst;
  reg [6:0] T_26182_6_pop1;
  reg [6:0] T_26182_6_pop2;
  reg [6:0] T_26182_6_pop3;
  reg  T_26182_6_prs1_busy;
  reg  T_26182_6_prs2_busy;
  reg  T_26182_6_prs3_busy;
  reg [6:0] T_26182_6_stale_pdst;
  reg  T_26182_6_exception;
  reg [63:0] T_26182_6_exc_cause;
  reg  T_26182_6_bypassable;
  reg [3:0] T_26182_6_mem_cmd;
  reg [2:0] T_26182_6_mem_typ;
  reg  T_26182_6_is_fence;
  reg  T_26182_6_is_fencei;
  reg  T_26182_6_is_store;
  reg  T_26182_6_is_amo;
  reg  T_26182_6_is_load;
  reg  T_26182_6_is_unique;
  reg  T_26182_6_flush_on_commit;
  reg [5:0] T_26182_6_ldst;
  reg [5:0] T_26182_6_lrs1;
  reg [5:0] T_26182_6_lrs2;
  reg [5:0] T_26182_6_lrs3;
  reg  T_26182_6_ldst_val;
  reg [1:0] T_26182_6_dst_rtype;
  reg [1:0] T_26182_6_lrs1_rtype;
  reg [1:0] T_26182_6_lrs2_rtype;
  reg  T_26182_6_frs3_en;
  reg  T_26182_6_fp_val;
  reg  T_26182_6_fp_single;
  reg  T_26182_6_xcpt_if;
  reg  T_26182_6_replay_if;
  reg [63:0] T_26182_6_debug_wdata;
  reg [31:0] T_26182_6_debug_events_fetch_seq;
  reg  T_26182_7_valid;
  reg [1:0] T_26182_7_iw_state;
  reg [8:0] T_26182_7_uopc;
  reg [31:0] T_26182_7_inst;
  reg [39:0] T_26182_7_pc;
  reg [7:0] T_26182_7_fu_code;
  reg [3:0] T_26182_7_ctrl_br_type;
  reg [1:0] T_26182_7_ctrl_op1_sel;
  reg [2:0] T_26182_7_ctrl_op2_sel;
  reg [2:0] T_26182_7_ctrl_imm_sel;
  reg [3:0] T_26182_7_ctrl_op_fcn;
  reg  T_26182_7_ctrl_fcn_dw;
  reg  T_26182_7_ctrl_rf_wen;
  reg [2:0] T_26182_7_ctrl_csr_cmd;
  reg  T_26182_7_ctrl_is_load;
  reg  T_26182_7_ctrl_is_sta;
  reg  T_26182_7_ctrl_is_std;
  reg [1:0] T_26182_7_wakeup_delay;
  reg  T_26182_7_allocate_brtag;
  reg  T_26182_7_is_br_or_jmp;
  reg  T_26182_7_is_jump;
  reg  T_26182_7_is_jal;
  reg  T_26182_7_is_ret;
  reg  T_26182_7_is_call;
  reg [7:0] T_26182_7_br_mask;
  reg [2:0] T_26182_7_br_tag;
  reg  T_26182_7_br_prediction_bpd_predict_val;
  reg  T_26182_7_br_prediction_bpd_predict_taken;
  reg  T_26182_7_br_prediction_btb_hit;
  reg  T_26182_7_br_prediction_btb_predicted;
  reg  T_26182_7_br_prediction_is_br_or_jalr;
  reg  T_26182_7_stat_brjmp_mispredicted;
  reg  T_26182_7_stat_btb_made_pred;
  reg  T_26182_7_stat_btb_mispredicted;
  reg  T_26182_7_stat_bpd_made_pred;
  reg  T_26182_7_stat_bpd_mispredicted;
  reg [2:0] T_26182_7_fetch_pc_lob;
  reg [19:0] T_26182_7_imm_packed;
  reg [11:0] T_26182_7_csr_addr;
  reg [5:0] T_26182_7_rob_idx;
  reg [3:0] T_26182_7_ldq_idx;
  reg [3:0] T_26182_7_stq_idx;
  reg [4:0] T_26182_7_brob_idx;
  reg [6:0] T_26182_7_pdst;
  reg [6:0] T_26182_7_pop1;
  reg [6:0] T_26182_7_pop2;
  reg [6:0] T_26182_7_pop3;
  reg  T_26182_7_prs1_busy;
  reg  T_26182_7_prs2_busy;
  reg  T_26182_7_prs3_busy;
  reg [6:0] T_26182_7_stale_pdst;
  reg  T_26182_7_exception;
  reg [63:0] T_26182_7_exc_cause;
  reg  T_26182_7_bypassable;
  reg [3:0] T_26182_7_mem_cmd;
  reg [2:0] T_26182_7_mem_typ;
  reg  T_26182_7_is_fence;
  reg  T_26182_7_is_fencei;
  reg  T_26182_7_is_store;
  reg  T_26182_7_is_amo;
  reg  T_26182_7_is_load;
  reg  T_26182_7_is_unique;
  reg  T_26182_7_flush_on_commit;
  reg [5:0] T_26182_7_ldst;
  reg [5:0] T_26182_7_lrs1;
  reg [5:0] T_26182_7_lrs2;
  reg [5:0] T_26182_7_lrs3;
  reg  T_26182_7_ldst_val;
  reg [1:0] T_26182_7_dst_rtype;
  reg [1:0] T_26182_7_lrs1_rtype;
  reg [1:0] T_26182_7_lrs2_rtype;
  reg  T_26182_7_frs3_en;
  reg  T_26182_7_fp_val;
  reg  T_26182_7_fp_single;
  reg  T_26182_7_xcpt_if;
  reg  T_26182_7_replay_if;
  reg [63:0] T_26182_7_debug_wdata;
  reg [31:0] T_26182_7_debug_events_fetch_seq;
  reg  T_26182_8_valid;
  reg [1:0] T_26182_8_iw_state;
  reg [8:0] T_26182_8_uopc;
  reg [31:0] T_26182_8_inst;
  reg [39:0] T_26182_8_pc;
  reg [7:0] T_26182_8_fu_code;
  reg [3:0] T_26182_8_ctrl_br_type;
  reg [1:0] T_26182_8_ctrl_op1_sel;
  reg [2:0] T_26182_8_ctrl_op2_sel;
  reg [2:0] T_26182_8_ctrl_imm_sel;
  reg [3:0] T_26182_8_ctrl_op_fcn;
  reg  T_26182_8_ctrl_fcn_dw;
  reg  T_26182_8_ctrl_rf_wen;
  reg [2:0] T_26182_8_ctrl_csr_cmd;
  reg  T_26182_8_ctrl_is_load;
  reg  T_26182_8_ctrl_is_sta;
  reg  T_26182_8_ctrl_is_std;
  reg [1:0] T_26182_8_wakeup_delay;
  reg  T_26182_8_allocate_brtag;
  reg  T_26182_8_is_br_or_jmp;
  reg  T_26182_8_is_jump;
  reg  T_26182_8_is_jal;
  reg  T_26182_8_is_ret;
  reg  T_26182_8_is_call;
  reg [7:0] T_26182_8_br_mask;
  reg [2:0] T_26182_8_br_tag;
  reg  T_26182_8_br_prediction_bpd_predict_val;
  reg  T_26182_8_br_prediction_bpd_predict_taken;
  reg  T_26182_8_br_prediction_btb_hit;
  reg  T_26182_8_br_prediction_btb_predicted;
  reg  T_26182_8_br_prediction_is_br_or_jalr;
  reg  T_26182_8_stat_brjmp_mispredicted;
  reg  T_26182_8_stat_btb_made_pred;
  reg  T_26182_8_stat_btb_mispredicted;
  reg  T_26182_8_stat_bpd_made_pred;
  reg  T_26182_8_stat_bpd_mispredicted;
  reg [2:0] T_26182_8_fetch_pc_lob;
  reg [19:0] T_26182_8_imm_packed;
  reg [11:0] T_26182_8_csr_addr;
  reg [5:0] T_26182_8_rob_idx;
  reg [3:0] T_26182_8_ldq_idx;
  reg [3:0] T_26182_8_stq_idx;
  reg [4:0] T_26182_8_brob_idx;
  reg [6:0] T_26182_8_pdst;
  reg [6:0] T_26182_8_pop1;
  reg [6:0] T_26182_8_pop2;
  reg [6:0] T_26182_8_pop3;
  reg  T_26182_8_prs1_busy;
  reg  T_26182_8_prs2_busy;
  reg  T_26182_8_prs3_busy;
  reg [6:0] T_26182_8_stale_pdst;
  reg  T_26182_8_exception;
  reg [63:0] T_26182_8_exc_cause;
  reg  T_26182_8_bypassable;
  reg [3:0] T_26182_8_mem_cmd;
  reg [2:0] T_26182_8_mem_typ;
  reg  T_26182_8_is_fence;
  reg  T_26182_8_is_fencei;
  reg  T_26182_8_is_store;
  reg  T_26182_8_is_amo;
  reg  T_26182_8_is_load;
  reg  T_26182_8_is_unique;
  reg  T_26182_8_flush_on_commit;
  reg [5:0] T_26182_8_ldst;
  reg [5:0] T_26182_8_lrs1;
  reg [5:0] T_26182_8_lrs2;
  reg [5:0] T_26182_8_lrs3;
  reg  T_26182_8_ldst_val;
  reg [1:0] T_26182_8_dst_rtype;
  reg [1:0] T_26182_8_lrs1_rtype;
  reg [1:0] T_26182_8_lrs2_rtype;
  reg  T_26182_8_frs3_en;
  reg  T_26182_8_fp_val;
  reg  T_26182_8_fp_single;
  reg  T_26182_8_xcpt_if;
  reg  T_26182_8_replay_if;
  reg [63:0] T_26182_8_debug_wdata;
  reg [31:0] T_26182_8_debug_events_fetch_seq;
  reg  T_26182_9_valid;
  reg [1:0] T_26182_9_iw_state;
  reg [8:0] T_26182_9_uopc;
  reg [31:0] T_26182_9_inst;
  reg [39:0] T_26182_9_pc;
  reg [7:0] T_26182_9_fu_code;
  reg [3:0] T_26182_9_ctrl_br_type;
  reg [1:0] T_26182_9_ctrl_op1_sel;
  reg [2:0] T_26182_9_ctrl_op2_sel;
  reg [2:0] T_26182_9_ctrl_imm_sel;
  reg [3:0] T_26182_9_ctrl_op_fcn;
  reg  T_26182_9_ctrl_fcn_dw;
  reg  T_26182_9_ctrl_rf_wen;
  reg [2:0] T_26182_9_ctrl_csr_cmd;
  reg  T_26182_9_ctrl_is_load;
  reg  T_26182_9_ctrl_is_sta;
  reg  T_26182_9_ctrl_is_std;
  reg [1:0] T_26182_9_wakeup_delay;
  reg  T_26182_9_allocate_brtag;
  reg  T_26182_9_is_br_or_jmp;
  reg  T_26182_9_is_jump;
  reg  T_26182_9_is_jal;
  reg  T_26182_9_is_ret;
  reg  T_26182_9_is_call;
  reg [7:0] T_26182_9_br_mask;
  reg [2:0] T_26182_9_br_tag;
  reg  T_26182_9_br_prediction_bpd_predict_val;
  reg  T_26182_9_br_prediction_bpd_predict_taken;
  reg  T_26182_9_br_prediction_btb_hit;
  reg  T_26182_9_br_prediction_btb_predicted;
  reg  T_26182_9_br_prediction_is_br_or_jalr;
  reg  T_26182_9_stat_brjmp_mispredicted;
  reg  T_26182_9_stat_btb_made_pred;
  reg  T_26182_9_stat_btb_mispredicted;
  reg  T_26182_9_stat_bpd_made_pred;
  reg  T_26182_9_stat_bpd_mispredicted;
  reg [2:0] T_26182_9_fetch_pc_lob;
  reg [19:0] T_26182_9_imm_packed;
  reg [11:0] T_26182_9_csr_addr;
  reg [5:0] T_26182_9_rob_idx;
  reg [3:0] T_26182_9_ldq_idx;
  reg [3:0] T_26182_9_stq_idx;
  reg [4:0] T_26182_9_brob_idx;
  reg [6:0] T_26182_9_pdst;
  reg [6:0] T_26182_9_pop1;
  reg [6:0] T_26182_9_pop2;
  reg [6:0] T_26182_9_pop3;
  reg  T_26182_9_prs1_busy;
  reg  T_26182_9_prs2_busy;
  reg  T_26182_9_prs3_busy;
  reg [6:0] T_26182_9_stale_pdst;
  reg  T_26182_9_exception;
  reg [63:0] T_26182_9_exc_cause;
  reg  T_26182_9_bypassable;
  reg [3:0] T_26182_9_mem_cmd;
  reg [2:0] T_26182_9_mem_typ;
  reg  T_26182_9_is_fence;
  reg  T_26182_9_is_fencei;
  reg  T_26182_9_is_store;
  reg  T_26182_9_is_amo;
  reg  T_26182_9_is_load;
  reg  T_26182_9_is_unique;
  reg  T_26182_9_flush_on_commit;
  reg [5:0] T_26182_9_ldst;
  reg [5:0] T_26182_9_lrs1;
  reg [5:0] T_26182_9_lrs2;
  reg [5:0] T_26182_9_lrs3;
  reg  T_26182_9_ldst_val;
  reg [1:0] T_26182_9_dst_rtype;
  reg [1:0] T_26182_9_lrs1_rtype;
  reg [1:0] T_26182_9_lrs2_rtype;
  reg  T_26182_9_frs3_en;
  reg  T_26182_9_fp_val;
  reg  T_26182_9_fp_single;
  reg  T_26182_9_xcpt_if;
  reg  T_26182_9_replay_if;
  reg [63:0] T_26182_9_debug_wdata;
  reg [31:0] T_26182_9_debug_events_fetch_seq;
  reg  T_26182_10_valid;
  reg [1:0] T_26182_10_iw_state;
  reg [8:0] T_26182_10_uopc;
  reg [31:0] T_26182_10_inst;
  reg [39:0] T_26182_10_pc;
  reg [7:0] T_26182_10_fu_code;
  reg [3:0] T_26182_10_ctrl_br_type;
  reg [1:0] T_26182_10_ctrl_op1_sel;
  reg [2:0] T_26182_10_ctrl_op2_sel;
  reg [2:0] T_26182_10_ctrl_imm_sel;
  reg [3:0] T_26182_10_ctrl_op_fcn;
  reg  T_26182_10_ctrl_fcn_dw;
  reg  T_26182_10_ctrl_rf_wen;
  reg [2:0] T_26182_10_ctrl_csr_cmd;
  reg  T_26182_10_ctrl_is_load;
  reg  T_26182_10_ctrl_is_sta;
  reg  T_26182_10_ctrl_is_std;
  reg [1:0] T_26182_10_wakeup_delay;
  reg  T_26182_10_allocate_brtag;
  reg  T_26182_10_is_br_or_jmp;
  reg  T_26182_10_is_jump;
  reg  T_26182_10_is_jal;
  reg  T_26182_10_is_ret;
  reg  T_26182_10_is_call;
  reg [7:0] T_26182_10_br_mask;
  reg [2:0] T_26182_10_br_tag;
  reg  T_26182_10_br_prediction_bpd_predict_val;
  reg  T_26182_10_br_prediction_bpd_predict_taken;
  reg  T_26182_10_br_prediction_btb_hit;
  reg  T_26182_10_br_prediction_btb_predicted;
  reg  T_26182_10_br_prediction_is_br_or_jalr;
  reg  T_26182_10_stat_brjmp_mispredicted;
  reg  T_26182_10_stat_btb_made_pred;
  reg  T_26182_10_stat_btb_mispredicted;
  reg  T_26182_10_stat_bpd_made_pred;
  reg  T_26182_10_stat_bpd_mispredicted;
  reg [2:0] T_26182_10_fetch_pc_lob;
  reg [19:0] T_26182_10_imm_packed;
  reg [11:0] T_26182_10_csr_addr;
  reg [5:0] T_26182_10_rob_idx;
  reg [3:0] T_26182_10_ldq_idx;
  reg [3:0] T_26182_10_stq_idx;
  reg [4:0] T_26182_10_brob_idx;
  reg [6:0] T_26182_10_pdst;
  reg [6:0] T_26182_10_pop1;
  reg [6:0] T_26182_10_pop2;
  reg [6:0] T_26182_10_pop3;
  reg  T_26182_10_prs1_busy;
  reg  T_26182_10_prs2_busy;
  reg  T_26182_10_prs3_busy;
  reg [6:0] T_26182_10_stale_pdst;
  reg  T_26182_10_exception;
  reg [63:0] T_26182_10_exc_cause;
  reg  T_26182_10_bypassable;
  reg [3:0] T_26182_10_mem_cmd;
  reg [2:0] T_26182_10_mem_typ;
  reg  T_26182_10_is_fence;
  reg  T_26182_10_is_fencei;
  reg  T_26182_10_is_store;
  reg  T_26182_10_is_amo;
  reg  T_26182_10_is_load;
  reg  T_26182_10_is_unique;
  reg  T_26182_10_flush_on_commit;
  reg [5:0] T_26182_10_ldst;
  reg [5:0] T_26182_10_lrs1;
  reg [5:0] T_26182_10_lrs2;
  reg [5:0] T_26182_10_lrs3;
  reg  T_26182_10_ldst_val;
  reg [1:0] T_26182_10_dst_rtype;
  reg [1:0] T_26182_10_lrs1_rtype;
  reg [1:0] T_26182_10_lrs2_rtype;
  reg  T_26182_10_frs3_en;
  reg  T_26182_10_fp_val;
  reg  T_26182_10_fp_single;
  reg  T_26182_10_xcpt_if;
  reg  T_26182_10_replay_if;
  reg [63:0] T_26182_10_debug_wdata;
  reg [31:0] T_26182_10_debug_events_fetch_seq;
  reg  T_26182_11_valid;
  reg [1:0] T_26182_11_iw_state;
  reg [8:0] T_26182_11_uopc;
  reg [31:0] T_26182_11_inst;
  reg [39:0] T_26182_11_pc;
  reg [7:0] T_26182_11_fu_code;
  reg [3:0] T_26182_11_ctrl_br_type;
  reg [1:0] T_26182_11_ctrl_op1_sel;
  reg [2:0] T_26182_11_ctrl_op2_sel;
  reg [2:0] T_26182_11_ctrl_imm_sel;
  reg [3:0] T_26182_11_ctrl_op_fcn;
  reg  T_26182_11_ctrl_fcn_dw;
  reg  T_26182_11_ctrl_rf_wen;
  reg [2:0] T_26182_11_ctrl_csr_cmd;
  reg  T_26182_11_ctrl_is_load;
  reg  T_26182_11_ctrl_is_sta;
  reg  T_26182_11_ctrl_is_std;
  reg [1:0] T_26182_11_wakeup_delay;
  reg  T_26182_11_allocate_brtag;
  reg  T_26182_11_is_br_or_jmp;
  reg  T_26182_11_is_jump;
  reg  T_26182_11_is_jal;
  reg  T_26182_11_is_ret;
  reg  T_26182_11_is_call;
  reg [7:0] T_26182_11_br_mask;
  reg [2:0] T_26182_11_br_tag;
  reg  T_26182_11_br_prediction_bpd_predict_val;
  reg  T_26182_11_br_prediction_bpd_predict_taken;
  reg  T_26182_11_br_prediction_btb_hit;
  reg  T_26182_11_br_prediction_btb_predicted;
  reg  T_26182_11_br_prediction_is_br_or_jalr;
  reg  T_26182_11_stat_brjmp_mispredicted;
  reg  T_26182_11_stat_btb_made_pred;
  reg  T_26182_11_stat_btb_mispredicted;
  reg  T_26182_11_stat_bpd_made_pred;
  reg  T_26182_11_stat_bpd_mispredicted;
  reg [2:0] T_26182_11_fetch_pc_lob;
  reg [19:0] T_26182_11_imm_packed;
  reg [11:0] T_26182_11_csr_addr;
  reg [5:0] T_26182_11_rob_idx;
  reg [3:0] T_26182_11_ldq_idx;
  reg [3:0] T_26182_11_stq_idx;
  reg [4:0] T_26182_11_brob_idx;
  reg [6:0] T_26182_11_pdst;
  reg [6:0] T_26182_11_pop1;
  reg [6:0] T_26182_11_pop2;
  reg [6:0] T_26182_11_pop3;
  reg  T_26182_11_prs1_busy;
  reg  T_26182_11_prs2_busy;
  reg  T_26182_11_prs3_busy;
  reg [6:0] T_26182_11_stale_pdst;
  reg  T_26182_11_exception;
  reg [63:0] T_26182_11_exc_cause;
  reg  T_26182_11_bypassable;
  reg [3:0] T_26182_11_mem_cmd;
  reg [2:0] T_26182_11_mem_typ;
  reg  T_26182_11_is_fence;
  reg  T_26182_11_is_fencei;
  reg  T_26182_11_is_store;
  reg  T_26182_11_is_amo;
  reg  T_26182_11_is_load;
  reg  T_26182_11_is_unique;
  reg  T_26182_11_flush_on_commit;
  reg [5:0] T_26182_11_ldst;
  reg [5:0] T_26182_11_lrs1;
  reg [5:0] T_26182_11_lrs2;
  reg [5:0] T_26182_11_lrs3;
  reg  T_26182_11_ldst_val;
  reg [1:0] T_26182_11_dst_rtype;
  reg [1:0] T_26182_11_lrs1_rtype;
  reg [1:0] T_26182_11_lrs2_rtype;
  reg  T_26182_11_frs3_en;
  reg  T_26182_11_fp_val;
  reg  T_26182_11_fp_single;
  reg  T_26182_11_xcpt_if;
  reg  T_26182_11_replay_if;
  reg [63:0] T_26182_11_debug_wdata;
  reg [31:0] T_26182_11_debug_events_fetch_seq;
  reg  T_26182_12_valid;
  reg [1:0] T_26182_12_iw_state;
  reg [8:0] T_26182_12_uopc;
  reg [31:0] T_26182_12_inst;
  reg [39:0] T_26182_12_pc;
  reg [7:0] T_26182_12_fu_code;
  reg [3:0] T_26182_12_ctrl_br_type;
  reg [1:0] T_26182_12_ctrl_op1_sel;
  reg [2:0] T_26182_12_ctrl_op2_sel;
  reg [2:0] T_26182_12_ctrl_imm_sel;
  reg [3:0] T_26182_12_ctrl_op_fcn;
  reg  T_26182_12_ctrl_fcn_dw;
  reg  T_26182_12_ctrl_rf_wen;
  reg [2:0] T_26182_12_ctrl_csr_cmd;
  reg  T_26182_12_ctrl_is_load;
  reg  T_26182_12_ctrl_is_sta;
  reg  T_26182_12_ctrl_is_std;
  reg [1:0] T_26182_12_wakeup_delay;
  reg  T_26182_12_allocate_brtag;
  reg  T_26182_12_is_br_or_jmp;
  reg  T_26182_12_is_jump;
  reg  T_26182_12_is_jal;
  reg  T_26182_12_is_ret;
  reg  T_26182_12_is_call;
  reg [7:0] T_26182_12_br_mask;
  reg [2:0] T_26182_12_br_tag;
  reg  T_26182_12_br_prediction_bpd_predict_val;
  reg  T_26182_12_br_prediction_bpd_predict_taken;
  reg  T_26182_12_br_prediction_btb_hit;
  reg  T_26182_12_br_prediction_btb_predicted;
  reg  T_26182_12_br_prediction_is_br_or_jalr;
  reg  T_26182_12_stat_brjmp_mispredicted;
  reg  T_26182_12_stat_btb_made_pred;
  reg  T_26182_12_stat_btb_mispredicted;
  reg  T_26182_12_stat_bpd_made_pred;
  reg  T_26182_12_stat_bpd_mispredicted;
  reg [2:0] T_26182_12_fetch_pc_lob;
  reg [19:0] T_26182_12_imm_packed;
  reg [11:0] T_26182_12_csr_addr;
  reg [5:0] T_26182_12_rob_idx;
  reg [3:0] T_26182_12_ldq_idx;
  reg [3:0] T_26182_12_stq_idx;
  reg [4:0] T_26182_12_brob_idx;
  reg [6:0] T_26182_12_pdst;
  reg [6:0] T_26182_12_pop1;
  reg [6:0] T_26182_12_pop2;
  reg [6:0] T_26182_12_pop3;
  reg  T_26182_12_prs1_busy;
  reg  T_26182_12_prs2_busy;
  reg  T_26182_12_prs3_busy;
  reg [6:0] T_26182_12_stale_pdst;
  reg  T_26182_12_exception;
  reg [63:0] T_26182_12_exc_cause;
  reg  T_26182_12_bypassable;
  reg [3:0] T_26182_12_mem_cmd;
  reg [2:0] T_26182_12_mem_typ;
  reg  T_26182_12_is_fence;
  reg  T_26182_12_is_fencei;
  reg  T_26182_12_is_store;
  reg  T_26182_12_is_amo;
  reg  T_26182_12_is_load;
  reg  T_26182_12_is_unique;
  reg  T_26182_12_flush_on_commit;
  reg [5:0] T_26182_12_ldst;
  reg [5:0] T_26182_12_lrs1;
  reg [5:0] T_26182_12_lrs2;
  reg [5:0] T_26182_12_lrs3;
  reg  T_26182_12_ldst_val;
  reg [1:0] T_26182_12_dst_rtype;
  reg [1:0] T_26182_12_lrs1_rtype;
  reg [1:0] T_26182_12_lrs2_rtype;
  reg  T_26182_12_frs3_en;
  reg  T_26182_12_fp_val;
  reg  T_26182_12_fp_single;
  reg  T_26182_12_xcpt_if;
  reg  T_26182_12_replay_if;
  reg [63:0] T_26182_12_debug_wdata;
  reg [31:0] T_26182_12_debug_events_fetch_seq;
  reg  T_26182_13_valid;
  reg [1:0] T_26182_13_iw_state;
  reg [8:0] T_26182_13_uopc;
  reg [31:0] T_26182_13_inst;
  reg [39:0] T_26182_13_pc;
  reg [7:0] T_26182_13_fu_code;
  reg [3:0] T_26182_13_ctrl_br_type;
  reg [1:0] T_26182_13_ctrl_op1_sel;
  reg [2:0] T_26182_13_ctrl_op2_sel;
  reg [2:0] T_26182_13_ctrl_imm_sel;
  reg [3:0] T_26182_13_ctrl_op_fcn;
  reg  T_26182_13_ctrl_fcn_dw;
  reg  T_26182_13_ctrl_rf_wen;
  reg [2:0] T_26182_13_ctrl_csr_cmd;
  reg  T_26182_13_ctrl_is_load;
  reg  T_26182_13_ctrl_is_sta;
  reg  T_26182_13_ctrl_is_std;
  reg [1:0] T_26182_13_wakeup_delay;
  reg  T_26182_13_allocate_brtag;
  reg  T_26182_13_is_br_or_jmp;
  reg  T_26182_13_is_jump;
  reg  T_26182_13_is_jal;
  reg  T_26182_13_is_ret;
  reg  T_26182_13_is_call;
  reg [7:0] T_26182_13_br_mask;
  reg [2:0] T_26182_13_br_tag;
  reg  T_26182_13_br_prediction_bpd_predict_val;
  reg  T_26182_13_br_prediction_bpd_predict_taken;
  reg  T_26182_13_br_prediction_btb_hit;
  reg  T_26182_13_br_prediction_btb_predicted;
  reg  T_26182_13_br_prediction_is_br_or_jalr;
  reg  T_26182_13_stat_brjmp_mispredicted;
  reg  T_26182_13_stat_btb_made_pred;
  reg  T_26182_13_stat_btb_mispredicted;
  reg  T_26182_13_stat_bpd_made_pred;
  reg  T_26182_13_stat_bpd_mispredicted;
  reg [2:0] T_26182_13_fetch_pc_lob;
  reg [19:0] T_26182_13_imm_packed;
  reg [11:0] T_26182_13_csr_addr;
  reg [5:0] T_26182_13_rob_idx;
  reg [3:0] T_26182_13_ldq_idx;
  reg [3:0] T_26182_13_stq_idx;
  reg [4:0] T_26182_13_brob_idx;
  reg [6:0] T_26182_13_pdst;
  reg [6:0] T_26182_13_pop1;
  reg [6:0] T_26182_13_pop2;
  reg [6:0] T_26182_13_pop3;
  reg  T_26182_13_prs1_busy;
  reg  T_26182_13_prs2_busy;
  reg  T_26182_13_prs3_busy;
  reg [6:0] T_26182_13_stale_pdst;
  reg  T_26182_13_exception;
  reg [63:0] T_26182_13_exc_cause;
  reg  T_26182_13_bypassable;
  reg [3:0] T_26182_13_mem_cmd;
  reg [2:0] T_26182_13_mem_typ;
  reg  T_26182_13_is_fence;
  reg  T_26182_13_is_fencei;
  reg  T_26182_13_is_store;
  reg  T_26182_13_is_amo;
  reg  T_26182_13_is_load;
  reg  T_26182_13_is_unique;
  reg  T_26182_13_flush_on_commit;
  reg [5:0] T_26182_13_ldst;
  reg [5:0] T_26182_13_lrs1;
  reg [5:0] T_26182_13_lrs2;
  reg [5:0] T_26182_13_lrs3;
  reg  T_26182_13_ldst_val;
  reg [1:0] T_26182_13_dst_rtype;
  reg [1:0] T_26182_13_lrs1_rtype;
  reg [1:0] T_26182_13_lrs2_rtype;
  reg  T_26182_13_frs3_en;
  reg  T_26182_13_fp_val;
  reg  T_26182_13_fp_single;
  reg  T_26182_13_xcpt_if;
  reg  T_26182_13_replay_if;
  reg [63:0] T_26182_13_debug_wdata;
  reg [31:0] T_26182_13_debug_events_fetch_seq;
  reg  T_26182_14_valid;
  reg [1:0] T_26182_14_iw_state;
  reg [8:0] T_26182_14_uopc;
  reg [31:0] T_26182_14_inst;
  reg [39:0] T_26182_14_pc;
  reg [7:0] T_26182_14_fu_code;
  reg [3:0] T_26182_14_ctrl_br_type;
  reg [1:0] T_26182_14_ctrl_op1_sel;
  reg [2:0] T_26182_14_ctrl_op2_sel;
  reg [2:0] T_26182_14_ctrl_imm_sel;
  reg [3:0] T_26182_14_ctrl_op_fcn;
  reg  T_26182_14_ctrl_fcn_dw;
  reg  T_26182_14_ctrl_rf_wen;
  reg [2:0] T_26182_14_ctrl_csr_cmd;
  reg  T_26182_14_ctrl_is_load;
  reg  T_26182_14_ctrl_is_sta;
  reg  T_26182_14_ctrl_is_std;
  reg [1:0] T_26182_14_wakeup_delay;
  reg  T_26182_14_allocate_brtag;
  reg  T_26182_14_is_br_or_jmp;
  reg  T_26182_14_is_jump;
  reg  T_26182_14_is_jal;
  reg  T_26182_14_is_ret;
  reg  T_26182_14_is_call;
  reg [7:0] T_26182_14_br_mask;
  reg [2:0] T_26182_14_br_tag;
  reg  T_26182_14_br_prediction_bpd_predict_val;
  reg  T_26182_14_br_prediction_bpd_predict_taken;
  reg  T_26182_14_br_prediction_btb_hit;
  reg  T_26182_14_br_prediction_btb_predicted;
  reg  T_26182_14_br_prediction_is_br_or_jalr;
  reg  T_26182_14_stat_brjmp_mispredicted;
  reg  T_26182_14_stat_btb_made_pred;
  reg  T_26182_14_stat_btb_mispredicted;
  reg  T_26182_14_stat_bpd_made_pred;
  reg  T_26182_14_stat_bpd_mispredicted;
  reg [2:0] T_26182_14_fetch_pc_lob;
  reg [19:0] T_26182_14_imm_packed;
  reg [11:0] T_26182_14_csr_addr;
  reg [5:0] T_26182_14_rob_idx;
  reg [3:0] T_26182_14_ldq_idx;
  reg [3:0] T_26182_14_stq_idx;
  reg [4:0] T_26182_14_brob_idx;
  reg [6:0] T_26182_14_pdst;
  reg [6:0] T_26182_14_pop1;
  reg [6:0] T_26182_14_pop2;
  reg [6:0] T_26182_14_pop3;
  reg  T_26182_14_prs1_busy;
  reg  T_26182_14_prs2_busy;
  reg  T_26182_14_prs3_busy;
  reg [6:0] T_26182_14_stale_pdst;
  reg  T_26182_14_exception;
  reg [63:0] T_26182_14_exc_cause;
  reg  T_26182_14_bypassable;
  reg [3:0] T_26182_14_mem_cmd;
  reg [2:0] T_26182_14_mem_typ;
  reg  T_26182_14_is_fence;
  reg  T_26182_14_is_fencei;
  reg  T_26182_14_is_store;
  reg  T_26182_14_is_amo;
  reg  T_26182_14_is_load;
  reg  T_26182_14_is_unique;
  reg  T_26182_14_flush_on_commit;
  reg [5:0] T_26182_14_ldst;
  reg [5:0] T_26182_14_lrs1;
  reg [5:0] T_26182_14_lrs2;
  reg [5:0] T_26182_14_lrs3;
  reg  T_26182_14_ldst_val;
  reg [1:0] T_26182_14_dst_rtype;
  reg [1:0] T_26182_14_lrs1_rtype;
  reg [1:0] T_26182_14_lrs2_rtype;
  reg  T_26182_14_frs3_en;
  reg  T_26182_14_fp_val;
  reg  T_26182_14_fp_single;
  reg  T_26182_14_xcpt_if;
  reg  T_26182_14_replay_if;
  reg [63:0] T_26182_14_debug_wdata;
  reg [31:0] T_26182_14_debug_events_fetch_seq;
  reg  T_26182_15_valid;
  reg [1:0] T_26182_15_iw_state;
  reg [8:0] T_26182_15_uopc;
  reg [31:0] T_26182_15_inst;
  reg [39:0] T_26182_15_pc;
  reg [7:0] T_26182_15_fu_code;
  reg [3:0] T_26182_15_ctrl_br_type;
  reg [1:0] T_26182_15_ctrl_op1_sel;
  reg [2:0] T_26182_15_ctrl_op2_sel;
  reg [2:0] T_26182_15_ctrl_imm_sel;
  reg [3:0] T_26182_15_ctrl_op_fcn;
  reg  T_26182_15_ctrl_fcn_dw;
  reg  T_26182_15_ctrl_rf_wen;
  reg [2:0] T_26182_15_ctrl_csr_cmd;
  reg  T_26182_15_ctrl_is_load;
  reg  T_26182_15_ctrl_is_sta;
  reg  T_26182_15_ctrl_is_std;
  reg [1:0] T_26182_15_wakeup_delay;
  reg  T_26182_15_allocate_brtag;
  reg  T_26182_15_is_br_or_jmp;
  reg  T_26182_15_is_jump;
  reg  T_26182_15_is_jal;
  reg  T_26182_15_is_ret;
  reg  T_26182_15_is_call;
  reg [7:0] T_26182_15_br_mask;
  reg [2:0] T_26182_15_br_tag;
  reg  T_26182_15_br_prediction_bpd_predict_val;
  reg  T_26182_15_br_prediction_bpd_predict_taken;
  reg  T_26182_15_br_prediction_btb_hit;
  reg  T_26182_15_br_prediction_btb_predicted;
  reg  T_26182_15_br_prediction_is_br_or_jalr;
  reg  T_26182_15_stat_brjmp_mispredicted;
  reg  T_26182_15_stat_btb_made_pred;
  reg  T_26182_15_stat_btb_mispredicted;
  reg  T_26182_15_stat_bpd_made_pred;
  reg  T_26182_15_stat_bpd_mispredicted;
  reg [2:0] T_26182_15_fetch_pc_lob;
  reg [19:0] T_26182_15_imm_packed;
  reg [11:0] T_26182_15_csr_addr;
  reg [5:0] T_26182_15_rob_idx;
  reg [3:0] T_26182_15_ldq_idx;
  reg [3:0] T_26182_15_stq_idx;
  reg [4:0] T_26182_15_brob_idx;
  reg [6:0] T_26182_15_pdst;
  reg [6:0] T_26182_15_pop1;
  reg [6:0] T_26182_15_pop2;
  reg [6:0] T_26182_15_pop3;
  reg  T_26182_15_prs1_busy;
  reg  T_26182_15_prs2_busy;
  reg  T_26182_15_prs3_busy;
  reg [6:0] T_26182_15_stale_pdst;
  reg  T_26182_15_exception;
  reg [63:0] T_26182_15_exc_cause;
  reg  T_26182_15_bypassable;
  reg [3:0] T_26182_15_mem_cmd;
  reg [2:0] T_26182_15_mem_typ;
  reg  T_26182_15_is_fence;
  reg  T_26182_15_is_fencei;
  reg  T_26182_15_is_store;
  reg  T_26182_15_is_amo;
  reg  T_26182_15_is_load;
  reg  T_26182_15_is_unique;
  reg  T_26182_15_flush_on_commit;
  reg [5:0] T_26182_15_ldst;
  reg [5:0] T_26182_15_lrs1;
  reg [5:0] T_26182_15_lrs2;
  reg [5:0] T_26182_15_lrs3;
  reg  T_26182_15_ldst_val;
  reg [1:0] T_26182_15_dst_rtype;
  reg [1:0] T_26182_15_lrs1_rtype;
  reg [1:0] T_26182_15_lrs2_rtype;
  reg  T_26182_15_frs3_en;
  reg  T_26182_15_fp_val;
  reg  T_26182_15_fp_single;
  reg  T_26182_15_xcpt_if;
  reg  T_26182_15_replay_if;
  reg [63:0] T_26182_15_debug_wdata;
  reg [31:0] T_26182_15_debug_events_fetch_seq;
  reg  T_26182_16_valid;
  reg [1:0] T_26182_16_iw_state;
  reg [8:0] T_26182_16_uopc;
  reg [31:0] T_26182_16_inst;
  reg [39:0] T_26182_16_pc;
  reg [7:0] T_26182_16_fu_code;
  reg [3:0] T_26182_16_ctrl_br_type;
  reg [1:0] T_26182_16_ctrl_op1_sel;
  reg [2:0] T_26182_16_ctrl_op2_sel;
  reg [2:0] T_26182_16_ctrl_imm_sel;
  reg [3:0] T_26182_16_ctrl_op_fcn;
  reg  T_26182_16_ctrl_fcn_dw;
  reg  T_26182_16_ctrl_rf_wen;
  reg [2:0] T_26182_16_ctrl_csr_cmd;
  reg  T_26182_16_ctrl_is_load;
  reg  T_26182_16_ctrl_is_sta;
  reg  T_26182_16_ctrl_is_std;
  reg [1:0] T_26182_16_wakeup_delay;
  reg  T_26182_16_allocate_brtag;
  reg  T_26182_16_is_br_or_jmp;
  reg  T_26182_16_is_jump;
  reg  T_26182_16_is_jal;
  reg  T_26182_16_is_ret;
  reg  T_26182_16_is_call;
  reg [7:0] T_26182_16_br_mask;
  reg [2:0] T_26182_16_br_tag;
  reg  T_26182_16_br_prediction_bpd_predict_val;
  reg  T_26182_16_br_prediction_bpd_predict_taken;
  reg  T_26182_16_br_prediction_btb_hit;
  reg  T_26182_16_br_prediction_btb_predicted;
  reg  T_26182_16_br_prediction_is_br_or_jalr;
  reg  T_26182_16_stat_brjmp_mispredicted;
  reg  T_26182_16_stat_btb_made_pred;
  reg  T_26182_16_stat_btb_mispredicted;
  reg  T_26182_16_stat_bpd_made_pred;
  reg  T_26182_16_stat_bpd_mispredicted;
  reg [2:0] T_26182_16_fetch_pc_lob;
  reg [19:0] T_26182_16_imm_packed;
  reg [11:0] T_26182_16_csr_addr;
  reg [5:0] T_26182_16_rob_idx;
  reg [3:0] T_26182_16_ldq_idx;
  reg [3:0] T_26182_16_stq_idx;
  reg [4:0] T_26182_16_brob_idx;
  reg [6:0] T_26182_16_pdst;
  reg [6:0] T_26182_16_pop1;
  reg [6:0] T_26182_16_pop2;
  reg [6:0] T_26182_16_pop3;
  reg  T_26182_16_prs1_busy;
  reg  T_26182_16_prs2_busy;
  reg  T_26182_16_prs3_busy;
  reg [6:0] T_26182_16_stale_pdst;
  reg  T_26182_16_exception;
  reg [63:0] T_26182_16_exc_cause;
  reg  T_26182_16_bypassable;
  reg [3:0] T_26182_16_mem_cmd;
  reg [2:0] T_26182_16_mem_typ;
  reg  T_26182_16_is_fence;
  reg  T_26182_16_is_fencei;
  reg  T_26182_16_is_store;
  reg  T_26182_16_is_amo;
  reg  T_26182_16_is_load;
  reg  T_26182_16_is_unique;
  reg  T_26182_16_flush_on_commit;
  reg [5:0] T_26182_16_ldst;
  reg [5:0] T_26182_16_lrs1;
  reg [5:0] T_26182_16_lrs2;
  reg [5:0] T_26182_16_lrs3;
  reg  T_26182_16_ldst_val;
  reg [1:0] T_26182_16_dst_rtype;
  reg [1:0] T_26182_16_lrs1_rtype;
  reg [1:0] T_26182_16_lrs2_rtype;
  reg  T_26182_16_frs3_en;
  reg  T_26182_16_fp_val;
  reg  T_26182_16_fp_single;
  reg  T_26182_16_xcpt_if;
  reg  T_26182_16_replay_if;
  reg [63:0] T_26182_16_debug_wdata;
  reg [31:0] T_26182_16_debug_events_fetch_seq;
  reg  T_26182_17_valid;
  reg [1:0] T_26182_17_iw_state;
  reg [8:0] T_26182_17_uopc;
  reg [31:0] T_26182_17_inst;
  reg [39:0] T_26182_17_pc;
  reg [7:0] T_26182_17_fu_code;
  reg [3:0] T_26182_17_ctrl_br_type;
  reg [1:0] T_26182_17_ctrl_op1_sel;
  reg [2:0] T_26182_17_ctrl_op2_sel;
  reg [2:0] T_26182_17_ctrl_imm_sel;
  reg [3:0] T_26182_17_ctrl_op_fcn;
  reg  T_26182_17_ctrl_fcn_dw;
  reg  T_26182_17_ctrl_rf_wen;
  reg [2:0] T_26182_17_ctrl_csr_cmd;
  reg  T_26182_17_ctrl_is_load;
  reg  T_26182_17_ctrl_is_sta;
  reg  T_26182_17_ctrl_is_std;
  reg [1:0] T_26182_17_wakeup_delay;
  reg  T_26182_17_allocate_brtag;
  reg  T_26182_17_is_br_or_jmp;
  reg  T_26182_17_is_jump;
  reg  T_26182_17_is_jal;
  reg  T_26182_17_is_ret;
  reg  T_26182_17_is_call;
  reg [7:0] T_26182_17_br_mask;
  reg [2:0] T_26182_17_br_tag;
  reg  T_26182_17_br_prediction_bpd_predict_val;
  reg  T_26182_17_br_prediction_bpd_predict_taken;
  reg  T_26182_17_br_prediction_btb_hit;
  reg  T_26182_17_br_prediction_btb_predicted;
  reg  T_26182_17_br_prediction_is_br_or_jalr;
  reg  T_26182_17_stat_brjmp_mispredicted;
  reg  T_26182_17_stat_btb_made_pred;
  reg  T_26182_17_stat_btb_mispredicted;
  reg  T_26182_17_stat_bpd_made_pred;
  reg  T_26182_17_stat_bpd_mispredicted;
  reg [2:0] T_26182_17_fetch_pc_lob;
  reg [19:0] T_26182_17_imm_packed;
  reg [11:0] T_26182_17_csr_addr;
  reg [5:0] T_26182_17_rob_idx;
  reg [3:0] T_26182_17_ldq_idx;
  reg [3:0] T_26182_17_stq_idx;
  reg [4:0] T_26182_17_brob_idx;
  reg [6:0] T_26182_17_pdst;
  reg [6:0] T_26182_17_pop1;
  reg [6:0] T_26182_17_pop2;
  reg [6:0] T_26182_17_pop3;
  reg  T_26182_17_prs1_busy;
  reg  T_26182_17_prs2_busy;
  reg  T_26182_17_prs3_busy;
  reg [6:0] T_26182_17_stale_pdst;
  reg  T_26182_17_exception;
  reg [63:0] T_26182_17_exc_cause;
  reg  T_26182_17_bypassable;
  reg [3:0] T_26182_17_mem_cmd;
  reg [2:0] T_26182_17_mem_typ;
  reg  T_26182_17_is_fence;
  reg  T_26182_17_is_fencei;
  reg  T_26182_17_is_store;
  reg  T_26182_17_is_amo;
  reg  T_26182_17_is_load;
  reg  T_26182_17_is_unique;
  reg  T_26182_17_flush_on_commit;
  reg [5:0] T_26182_17_ldst;
  reg [5:0] T_26182_17_lrs1;
  reg [5:0] T_26182_17_lrs2;
  reg [5:0] T_26182_17_lrs3;
  reg  T_26182_17_ldst_val;
  reg [1:0] T_26182_17_dst_rtype;
  reg [1:0] T_26182_17_lrs1_rtype;
  reg [1:0] T_26182_17_lrs2_rtype;
  reg  T_26182_17_frs3_en;
  reg  T_26182_17_fp_val;
  reg  T_26182_17_fp_single;
  reg  T_26182_17_xcpt_if;
  reg  T_26182_17_replay_if;
  reg [63:0] T_26182_17_debug_wdata;
  reg [31:0] T_26182_17_debug_events_fetch_seq;
  reg  T_26182_18_valid;
  reg [1:0] T_26182_18_iw_state;
  reg [8:0] T_26182_18_uopc;
  reg [31:0] T_26182_18_inst;
  reg [39:0] T_26182_18_pc;
  reg [7:0] T_26182_18_fu_code;
  reg [3:0] T_26182_18_ctrl_br_type;
  reg [1:0] T_26182_18_ctrl_op1_sel;
  reg [2:0] T_26182_18_ctrl_op2_sel;
  reg [2:0] T_26182_18_ctrl_imm_sel;
  reg [3:0] T_26182_18_ctrl_op_fcn;
  reg  T_26182_18_ctrl_fcn_dw;
  reg  T_26182_18_ctrl_rf_wen;
  reg [2:0] T_26182_18_ctrl_csr_cmd;
  reg  T_26182_18_ctrl_is_load;
  reg  T_26182_18_ctrl_is_sta;
  reg  T_26182_18_ctrl_is_std;
  reg [1:0] T_26182_18_wakeup_delay;
  reg  T_26182_18_allocate_brtag;
  reg  T_26182_18_is_br_or_jmp;
  reg  T_26182_18_is_jump;
  reg  T_26182_18_is_jal;
  reg  T_26182_18_is_ret;
  reg  T_26182_18_is_call;
  reg [7:0] T_26182_18_br_mask;
  reg [2:0] T_26182_18_br_tag;
  reg  T_26182_18_br_prediction_bpd_predict_val;
  reg  T_26182_18_br_prediction_bpd_predict_taken;
  reg  T_26182_18_br_prediction_btb_hit;
  reg  T_26182_18_br_prediction_btb_predicted;
  reg  T_26182_18_br_prediction_is_br_or_jalr;
  reg  T_26182_18_stat_brjmp_mispredicted;
  reg  T_26182_18_stat_btb_made_pred;
  reg  T_26182_18_stat_btb_mispredicted;
  reg  T_26182_18_stat_bpd_made_pred;
  reg  T_26182_18_stat_bpd_mispredicted;
  reg [2:0] T_26182_18_fetch_pc_lob;
  reg [19:0] T_26182_18_imm_packed;
  reg [11:0] T_26182_18_csr_addr;
  reg [5:0] T_26182_18_rob_idx;
  reg [3:0] T_26182_18_ldq_idx;
  reg [3:0] T_26182_18_stq_idx;
  reg [4:0] T_26182_18_brob_idx;
  reg [6:0] T_26182_18_pdst;
  reg [6:0] T_26182_18_pop1;
  reg [6:0] T_26182_18_pop2;
  reg [6:0] T_26182_18_pop3;
  reg  T_26182_18_prs1_busy;
  reg  T_26182_18_prs2_busy;
  reg  T_26182_18_prs3_busy;
  reg [6:0] T_26182_18_stale_pdst;
  reg  T_26182_18_exception;
  reg [63:0] T_26182_18_exc_cause;
  reg  T_26182_18_bypassable;
  reg [3:0] T_26182_18_mem_cmd;
  reg [2:0] T_26182_18_mem_typ;
  reg  T_26182_18_is_fence;
  reg  T_26182_18_is_fencei;
  reg  T_26182_18_is_store;
  reg  T_26182_18_is_amo;
  reg  T_26182_18_is_load;
  reg  T_26182_18_is_unique;
  reg  T_26182_18_flush_on_commit;
  reg [5:0] T_26182_18_ldst;
  reg [5:0] T_26182_18_lrs1;
  reg [5:0] T_26182_18_lrs2;
  reg [5:0] T_26182_18_lrs3;
  reg  T_26182_18_ldst_val;
  reg [1:0] T_26182_18_dst_rtype;
  reg [1:0] T_26182_18_lrs1_rtype;
  reg [1:0] T_26182_18_lrs2_rtype;
  reg  T_26182_18_frs3_en;
  reg  T_26182_18_fp_val;
  reg  T_26182_18_fp_single;
  reg  T_26182_18_xcpt_if;
  reg  T_26182_18_replay_if;
  reg [63:0] T_26182_18_debug_wdata;
  reg [31:0] T_26182_18_debug_events_fetch_seq;
  reg  T_26182_19_valid;
  reg [1:0] T_26182_19_iw_state;
  reg [8:0] T_26182_19_uopc;
  reg [31:0] T_26182_19_inst;
  reg [39:0] T_26182_19_pc;
  reg [7:0] T_26182_19_fu_code;
  reg [3:0] T_26182_19_ctrl_br_type;
  reg [1:0] T_26182_19_ctrl_op1_sel;
  reg [2:0] T_26182_19_ctrl_op2_sel;
  reg [2:0] T_26182_19_ctrl_imm_sel;
  reg [3:0] T_26182_19_ctrl_op_fcn;
  reg  T_26182_19_ctrl_fcn_dw;
  reg  T_26182_19_ctrl_rf_wen;
  reg [2:0] T_26182_19_ctrl_csr_cmd;
  reg  T_26182_19_ctrl_is_load;
  reg  T_26182_19_ctrl_is_sta;
  reg  T_26182_19_ctrl_is_std;
  reg [1:0] T_26182_19_wakeup_delay;
  reg  T_26182_19_allocate_brtag;
  reg  T_26182_19_is_br_or_jmp;
  reg  T_26182_19_is_jump;
  reg  T_26182_19_is_jal;
  reg  T_26182_19_is_ret;
  reg  T_26182_19_is_call;
  reg [7:0] T_26182_19_br_mask;
  reg [2:0] T_26182_19_br_tag;
  reg  T_26182_19_br_prediction_bpd_predict_val;
  reg  T_26182_19_br_prediction_bpd_predict_taken;
  reg  T_26182_19_br_prediction_btb_hit;
  reg  T_26182_19_br_prediction_btb_predicted;
  reg  T_26182_19_br_prediction_is_br_or_jalr;
  reg  T_26182_19_stat_brjmp_mispredicted;
  reg  T_26182_19_stat_btb_made_pred;
  reg  T_26182_19_stat_btb_mispredicted;
  reg  T_26182_19_stat_bpd_made_pred;
  reg  T_26182_19_stat_bpd_mispredicted;
  reg [2:0] T_26182_19_fetch_pc_lob;
  reg [19:0] T_26182_19_imm_packed;
  reg [11:0] T_26182_19_csr_addr;
  reg [5:0] T_26182_19_rob_idx;
  reg [3:0] T_26182_19_ldq_idx;
  reg [3:0] T_26182_19_stq_idx;
  reg [4:0] T_26182_19_brob_idx;
  reg [6:0] T_26182_19_pdst;
  reg [6:0] T_26182_19_pop1;
  reg [6:0] T_26182_19_pop2;
  reg [6:0] T_26182_19_pop3;
  reg  T_26182_19_prs1_busy;
  reg  T_26182_19_prs2_busy;
  reg  T_26182_19_prs3_busy;
  reg [6:0] T_26182_19_stale_pdst;
  reg  T_26182_19_exception;
  reg [63:0] T_26182_19_exc_cause;
  reg  T_26182_19_bypassable;
  reg [3:0] T_26182_19_mem_cmd;
  reg [2:0] T_26182_19_mem_typ;
  reg  T_26182_19_is_fence;
  reg  T_26182_19_is_fencei;
  reg  T_26182_19_is_store;
  reg  T_26182_19_is_amo;
  reg  T_26182_19_is_load;
  reg  T_26182_19_is_unique;
  reg  T_26182_19_flush_on_commit;
  reg [5:0] T_26182_19_ldst;
  reg [5:0] T_26182_19_lrs1;
  reg [5:0] T_26182_19_lrs2;
  reg [5:0] T_26182_19_lrs3;
  reg  T_26182_19_ldst_val;
  reg [1:0] T_26182_19_dst_rtype;
  reg [1:0] T_26182_19_lrs1_rtype;
  reg [1:0] T_26182_19_lrs2_rtype;
  reg  T_26182_19_frs3_en;
  reg  T_26182_19_fp_val;
  reg  T_26182_19_fp_single;
  reg  T_26182_19_xcpt_if;
  reg  T_26182_19_replay_if;
  reg [63:0] T_26182_19_debug_wdata;
  reg [31:0] T_26182_19_debug_events_fetch_seq;
  reg  T_26182_20_valid;
  reg [1:0] T_26182_20_iw_state;
  reg [8:0] T_26182_20_uopc;
  reg [31:0] T_26182_20_inst;
  reg [39:0] T_26182_20_pc;
  reg [7:0] T_26182_20_fu_code;
  reg [3:0] T_26182_20_ctrl_br_type;
  reg [1:0] T_26182_20_ctrl_op1_sel;
  reg [2:0] T_26182_20_ctrl_op2_sel;
  reg [2:0] T_26182_20_ctrl_imm_sel;
  reg [3:0] T_26182_20_ctrl_op_fcn;
  reg  T_26182_20_ctrl_fcn_dw;
  reg  T_26182_20_ctrl_rf_wen;
  reg [2:0] T_26182_20_ctrl_csr_cmd;
  reg  T_26182_20_ctrl_is_load;
  reg  T_26182_20_ctrl_is_sta;
  reg  T_26182_20_ctrl_is_std;
  reg [1:0] T_26182_20_wakeup_delay;
  reg  T_26182_20_allocate_brtag;
  reg  T_26182_20_is_br_or_jmp;
  reg  T_26182_20_is_jump;
  reg  T_26182_20_is_jal;
  reg  T_26182_20_is_ret;
  reg  T_26182_20_is_call;
  reg [7:0] T_26182_20_br_mask;
  reg [2:0] T_26182_20_br_tag;
  reg  T_26182_20_br_prediction_bpd_predict_val;
  reg  T_26182_20_br_prediction_bpd_predict_taken;
  reg  T_26182_20_br_prediction_btb_hit;
  reg  T_26182_20_br_prediction_btb_predicted;
  reg  T_26182_20_br_prediction_is_br_or_jalr;
  reg  T_26182_20_stat_brjmp_mispredicted;
  reg  T_26182_20_stat_btb_made_pred;
  reg  T_26182_20_stat_btb_mispredicted;
  reg  T_26182_20_stat_bpd_made_pred;
  reg  T_26182_20_stat_bpd_mispredicted;
  reg [2:0] T_26182_20_fetch_pc_lob;
  reg [19:0] T_26182_20_imm_packed;
  reg [11:0] T_26182_20_csr_addr;
  reg [5:0] T_26182_20_rob_idx;
  reg [3:0] T_26182_20_ldq_idx;
  reg [3:0] T_26182_20_stq_idx;
  reg [4:0] T_26182_20_brob_idx;
  reg [6:0] T_26182_20_pdst;
  reg [6:0] T_26182_20_pop1;
  reg [6:0] T_26182_20_pop2;
  reg [6:0] T_26182_20_pop3;
  reg  T_26182_20_prs1_busy;
  reg  T_26182_20_prs2_busy;
  reg  T_26182_20_prs3_busy;
  reg [6:0] T_26182_20_stale_pdst;
  reg  T_26182_20_exception;
  reg [63:0] T_26182_20_exc_cause;
  reg  T_26182_20_bypassable;
  reg [3:0] T_26182_20_mem_cmd;
  reg [2:0] T_26182_20_mem_typ;
  reg  T_26182_20_is_fence;
  reg  T_26182_20_is_fencei;
  reg  T_26182_20_is_store;
  reg  T_26182_20_is_amo;
  reg  T_26182_20_is_load;
  reg  T_26182_20_is_unique;
  reg  T_26182_20_flush_on_commit;
  reg [5:0] T_26182_20_ldst;
  reg [5:0] T_26182_20_lrs1;
  reg [5:0] T_26182_20_lrs2;
  reg [5:0] T_26182_20_lrs3;
  reg  T_26182_20_ldst_val;
  reg [1:0] T_26182_20_dst_rtype;
  reg [1:0] T_26182_20_lrs1_rtype;
  reg [1:0] T_26182_20_lrs2_rtype;
  reg  T_26182_20_frs3_en;
  reg  T_26182_20_fp_val;
  reg  T_26182_20_fp_single;
  reg  T_26182_20_xcpt_if;
  reg  T_26182_20_replay_if;
  reg [63:0] T_26182_20_debug_wdata;
  reg [31:0] T_26182_20_debug_events_fetch_seq;
  reg  T_26182_21_valid;
  reg [1:0] T_26182_21_iw_state;
  reg [8:0] T_26182_21_uopc;
  reg [31:0] T_26182_21_inst;
  reg [39:0] T_26182_21_pc;
  reg [7:0] T_26182_21_fu_code;
  reg [3:0] T_26182_21_ctrl_br_type;
  reg [1:0] T_26182_21_ctrl_op1_sel;
  reg [2:0] T_26182_21_ctrl_op2_sel;
  reg [2:0] T_26182_21_ctrl_imm_sel;
  reg [3:0] T_26182_21_ctrl_op_fcn;
  reg  T_26182_21_ctrl_fcn_dw;
  reg  T_26182_21_ctrl_rf_wen;
  reg [2:0] T_26182_21_ctrl_csr_cmd;
  reg  T_26182_21_ctrl_is_load;
  reg  T_26182_21_ctrl_is_sta;
  reg  T_26182_21_ctrl_is_std;
  reg [1:0] T_26182_21_wakeup_delay;
  reg  T_26182_21_allocate_brtag;
  reg  T_26182_21_is_br_or_jmp;
  reg  T_26182_21_is_jump;
  reg  T_26182_21_is_jal;
  reg  T_26182_21_is_ret;
  reg  T_26182_21_is_call;
  reg [7:0] T_26182_21_br_mask;
  reg [2:0] T_26182_21_br_tag;
  reg  T_26182_21_br_prediction_bpd_predict_val;
  reg  T_26182_21_br_prediction_bpd_predict_taken;
  reg  T_26182_21_br_prediction_btb_hit;
  reg  T_26182_21_br_prediction_btb_predicted;
  reg  T_26182_21_br_prediction_is_br_or_jalr;
  reg  T_26182_21_stat_brjmp_mispredicted;
  reg  T_26182_21_stat_btb_made_pred;
  reg  T_26182_21_stat_btb_mispredicted;
  reg  T_26182_21_stat_bpd_made_pred;
  reg  T_26182_21_stat_bpd_mispredicted;
  reg [2:0] T_26182_21_fetch_pc_lob;
  reg [19:0] T_26182_21_imm_packed;
  reg [11:0] T_26182_21_csr_addr;
  reg [5:0] T_26182_21_rob_idx;
  reg [3:0] T_26182_21_ldq_idx;
  reg [3:0] T_26182_21_stq_idx;
  reg [4:0] T_26182_21_brob_idx;
  reg [6:0] T_26182_21_pdst;
  reg [6:0] T_26182_21_pop1;
  reg [6:0] T_26182_21_pop2;
  reg [6:0] T_26182_21_pop3;
  reg  T_26182_21_prs1_busy;
  reg  T_26182_21_prs2_busy;
  reg  T_26182_21_prs3_busy;
  reg [6:0] T_26182_21_stale_pdst;
  reg  T_26182_21_exception;
  reg [63:0] T_26182_21_exc_cause;
  reg  T_26182_21_bypassable;
  reg [3:0] T_26182_21_mem_cmd;
  reg [2:0] T_26182_21_mem_typ;
  reg  T_26182_21_is_fence;
  reg  T_26182_21_is_fencei;
  reg  T_26182_21_is_store;
  reg  T_26182_21_is_amo;
  reg  T_26182_21_is_load;
  reg  T_26182_21_is_unique;
  reg  T_26182_21_flush_on_commit;
  reg [5:0] T_26182_21_ldst;
  reg [5:0] T_26182_21_lrs1;
  reg [5:0] T_26182_21_lrs2;
  reg [5:0] T_26182_21_lrs3;
  reg  T_26182_21_ldst_val;
  reg [1:0] T_26182_21_dst_rtype;
  reg [1:0] T_26182_21_lrs1_rtype;
  reg [1:0] T_26182_21_lrs2_rtype;
  reg  T_26182_21_frs3_en;
  reg  T_26182_21_fp_val;
  reg  T_26182_21_fp_single;
  reg  T_26182_21_xcpt_if;
  reg  T_26182_21_replay_if;
  reg [63:0] T_26182_21_debug_wdata;
  reg [31:0] T_26182_21_debug_events_fetch_seq;
  reg  T_26182_22_valid;
  reg [1:0] T_26182_22_iw_state;
  reg [8:0] T_26182_22_uopc;
  reg [31:0] T_26182_22_inst;
  reg [39:0] T_26182_22_pc;
  reg [7:0] T_26182_22_fu_code;
  reg [3:0] T_26182_22_ctrl_br_type;
  reg [1:0] T_26182_22_ctrl_op1_sel;
  reg [2:0] T_26182_22_ctrl_op2_sel;
  reg [2:0] T_26182_22_ctrl_imm_sel;
  reg [3:0] T_26182_22_ctrl_op_fcn;
  reg  T_26182_22_ctrl_fcn_dw;
  reg  T_26182_22_ctrl_rf_wen;
  reg [2:0] T_26182_22_ctrl_csr_cmd;
  reg  T_26182_22_ctrl_is_load;
  reg  T_26182_22_ctrl_is_sta;
  reg  T_26182_22_ctrl_is_std;
  reg [1:0] T_26182_22_wakeup_delay;
  reg  T_26182_22_allocate_brtag;
  reg  T_26182_22_is_br_or_jmp;
  reg  T_26182_22_is_jump;
  reg  T_26182_22_is_jal;
  reg  T_26182_22_is_ret;
  reg  T_26182_22_is_call;
  reg [7:0] T_26182_22_br_mask;
  reg [2:0] T_26182_22_br_tag;
  reg  T_26182_22_br_prediction_bpd_predict_val;
  reg  T_26182_22_br_prediction_bpd_predict_taken;
  reg  T_26182_22_br_prediction_btb_hit;
  reg  T_26182_22_br_prediction_btb_predicted;
  reg  T_26182_22_br_prediction_is_br_or_jalr;
  reg  T_26182_22_stat_brjmp_mispredicted;
  reg  T_26182_22_stat_btb_made_pred;
  reg  T_26182_22_stat_btb_mispredicted;
  reg  T_26182_22_stat_bpd_made_pred;
  reg  T_26182_22_stat_bpd_mispredicted;
  reg [2:0] T_26182_22_fetch_pc_lob;
  reg [19:0] T_26182_22_imm_packed;
  reg [11:0] T_26182_22_csr_addr;
  reg [5:0] T_26182_22_rob_idx;
  reg [3:0] T_26182_22_ldq_idx;
  reg [3:0] T_26182_22_stq_idx;
  reg [4:0] T_26182_22_brob_idx;
  reg [6:0] T_26182_22_pdst;
  reg [6:0] T_26182_22_pop1;
  reg [6:0] T_26182_22_pop2;
  reg [6:0] T_26182_22_pop3;
  reg  T_26182_22_prs1_busy;
  reg  T_26182_22_prs2_busy;
  reg  T_26182_22_prs3_busy;
  reg [6:0] T_26182_22_stale_pdst;
  reg  T_26182_22_exception;
  reg [63:0] T_26182_22_exc_cause;
  reg  T_26182_22_bypassable;
  reg [3:0] T_26182_22_mem_cmd;
  reg [2:0] T_26182_22_mem_typ;
  reg  T_26182_22_is_fence;
  reg  T_26182_22_is_fencei;
  reg  T_26182_22_is_store;
  reg  T_26182_22_is_amo;
  reg  T_26182_22_is_load;
  reg  T_26182_22_is_unique;
  reg  T_26182_22_flush_on_commit;
  reg [5:0] T_26182_22_ldst;
  reg [5:0] T_26182_22_lrs1;
  reg [5:0] T_26182_22_lrs2;
  reg [5:0] T_26182_22_lrs3;
  reg  T_26182_22_ldst_val;
  reg [1:0] T_26182_22_dst_rtype;
  reg [1:0] T_26182_22_lrs1_rtype;
  reg [1:0] T_26182_22_lrs2_rtype;
  reg  T_26182_22_frs3_en;
  reg  T_26182_22_fp_val;
  reg  T_26182_22_fp_single;
  reg  T_26182_22_xcpt_if;
  reg  T_26182_22_replay_if;
  reg [63:0] T_26182_22_debug_wdata;
  reg [31:0] T_26182_22_debug_events_fetch_seq;
  reg  T_26182_23_valid;
  reg [1:0] T_26182_23_iw_state;
  reg [8:0] T_26182_23_uopc;
  reg [31:0] T_26182_23_inst;
  reg [39:0] T_26182_23_pc;
  reg [7:0] T_26182_23_fu_code;
  reg [3:0] T_26182_23_ctrl_br_type;
  reg [1:0] T_26182_23_ctrl_op1_sel;
  reg [2:0] T_26182_23_ctrl_op2_sel;
  reg [2:0] T_26182_23_ctrl_imm_sel;
  reg [3:0] T_26182_23_ctrl_op_fcn;
  reg  T_26182_23_ctrl_fcn_dw;
  reg  T_26182_23_ctrl_rf_wen;
  reg [2:0] T_26182_23_ctrl_csr_cmd;
  reg  T_26182_23_ctrl_is_load;
  reg  T_26182_23_ctrl_is_sta;
  reg  T_26182_23_ctrl_is_std;
  reg [1:0] T_26182_23_wakeup_delay;
  reg  T_26182_23_allocate_brtag;
  reg  T_26182_23_is_br_or_jmp;
  reg  T_26182_23_is_jump;
  reg  T_26182_23_is_jal;
  reg  T_26182_23_is_ret;
  reg  T_26182_23_is_call;
  reg [7:0] T_26182_23_br_mask;
  reg [2:0] T_26182_23_br_tag;
  reg  T_26182_23_br_prediction_bpd_predict_val;
  reg  T_26182_23_br_prediction_bpd_predict_taken;
  reg  T_26182_23_br_prediction_btb_hit;
  reg  T_26182_23_br_prediction_btb_predicted;
  reg  T_26182_23_br_prediction_is_br_or_jalr;
  reg  T_26182_23_stat_brjmp_mispredicted;
  reg  T_26182_23_stat_btb_made_pred;
  reg  T_26182_23_stat_btb_mispredicted;
  reg  T_26182_23_stat_bpd_made_pred;
  reg  T_26182_23_stat_bpd_mispredicted;
  reg [2:0] T_26182_23_fetch_pc_lob;
  reg [19:0] T_26182_23_imm_packed;
  reg [11:0] T_26182_23_csr_addr;
  reg [5:0] T_26182_23_rob_idx;
  reg [3:0] T_26182_23_ldq_idx;
  reg [3:0] T_26182_23_stq_idx;
  reg [4:0] T_26182_23_brob_idx;
  reg [6:0] T_26182_23_pdst;
  reg [6:0] T_26182_23_pop1;
  reg [6:0] T_26182_23_pop2;
  reg [6:0] T_26182_23_pop3;
  reg  T_26182_23_prs1_busy;
  reg  T_26182_23_prs2_busy;
  reg  T_26182_23_prs3_busy;
  reg [6:0] T_26182_23_stale_pdst;
  reg  T_26182_23_exception;
  reg [63:0] T_26182_23_exc_cause;
  reg  T_26182_23_bypassable;
  reg [3:0] T_26182_23_mem_cmd;
  reg [2:0] T_26182_23_mem_typ;
  reg  T_26182_23_is_fence;
  reg  T_26182_23_is_fencei;
  reg  T_26182_23_is_store;
  reg  T_26182_23_is_amo;
  reg  T_26182_23_is_load;
  reg  T_26182_23_is_unique;
  reg  T_26182_23_flush_on_commit;
  reg [5:0] T_26182_23_ldst;
  reg [5:0] T_26182_23_lrs1;
  reg [5:0] T_26182_23_lrs2;
  reg [5:0] T_26182_23_lrs3;
  reg  T_26182_23_ldst_val;
  reg [1:0] T_26182_23_dst_rtype;
  reg [1:0] T_26182_23_lrs1_rtype;
  reg [1:0] T_26182_23_lrs2_rtype;
  reg  T_26182_23_frs3_en;
  reg  T_26182_23_fp_val;
  reg  T_26182_23_fp_single;
  reg  T_26182_23_xcpt_if;
  reg  T_26182_23_replay_if;
  reg [63:0] T_26182_23_debug_wdata;
  reg [31:0] T_26182_23_debug_events_fetch_seq;
  wire  _GEN_33 = 5'h0 == rob_tail | T_23706_0; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_34 = 5'h1 == rob_tail | T_23706_1; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_35 = 5'h2 == rob_tail | T_23706_2; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_36 = 5'h3 == rob_tail | T_23706_3; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_37 = 5'h4 == rob_tail | T_23706_4; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_38 = 5'h5 == rob_tail | T_23706_5; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_39 = 5'h6 == rob_tail | T_23706_6; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_40 = 5'h7 == rob_tail | T_23706_7; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_41 = 5'h8 == rob_tail | T_23706_8; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_42 = 5'h9 == rob_tail | T_23706_9; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_43 = 5'ha == rob_tail | T_23706_10; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_44 = 5'hb == rob_tail | T_23706_11; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_45 = 5'hc == rob_tail | T_23706_12; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_46 = 5'hd == rob_tail | T_23706_13; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_47 = 5'he == rob_tail | T_23706_14; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_48 = 5'hf == rob_tail | T_23706_15; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_49 = 5'h10 == rob_tail | T_23706_16; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_50 = 5'h11 == rob_tail | T_23706_17; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_51 = 5'h12 == rob_tail | T_23706_18; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_52 = 5'h13 == rob_tail | T_23706_19; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_53 = 5'h14 == rob_tail | T_23706_20; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_54 = 5'h15 == rob_tail | T_23706_21; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_55 = 5'h16 == rob_tail | T_23706_22; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_56 = 5'h17 == rob_tail | T_23706_23; // @[rob.scala 347:34 rob.scala 347:34]
  wire [31:0] _GEN_129 = 5'h0 == rob_tail ? io_dis_uops_0_inst : T_26182_0_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_130 = 5'h1 == rob_tail ? io_dis_uops_0_inst : T_26182_1_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_131 = 5'h2 == rob_tail ? io_dis_uops_0_inst : T_26182_2_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_132 = 5'h3 == rob_tail ? io_dis_uops_0_inst : T_26182_3_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_133 = 5'h4 == rob_tail ? io_dis_uops_0_inst : T_26182_4_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_134 = 5'h5 == rob_tail ? io_dis_uops_0_inst : T_26182_5_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_135 = 5'h6 == rob_tail ? io_dis_uops_0_inst : T_26182_6_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_136 = 5'h7 == rob_tail ? io_dis_uops_0_inst : T_26182_7_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_137 = 5'h8 == rob_tail ? io_dis_uops_0_inst : T_26182_8_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_138 = 5'h9 == rob_tail ? io_dis_uops_0_inst : T_26182_9_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_139 = 5'ha == rob_tail ? io_dis_uops_0_inst : T_26182_10_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_140 = 5'hb == rob_tail ? io_dis_uops_0_inst : T_26182_11_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_141 = 5'hc == rob_tail ? io_dis_uops_0_inst : T_26182_12_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_142 = 5'hd == rob_tail ? io_dis_uops_0_inst : T_26182_13_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_143 = 5'he == rob_tail ? io_dis_uops_0_inst : T_26182_14_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_144 = 5'hf == rob_tail ? io_dis_uops_0_inst : T_26182_15_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_145 = 5'h10 == rob_tail ? io_dis_uops_0_inst : T_26182_16_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_146 = 5'h11 == rob_tail ? io_dis_uops_0_inst : T_26182_17_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_147 = 5'h12 == rob_tail ? io_dis_uops_0_inst : T_26182_18_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_148 = 5'h13 == rob_tail ? io_dis_uops_0_inst : T_26182_19_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_149 = 5'h14 == rob_tail ? io_dis_uops_0_inst : T_26182_20_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_150 = 5'h15 == rob_tail ? io_dis_uops_0_inst : T_26182_21_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_151 = 5'h16 == rob_tail ? io_dis_uops_0_inst : T_26182_22_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_152 = 5'h17 == rob_tail ? io_dis_uops_0_inst : T_26182_23_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_801 = 5'h0 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_0_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_802 = 5'h1 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_1_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_803 = 5'h2 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_2_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_804 = 5'h3 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_3_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_805 = 5'h4 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_4_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_806 = 5'h5 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_5_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_807 = 5'h6 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_6_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_808 = 5'h7 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_7_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_809 = 5'h8 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_8_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_810 = 5'h9 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_9_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_811 = 5'ha == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_10_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_812 = 5'hb == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_11_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_813 = 5'hc == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_12_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_814 = 5'hd == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_13_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_815 = 5'he == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_14_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_816 = 5'hf == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_15_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_817 = 5'h10 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_16_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_818 = 5'h11 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_17_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_819 = 5'h12 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_18_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_820 = 5'h13 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_19_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_821 = 5'h14 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_20_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_822 = 5'h15 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_21_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_823 = 5'h16 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_22_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_824 = 5'h17 == rob_tail ? io_dis_uops_0_stat_brjmp_mispredicted : T_26182_23_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_825 = 5'h0 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_0_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_826 = 5'h1 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_1_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_827 = 5'h2 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_2_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_828 = 5'h3 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_3_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_829 = 5'h4 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_4_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_830 = 5'h5 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_5_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_831 = 5'h6 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_6_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_832 = 5'h7 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_7_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_833 = 5'h8 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_8_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_834 = 5'h9 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_9_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_835 = 5'ha == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_10_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_836 = 5'hb == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_11_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_837 = 5'hc == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_12_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_838 = 5'hd == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_13_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_839 = 5'he == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_14_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_840 = 5'hf == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_15_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_841 = 5'h10 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_16_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_842 = 5'h11 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_17_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_843 = 5'h12 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_18_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_844 = 5'h13 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_19_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_845 = 5'h14 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_20_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_846 = 5'h15 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_21_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_847 = 5'h16 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_22_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_848 = 5'h17 == rob_tail ? io_dis_uops_0_stat_btb_made_pred : T_26182_23_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_849 = 5'h0 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_0_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_850 = 5'h1 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_1_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_851 = 5'h2 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_2_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_852 = 5'h3 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_3_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_853 = 5'h4 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_4_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_854 = 5'h5 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_5_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_855 = 5'h6 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_6_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_856 = 5'h7 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_7_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_857 = 5'h8 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_8_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_858 = 5'h9 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_9_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_859 = 5'ha == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_10_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_860 = 5'hb == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_11_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_861 = 5'hc == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_12_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_862 = 5'hd == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_13_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_863 = 5'he == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_14_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_864 = 5'hf == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_15_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_865 = 5'h10 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_16_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_866 = 5'h11 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_17_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_867 = 5'h12 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_18_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_868 = 5'h13 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_19_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_869 = 5'h14 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_20_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_870 = 5'h15 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_21_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_871 = 5'h16 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_22_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_872 = 5'h17 == rob_tail ? io_dis_uops_0_stat_btb_mispredicted : T_26182_23_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_873 = 5'h0 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_0_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_874 = 5'h1 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_1_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_875 = 5'h2 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_2_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_876 = 5'h3 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_3_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_877 = 5'h4 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_4_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_878 = 5'h5 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_5_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_879 = 5'h6 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_6_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_880 = 5'h7 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_7_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_881 = 5'h8 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_8_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_882 = 5'h9 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_9_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_883 = 5'ha == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_10_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_884 = 5'hb == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_11_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_885 = 5'hc == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_12_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_886 = 5'hd == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_13_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_887 = 5'he == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_14_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_888 = 5'hf == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_15_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_889 = 5'h10 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_16_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_890 = 5'h11 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_17_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_891 = 5'h12 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_18_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_892 = 5'h13 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_19_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_893 = 5'h14 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_20_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_894 = 5'h15 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_21_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_895 = 5'h16 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_22_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_896 = 5'h17 == rob_tail ? io_dis_uops_0_stat_bpd_made_pred : T_26182_23_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_897 = 5'h0 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_0_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_898 = 5'h1 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_1_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_899 = 5'h2 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_2_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_900 = 5'h3 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_3_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_901 = 5'h4 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_4_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_902 = 5'h5 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_5_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_903 = 5'h6 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_6_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_904 = 5'h7 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_7_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_905 = 5'h8 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_8_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_906 = 5'h9 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_9_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_907 = 5'ha == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_10_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_908 = 5'hb == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_11_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_909 = 5'hc == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_12_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_910 = 5'hd == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_13_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_911 = 5'he == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_14_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_912 = 5'hf == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_15_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_913 = 5'h10 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_16_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_914 = 5'h11 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_17_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_915 = 5'h12 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_18_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_916 = 5'h13 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_19_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_917 = 5'h14 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_20_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_918 = 5'h15 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_21_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_919 = 5'h16 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_22_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_920 = 5'h17 == rob_tail ? io_dis_uops_0_stat_bpd_mispredicted : T_26182_23_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1881 = 5'h0 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_0_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1882 = 5'h1 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_1_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1883 = 5'h2 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_2_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1884 = 5'h3 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_3_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1885 = 5'h4 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_4_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1886 = 5'h5 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_5_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1887 = 5'h6 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_6_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1888 = 5'h7 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_7_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1889 = 5'h8 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_8_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1890 = 5'h9 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_9_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1891 = 5'ha == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_10_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1892 = 5'hb == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_11_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1893 = 5'hc == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_12_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1894 = 5'hd == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_13_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1895 = 5'he == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_14_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1896 = 5'hf == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_15_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1897 = 5'h10 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_16_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1898 = 5'h11 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_17_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1899 = 5'h12 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_18_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1900 = 5'h13 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_19_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1901 = 5'h14 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_20_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1902 = 5'h15 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_21_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1903 = 5'h16 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_22_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_1904 = 5'h17 == rob_tail ? io_dis_uops_0_debug_wdata : T_26182_23_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_1929 = 5'h0 == rob_tail ? 1'h0 : _GEN_801; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1930 = 5'h1 == rob_tail ? 1'h0 : _GEN_802; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1931 = 5'h2 == rob_tail ? 1'h0 : _GEN_803; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1932 = 5'h3 == rob_tail ? 1'h0 : _GEN_804; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1933 = 5'h4 == rob_tail ? 1'h0 : _GEN_805; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1934 = 5'h5 == rob_tail ? 1'h0 : _GEN_806; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1935 = 5'h6 == rob_tail ? 1'h0 : _GEN_807; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1936 = 5'h7 == rob_tail ? 1'h0 : _GEN_808; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1937 = 5'h8 == rob_tail ? 1'h0 : _GEN_809; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1938 = 5'h9 == rob_tail ? 1'h0 : _GEN_810; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1939 = 5'ha == rob_tail ? 1'h0 : _GEN_811; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1940 = 5'hb == rob_tail ? 1'h0 : _GEN_812; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1941 = 5'hc == rob_tail ? 1'h0 : _GEN_813; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1942 = 5'hd == rob_tail ? 1'h0 : _GEN_814; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1943 = 5'he == rob_tail ? 1'h0 : _GEN_815; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1944 = 5'hf == rob_tail ? 1'h0 : _GEN_816; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1945 = 5'h10 == rob_tail ? 1'h0 : _GEN_817; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1946 = 5'h11 == rob_tail ? 1'h0 : _GEN_818; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1947 = 5'h12 == rob_tail ? 1'h0 : _GEN_819; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1948 = 5'h13 == rob_tail ? 1'h0 : _GEN_820; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1949 = 5'h14 == rob_tail ? 1'h0 : _GEN_821; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1950 = 5'h15 == rob_tail ? 1'h0 : _GEN_822; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1951 = 5'h16 == rob_tail ? 1'h0 : _GEN_823; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1952 = 5'h17 == rob_tail ? 1'h0 : _GEN_824; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_1953 = io_dis_valids_0 ? _GEN_33 : T_23706_0; // @[rob.scala 346:7]
  wire  _GEN_1954 = io_dis_valids_0 ? _GEN_34 : T_23706_1; // @[rob.scala 346:7]
  wire  _GEN_1955 = io_dis_valids_0 ? _GEN_35 : T_23706_2; // @[rob.scala 346:7]
  wire  _GEN_1956 = io_dis_valids_0 ? _GEN_36 : T_23706_3; // @[rob.scala 346:7]
  wire  _GEN_1957 = io_dis_valids_0 ? _GEN_37 : T_23706_4; // @[rob.scala 346:7]
  wire  _GEN_1958 = io_dis_valids_0 ? _GEN_38 : T_23706_5; // @[rob.scala 346:7]
  wire  _GEN_1959 = io_dis_valids_0 ? _GEN_39 : T_23706_6; // @[rob.scala 346:7]
  wire  _GEN_1960 = io_dis_valids_0 ? _GEN_40 : T_23706_7; // @[rob.scala 346:7]
  wire  _GEN_1961 = io_dis_valids_0 ? _GEN_41 : T_23706_8; // @[rob.scala 346:7]
  wire  _GEN_1962 = io_dis_valids_0 ? _GEN_42 : T_23706_9; // @[rob.scala 346:7]
  wire  _GEN_1963 = io_dis_valids_0 ? _GEN_43 : T_23706_10; // @[rob.scala 346:7]
  wire  _GEN_1964 = io_dis_valids_0 ? _GEN_44 : T_23706_11; // @[rob.scala 346:7]
  wire  _GEN_1965 = io_dis_valids_0 ? _GEN_45 : T_23706_12; // @[rob.scala 346:7]
  wire  _GEN_1966 = io_dis_valids_0 ? _GEN_46 : T_23706_13; // @[rob.scala 346:7]
  wire  _GEN_1967 = io_dis_valids_0 ? _GEN_47 : T_23706_14; // @[rob.scala 346:7]
  wire  _GEN_1968 = io_dis_valids_0 ? _GEN_48 : T_23706_15; // @[rob.scala 346:7]
  wire  _GEN_1969 = io_dis_valids_0 ? _GEN_49 : T_23706_16; // @[rob.scala 346:7]
  wire  _GEN_1970 = io_dis_valids_0 ? _GEN_50 : T_23706_17; // @[rob.scala 346:7]
  wire  _GEN_1971 = io_dis_valids_0 ? _GEN_51 : T_23706_18; // @[rob.scala 346:7]
  wire  _GEN_1972 = io_dis_valids_0 ? _GEN_52 : T_23706_19; // @[rob.scala 346:7]
  wire  _GEN_1973 = io_dis_valids_0 ? _GEN_53 : T_23706_20; // @[rob.scala 346:7]
  wire  _GEN_1974 = io_dis_valids_0 ? _GEN_54 : T_23706_21; // @[rob.scala 346:7]
  wire  _GEN_1975 = io_dis_valids_0 ? _GEN_55 : T_23706_22; // @[rob.scala 346:7]
  wire  _GEN_1976 = io_dis_valids_0 ? _GEN_56 : T_23706_23; // @[rob.scala 346:7]
  wire [31:0] _GEN_2054 = io_dis_valids_0 ? _GEN_129 : T_26182_0_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2055 = io_dis_valids_0 ? _GEN_130 : T_26182_1_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2056 = io_dis_valids_0 ? _GEN_131 : T_26182_2_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2057 = io_dis_valids_0 ? _GEN_132 : T_26182_3_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2058 = io_dis_valids_0 ? _GEN_133 : T_26182_4_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2059 = io_dis_valids_0 ? _GEN_134 : T_26182_5_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2060 = io_dis_valids_0 ? _GEN_135 : T_26182_6_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2061 = io_dis_valids_0 ? _GEN_136 : T_26182_7_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2062 = io_dis_valids_0 ? _GEN_137 : T_26182_8_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2063 = io_dis_valids_0 ? _GEN_138 : T_26182_9_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2064 = io_dis_valids_0 ? _GEN_139 : T_26182_10_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2065 = io_dis_valids_0 ? _GEN_140 : T_26182_11_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2066 = io_dis_valids_0 ? _GEN_141 : T_26182_12_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2067 = io_dis_valids_0 ? _GEN_142 : T_26182_13_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2068 = io_dis_valids_0 ? _GEN_143 : T_26182_14_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2069 = io_dis_valids_0 ? _GEN_144 : T_26182_15_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2070 = io_dis_valids_0 ? _GEN_145 : T_26182_16_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2071 = io_dis_valids_0 ? _GEN_146 : T_26182_17_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2072 = io_dis_valids_0 ? _GEN_147 : T_26182_18_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2073 = io_dis_valids_0 ? _GEN_148 : T_26182_19_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2074 = io_dis_valids_0 ? _GEN_149 : T_26182_20_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2075 = io_dis_valids_0 ? _GEN_150 : T_26182_21_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2076 = io_dis_valids_0 ? _GEN_151 : T_26182_22_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_2077 = io_dis_valids_0 ? _GEN_152 : T_26182_23_inst; // @[rob.scala 346:7]
  wire  _GEN_2726 = io_dis_valids_0 ? _GEN_1929 : T_26182_0_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2727 = io_dis_valids_0 ? _GEN_1930 : T_26182_1_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2728 = io_dis_valids_0 ? _GEN_1931 : T_26182_2_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2729 = io_dis_valids_0 ? _GEN_1932 : T_26182_3_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2730 = io_dis_valids_0 ? _GEN_1933 : T_26182_4_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2731 = io_dis_valids_0 ? _GEN_1934 : T_26182_5_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2732 = io_dis_valids_0 ? _GEN_1935 : T_26182_6_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2733 = io_dis_valids_0 ? _GEN_1936 : T_26182_7_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2734 = io_dis_valids_0 ? _GEN_1937 : T_26182_8_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2735 = io_dis_valids_0 ? _GEN_1938 : T_26182_9_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2736 = io_dis_valids_0 ? _GEN_1939 : T_26182_10_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2737 = io_dis_valids_0 ? _GEN_1940 : T_26182_11_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2738 = io_dis_valids_0 ? _GEN_1941 : T_26182_12_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2739 = io_dis_valids_0 ? _GEN_1942 : T_26182_13_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2740 = io_dis_valids_0 ? _GEN_1943 : T_26182_14_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2741 = io_dis_valids_0 ? _GEN_1944 : T_26182_15_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2742 = io_dis_valids_0 ? _GEN_1945 : T_26182_16_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2743 = io_dis_valids_0 ? _GEN_1946 : T_26182_17_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2744 = io_dis_valids_0 ? _GEN_1947 : T_26182_18_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2745 = io_dis_valids_0 ? _GEN_1948 : T_26182_19_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2746 = io_dis_valids_0 ? _GEN_1949 : T_26182_20_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2747 = io_dis_valids_0 ? _GEN_1950 : T_26182_21_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2748 = io_dis_valids_0 ? _GEN_1951 : T_26182_22_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2749 = io_dis_valids_0 ? _GEN_1952 : T_26182_23_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2750 = io_dis_valids_0 ? _GEN_825 : T_26182_0_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2751 = io_dis_valids_0 ? _GEN_826 : T_26182_1_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2752 = io_dis_valids_0 ? _GEN_827 : T_26182_2_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2753 = io_dis_valids_0 ? _GEN_828 : T_26182_3_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2754 = io_dis_valids_0 ? _GEN_829 : T_26182_4_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2755 = io_dis_valids_0 ? _GEN_830 : T_26182_5_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2756 = io_dis_valids_0 ? _GEN_831 : T_26182_6_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2757 = io_dis_valids_0 ? _GEN_832 : T_26182_7_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2758 = io_dis_valids_0 ? _GEN_833 : T_26182_8_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2759 = io_dis_valids_0 ? _GEN_834 : T_26182_9_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2760 = io_dis_valids_0 ? _GEN_835 : T_26182_10_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2761 = io_dis_valids_0 ? _GEN_836 : T_26182_11_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2762 = io_dis_valids_0 ? _GEN_837 : T_26182_12_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2763 = io_dis_valids_0 ? _GEN_838 : T_26182_13_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2764 = io_dis_valids_0 ? _GEN_839 : T_26182_14_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2765 = io_dis_valids_0 ? _GEN_840 : T_26182_15_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2766 = io_dis_valids_0 ? _GEN_841 : T_26182_16_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2767 = io_dis_valids_0 ? _GEN_842 : T_26182_17_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2768 = io_dis_valids_0 ? _GEN_843 : T_26182_18_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2769 = io_dis_valids_0 ? _GEN_844 : T_26182_19_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2770 = io_dis_valids_0 ? _GEN_845 : T_26182_20_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2771 = io_dis_valids_0 ? _GEN_846 : T_26182_21_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2772 = io_dis_valids_0 ? _GEN_847 : T_26182_22_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2773 = io_dis_valids_0 ? _GEN_848 : T_26182_23_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2774 = io_dis_valids_0 ? _GEN_849 : T_26182_0_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2775 = io_dis_valids_0 ? _GEN_850 : T_26182_1_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2776 = io_dis_valids_0 ? _GEN_851 : T_26182_2_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2777 = io_dis_valids_0 ? _GEN_852 : T_26182_3_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2778 = io_dis_valids_0 ? _GEN_853 : T_26182_4_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2779 = io_dis_valids_0 ? _GEN_854 : T_26182_5_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2780 = io_dis_valids_0 ? _GEN_855 : T_26182_6_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2781 = io_dis_valids_0 ? _GEN_856 : T_26182_7_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2782 = io_dis_valids_0 ? _GEN_857 : T_26182_8_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2783 = io_dis_valids_0 ? _GEN_858 : T_26182_9_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2784 = io_dis_valids_0 ? _GEN_859 : T_26182_10_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2785 = io_dis_valids_0 ? _GEN_860 : T_26182_11_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2786 = io_dis_valids_0 ? _GEN_861 : T_26182_12_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2787 = io_dis_valids_0 ? _GEN_862 : T_26182_13_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2788 = io_dis_valids_0 ? _GEN_863 : T_26182_14_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2789 = io_dis_valids_0 ? _GEN_864 : T_26182_15_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2790 = io_dis_valids_0 ? _GEN_865 : T_26182_16_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2791 = io_dis_valids_0 ? _GEN_866 : T_26182_17_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2792 = io_dis_valids_0 ? _GEN_867 : T_26182_18_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2793 = io_dis_valids_0 ? _GEN_868 : T_26182_19_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2794 = io_dis_valids_0 ? _GEN_869 : T_26182_20_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2795 = io_dis_valids_0 ? _GEN_870 : T_26182_21_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2796 = io_dis_valids_0 ? _GEN_871 : T_26182_22_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2797 = io_dis_valids_0 ? _GEN_872 : T_26182_23_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2798 = io_dis_valids_0 ? _GEN_873 : T_26182_0_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2799 = io_dis_valids_0 ? _GEN_874 : T_26182_1_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2800 = io_dis_valids_0 ? _GEN_875 : T_26182_2_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2801 = io_dis_valids_0 ? _GEN_876 : T_26182_3_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2802 = io_dis_valids_0 ? _GEN_877 : T_26182_4_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2803 = io_dis_valids_0 ? _GEN_878 : T_26182_5_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2804 = io_dis_valids_0 ? _GEN_879 : T_26182_6_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2805 = io_dis_valids_0 ? _GEN_880 : T_26182_7_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2806 = io_dis_valids_0 ? _GEN_881 : T_26182_8_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2807 = io_dis_valids_0 ? _GEN_882 : T_26182_9_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2808 = io_dis_valids_0 ? _GEN_883 : T_26182_10_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2809 = io_dis_valids_0 ? _GEN_884 : T_26182_11_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2810 = io_dis_valids_0 ? _GEN_885 : T_26182_12_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2811 = io_dis_valids_0 ? _GEN_886 : T_26182_13_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2812 = io_dis_valids_0 ? _GEN_887 : T_26182_14_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2813 = io_dis_valids_0 ? _GEN_888 : T_26182_15_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2814 = io_dis_valids_0 ? _GEN_889 : T_26182_16_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2815 = io_dis_valids_0 ? _GEN_890 : T_26182_17_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2816 = io_dis_valids_0 ? _GEN_891 : T_26182_18_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2817 = io_dis_valids_0 ? _GEN_892 : T_26182_19_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2818 = io_dis_valids_0 ? _GEN_893 : T_26182_20_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2819 = io_dis_valids_0 ? _GEN_894 : T_26182_21_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2820 = io_dis_valids_0 ? _GEN_895 : T_26182_22_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2821 = io_dis_valids_0 ? _GEN_896 : T_26182_23_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_2822 = io_dis_valids_0 ? _GEN_897 : T_26182_0_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2823 = io_dis_valids_0 ? _GEN_898 : T_26182_1_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2824 = io_dis_valids_0 ? _GEN_899 : T_26182_2_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2825 = io_dis_valids_0 ? _GEN_900 : T_26182_3_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2826 = io_dis_valids_0 ? _GEN_901 : T_26182_4_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2827 = io_dis_valids_0 ? _GEN_902 : T_26182_5_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2828 = io_dis_valids_0 ? _GEN_903 : T_26182_6_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2829 = io_dis_valids_0 ? _GEN_904 : T_26182_7_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2830 = io_dis_valids_0 ? _GEN_905 : T_26182_8_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2831 = io_dis_valids_0 ? _GEN_906 : T_26182_9_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2832 = io_dis_valids_0 ? _GEN_907 : T_26182_10_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2833 = io_dis_valids_0 ? _GEN_908 : T_26182_11_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2834 = io_dis_valids_0 ? _GEN_909 : T_26182_12_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2835 = io_dis_valids_0 ? _GEN_910 : T_26182_13_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2836 = io_dis_valids_0 ? _GEN_911 : T_26182_14_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2837 = io_dis_valids_0 ? _GEN_912 : T_26182_15_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2838 = io_dis_valids_0 ? _GEN_913 : T_26182_16_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2839 = io_dis_valids_0 ? _GEN_914 : T_26182_17_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2840 = io_dis_valids_0 ? _GEN_915 : T_26182_18_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2841 = io_dis_valids_0 ? _GEN_916 : T_26182_19_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2842 = io_dis_valids_0 ? _GEN_917 : T_26182_20_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2843 = io_dis_valids_0 ? _GEN_918 : T_26182_21_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2844 = io_dis_valids_0 ? _GEN_919 : T_26182_22_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_2845 = io_dis_valids_0 ? _GEN_920 : T_26182_23_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire [63:0] _GEN_3806 = io_dis_valids_0 ? _GEN_1881 : T_26182_0_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3807 = io_dis_valids_0 ? _GEN_1882 : T_26182_1_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3808 = io_dis_valids_0 ? _GEN_1883 : T_26182_2_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3809 = io_dis_valids_0 ? _GEN_1884 : T_26182_3_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3810 = io_dis_valids_0 ? _GEN_1885 : T_26182_4_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3811 = io_dis_valids_0 ? _GEN_1886 : T_26182_5_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3812 = io_dis_valids_0 ? _GEN_1887 : T_26182_6_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3813 = io_dis_valids_0 ? _GEN_1888 : T_26182_7_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3814 = io_dis_valids_0 ? _GEN_1889 : T_26182_8_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3815 = io_dis_valids_0 ? _GEN_1890 : T_26182_9_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3816 = io_dis_valids_0 ? _GEN_1891 : T_26182_10_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3817 = io_dis_valids_0 ? _GEN_1892 : T_26182_11_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3818 = io_dis_valids_0 ? _GEN_1893 : T_26182_12_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3819 = io_dis_valids_0 ? _GEN_1894 : T_26182_13_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3820 = io_dis_valids_0 ? _GEN_1895 : T_26182_14_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3821 = io_dis_valids_0 ? _GEN_1896 : T_26182_15_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3822 = io_dis_valids_0 ? _GEN_1897 : T_26182_16_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3823 = io_dis_valids_0 ? _GEN_1898 : T_26182_17_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3824 = io_dis_valids_0 ? _GEN_1899 : T_26182_18_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3825 = io_dis_valids_0 ? _GEN_1900 : T_26182_19_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3826 = io_dis_valids_0 ? _GEN_1901 : T_26182_20_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3827 = io_dis_valids_0 ? _GEN_1902 : T_26182_21_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3828 = io_dis_valids_0 ? _GEN_1903 : T_26182_22_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_3829 = io_dis_valids_0 ? _GEN_1904 : T_26182_23_debug_wdata; // @[rob.scala 346:7]
  wire  _GEN_3857 = 5'h1 == rob_tail ? T_23706_1 : T_23706_0; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3858 = 5'h2 == rob_tail ? T_23706_2 : _GEN_3857; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3859 = 5'h3 == rob_tail ? T_23706_3 : _GEN_3858; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3860 = 5'h4 == rob_tail ? T_23706_4 : _GEN_3859; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3861 = 5'h5 == rob_tail ? T_23706_5 : _GEN_3860; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3862 = 5'h6 == rob_tail ? T_23706_6 : _GEN_3861; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3863 = 5'h7 == rob_tail ? T_23706_7 : _GEN_3862; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3864 = 5'h8 == rob_tail ? T_23706_8 : _GEN_3863; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3865 = 5'h9 == rob_tail ? T_23706_9 : _GEN_3864; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3866 = 5'ha == rob_tail ? T_23706_10 : _GEN_3865; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3867 = 5'hb == rob_tail ? T_23706_11 : _GEN_3866; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3868 = 5'hc == rob_tail ? T_23706_12 : _GEN_3867; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3869 = 5'hd == rob_tail ? T_23706_13 : _GEN_3868; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3870 = 5'he == rob_tail ? T_23706_14 : _GEN_3869; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3871 = 5'hf == rob_tail ? T_23706_15 : _GEN_3870; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3872 = 5'h10 == rob_tail ? T_23706_16 : _GEN_3871; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3873 = 5'h11 == rob_tail ? T_23706_17 : _GEN_3872; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3874 = 5'h12 == rob_tail ? T_23706_18 : _GEN_3873; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3875 = 5'h13 == rob_tail ? T_23706_19 : _GEN_3874; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3876 = 5'h14 == rob_tail ? T_23706_20 : _GEN_3875; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3877 = 5'h15 == rob_tail ? T_23706_21 : _GEN_3876; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3878 = 5'h16 == rob_tail ? T_23706_22 : _GEN_3877; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_3879 = 5'h17 == rob_tail ? T_23706_23 : _GEN_3878; // @[rob.scala 355:47 rob.scala 355:47]
  wire  T_28498 = ~_GEN_3879; // @[rob.scala 355:47]
  wire  T_28499 = T_23559 & T_28498; // @[rob.scala 355:44]
  wire  T_28501 = ~io_dis_valids_0; // @[rob.scala 346:7]
  wire  T_28502 = T_28501 & T_28499; // @[rob.scala 356:7]
  wire [31:0] _GEN_3880 = 5'h0 == rob_tail ? 32'h4033 : _GEN_2054; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3881 = 5'h1 == rob_tail ? 32'h4033 : _GEN_2055; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3882 = 5'h2 == rob_tail ? 32'h4033 : _GEN_2056; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3883 = 5'h3 == rob_tail ? 32'h4033 : _GEN_2057; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3884 = 5'h4 == rob_tail ? 32'h4033 : _GEN_2058; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3885 = 5'h5 == rob_tail ? 32'h4033 : _GEN_2059; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3886 = 5'h6 == rob_tail ? 32'h4033 : _GEN_2060; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3887 = 5'h7 == rob_tail ? 32'h4033 : _GEN_2061; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3888 = 5'h8 == rob_tail ? 32'h4033 : _GEN_2062; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3889 = 5'h9 == rob_tail ? 32'h4033 : _GEN_2063; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3890 = 5'ha == rob_tail ? 32'h4033 : _GEN_2064; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3891 = 5'hb == rob_tail ? 32'h4033 : _GEN_2065; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3892 = 5'hc == rob_tail ? 32'h4033 : _GEN_2066; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3893 = 5'hd == rob_tail ? 32'h4033 : _GEN_2067; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3894 = 5'he == rob_tail ? 32'h4033 : _GEN_2068; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3895 = 5'hf == rob_tail ? 32'h4033 : _GEN_2069; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3896 = 5'h10 == rob_tail ? 32'h4033 : _GEN_2070; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3897 = 5'h11 == rob_tail ? 32'h4033 : _GEN_2071; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3898 = 5'h12 == rob_tail ? 32'h4033 : _GEN_2072; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3899 = 5'h13 == rob_tail ? 32'h4033 : _GEN_2073; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3900 = 5'h14 == rob_tail ? 32'h4033 : _GEN_2074; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3901 = 5'h15 == rob_tail ? 32'h4033 : _GEN_2075; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3902 = 5'h16 == rob_tail ? 32'h4033 : _GEN_2076; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3903 = 5'h17 == rob_tail ? 32'h4033 : _GEN_2077; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_3904 = T_28502 ? _GEN_3880 : _GEN_2054; // @[rob.scala 356:7]
  wire [31:0] _GEN_3905 = T_28502 ? _GEN_3881 : _GEN_2055; // @[rob.scala 356:7]
  wire [31:0] _GEN_3906 = T_28502 ? _GEN_3882 : _GEN_2056; // @[rob.scala 356:7]
  wire [31:0] _GEN_3907 = T_28502 ? _GEN_3883 : _GEN_2057; // @[rob.scala 356:7]
  wire [31:0] _GEN_3908 = T_28502 ? _GEN_3884 : _GEN_2058; // @[rob.scala 356:7]
  wire [31:0] _GEN_3909 = T_28502 ? _GEN_3885 : _GEN_2059; // @[rob.scala 356:7]
  wire [31:0] _GEN_3910 = T_28502 ? _GEN_3886 : _GEN_2060; // @[rob.scala 356:7]
  wire [31:0] _GEN_3911 = T_28502 ? _GEN_3887 : _GEN_2061; // @[rob.scala 356:7]
  wire [31:0] _GEN_3912 = T_28502 ? _GEN_3888 : _GEN_2062; // @[rob.scala 356:7]
  wire [31:0] _GEN_3913 = T_28502 ? _GEN_3889 : _GEN_2063; // @[rob.scala 356:7]
  wire [31:0] _GEN_3914 = T_28502 ? _GEN_3890 : _GEN_2064; // @[rob.scala 356:7]
  wire [31:0] _GEN_3915 = T_28502 ? _GEN_3891 : _GEN_2065; // @[rob.scala 356:7]
  wire [31:0] _GEN_3916 = T_28502 ? _GEN_3892 : _GEN_2066; // @[rob.scala 356:7]
  wire [31:0] _GEN_3917 = T_28502 ? _GEN_3893 : _GEN_2067; // @[rob.scala 356:7]
  wire [31:0] _GEN_3918 = T_28502 ? _GEN_3894 : _GEN_2068; // @[rob.scala 356:7]
  wire [31:0] _GEN_3919 = T_28502 ? _GEN_3895 : _GEN_2069; // @[rob.scala 356:7]
  wire [31:0] _GEN_3920 = T_28502 ? _GEN_3896 : _GEN_2070; // @[rob.scala 356:7]
  wire [31:0] _GEN_3921 = T_28502 ? _GEN_3897 : _GEN_2071; // @[rob.scala 356:7]
  wire [31:0] _GEN_3922 = T_28502 ? _GEN_3898 : _GEN_2072; // @[rob.scala 356:7]
  wire [31:0] _GEN_3923 = T_28502 ? _GEN_3899 : _GEN_2073; // @[rob.scala 356:7]
  wire [31:0] _GEN_3924 = T_28502 ? _GEN_3900 : _GEN_2074; // @[rob.scala 356:7]
  wire [31:0] _GEN_3925 = T_28502 ? _GEN_3901 : _GEN_2075; // @[rob.scala 356:7]
  wire [31:0] _GEN_3926 = T_28502 ? _GEN_3902 : _GEN_2076; // @[rob.scala 356:7]
  wire [31:0] _GEN_3927 = T_28502 ? _GEN_3903 : _GEN_2077; // @[rob.scala 356:7]
  wire [5:0] T_28589 = {{1'd0}, io_wb_resps_0_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_28590 = io_wb_resps_0_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_28592 = ~T_28590; // @[rob.scala 331:55]
  wire  T_28593 = io_wb_resps_0_valid & T_28592; // @[rob.scala 368:30]
  wire [5:0] T_28597 = {{1'd0}, io_wb_resps_1_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_28598 = io_wb_resps_1_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_28600 = ~T_28598; // @[rob.scala 331:55]
  wire  T_28601 = io_wb_resps_1_valid & T_28600; // @[rob.scala 368:30]
  wire [5:0] T_28605 = {{1'd0}, io_wb_resps_2_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_28606 = io_wb_resps_2_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_28608 = ~T_28606; // @[rob.scala 331:55]
  wire  T_28609 = io_wb_resps_2_valid & T_28608; // @[rob.scala 368:30]
  wire  T_28612 = io_lsu_clr_bsy_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_28614 = ~T_28612; // @[rob.scala 331:55]
  wire [5:0] T_28617 = {{1'd0}, io_lsu_clr_bsy_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_28620 = io_brinfo_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_28622 = ~T_28620; // @[rob.scala 331:55]
  wire  T_28623 = io_brinfo_valid & T_28622; // @[rob.scala 400:29]
  wire [5:0] T_28625 = {{1'd0}, io_brinfo_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_29059 = io_fflags_0_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_29061 = ~T_29059; // @[rob.scala 331:55]
  wire [5:0] T_29064 = {{1'd0}, io_fflags_0_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_29066 = io_fflags_1_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_29068 = ~T_29066; // @[rob.scala 331:55]
  wire [5:0] T_29071 = {{1'd0}, io_fflags_1_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_29073 = io_lxcpt_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_29075 = ~T_29073; // @[rob.scala 331:55]
  wire [5:0] T_29078 = {{1'd0}, io_lxcpt_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_29081 = io_bxcpt_bits_uop_rob_idx[0]; // @[rob.scala 227:38]
  wire  T_29083 = ~T_29081; // @[rob.scala 331:55]
  wire [5:0] T_29086 = {{1'd0}, io_bxcpt_bits_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire  T_29097 = rob_state == 2'h2; // @[rob.scala 443:23]
  wire [4:0] T_29096 = T_29097 ? rob_tail : rob_head; // @[rob.scala 444:7 rob.scala 445:18 rob.scala 442:15]
  wire  _GEN_4232 = 5'h1 == T_29096 ? T_23706_1 : T_23706_0; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4233 = 5'h2 == T_29096 ? T_23706_2 : _GEN_4232; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4234 = 5'h3 == T_29096 ? T_23706_3 : _GEN_4233; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4235 = 5'h4 == T_29096 ? T_23706_4 : _GEN_4234; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4236 = 5'h5 == T_29096 ? T_23706_5 : _GEN_4235; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4237 = 5'h6 == T_29096 ? T_23706_6 : _GEN_4236; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4238 = 5'h7 == T_29096 ? T_23706_7 : _GEN_4237; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4239 = 5'h8 == T_29096 ? T_23706_8 : _GEN_4238; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4240 = 5'h9 == T_29096 ? T_23706_9 : _GEN_4239; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4241 = 5'ha == T_29096 ? T_23706_10 : _GEN_4240; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4242 = 5'hb == T_29096 ? T_23706_11 : _GEN_4241; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4243 = 5'hc == T_29096 ? T_23706_12 : _GEN_4242; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4244 = 5'hd == T_29096 ? T_23706_13 : _GEN_4243; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4245 = 5'he == T_29096 ? T_23706_14 : _GEN_4244; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4246 = 5'hf == T_29096 ? T_23706_15 : _GEN_4245; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4247 = 5'h10 == T_29096 ? T_23706_16 : _GEN_4246; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4248 = 5'h11 == T_29096 ? T_23706_17 : _GEN_4247; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4249 = 5'h12 == T_29096 ? T_23706_18 : _GEN_4248; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4250 = 5'h13 == T_29096 ? T_23706_19 : _GEN_4249; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4251 = 5'h14 == T_29096 ? T_23706_20 : _GEN_4250; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4252 = 5'h15 == T_29096 ? T_23706_21 : _GEN_4251; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4253 = 5'h16 == T_29096 ? T_23706_22 : _GEN_4252; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_4254 = 5'h17 == T_29096 ? T_23706_23 : _GEN_4253; // @[rob.scala 451:58 rob.scala 451:58]
  wire  T_29099 = T_29097 & _GEN_4254; // @[rob.scala 451:58]
  wire  _GEN_4333 = 5'h1 == T_29096 ? T_26182_1_valid : T_26182_0_valid; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4334 = 5'h1 == T_29096 ? T_26182_1_iw_state : T_26182_0_iw_state; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4335 = 5'h1 == T_29096 ? T_26182_1_uopc : T_26182_0_uopc; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4336 = 5'h1 == T_29096 ? T_26182_1_inst : T_26182_0_inst; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4337 = 5'h1 == T_29096 ? T_26182_1_pc : T_26182_0_pc; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4338 = 5'h1 == T_29096 ? T_26182_1_fu_code : T_26182_0_fu_code; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4339 = 5'h1 == T_29096 ? T_26182_1_ctrl_br_type : T_26182_0_ctrl_br_type; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4340 = 5'h1 == T_29096 ? T_26182_1_ctrl_op1_sel : T_26182_0_ctrl_op1_sel; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4341 = 5'h1 == T_29096 ? T_26182_1_ctrl_op2_sel : T_26182_0_ctrl_op2_sel; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4342 = 5'h1 == T_29096 ? T_26182_1_ctrl_imm_sel : T_26182_0_ctrl_imm_sel; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4343 = 5'h1 == T_29096 ? T_26182_1_ctrl_op_fcn : T_26182_0_ctrl_op_fcn; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4344 = 5'h1 == T_29096 ? T_26182_1_ctrl_fcn_dw : T_26182_0_ctrl_fcn_dw; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4345 = 5'h1 == T_29096 ? T_26182_1_ctrl_rf_wen : T_26182_0_ctrl_rf_wen; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4346 = 5'h1 == T_29096 ? T_26182_1_ctrl_csr_cmd : T_26182_0_ctrl_csr_cmd; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4347 = 5'h1 == T_29096 ? T_26182_1_ctrl_is_load : T_26182_0_ctrl_is_load; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4348 = 5'h1 == T_29096 ? T_26182_1_ctrl_is_sta : T_26182_0_ctrl_is_sta; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4349 = 5'h1 == T_29096 ? T_26182_1_ctrl_is_std : T_26182_0_ctrl_is_std; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4350 = 5'h1 == T_29096 ? T_26182_1_wakeup_delay : T_26182_0_wakeup_delay; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4351 = 5'h1 == T_29096 ? T_26182_1_allocate_brtag : T_26182_0_allocate_brtag; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4352 = 5'h1 == T_29096 ? T_26182_1_is_br_or_jmp : T_26182_0_is_br_or_jmp; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4353 = 5'h1 == T_29096 ? T_26182_1_is_jump : T_26182_0_is_jump; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4354 = 5'h1 == T_29096 ? T_26182_1_is_jal : T_26182_0_is_jal; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4355 = 5'h1 == T_29096 ? T_26182_1_is_ret : T_26182_0_is_ret; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4356 = 5'h1 == T_29096 ? T_26182_1_is_call : T_26182_0_is_call; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4357 = 5'h1 == T_29096 ? T_26182_1_br_mask : T_26182_0_br_mask; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4358 = 5'h1 == T_29096 ? T_26182_1_br_tag : T_26182_0_br_tag; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4359 = 5'h1 == T_29096 ? T_26182_1_br_prediction_bpd_predict_val : T_26182_0_br_prediction_bpd_predict_val; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4360 = 5'h1 == T_29096 ? T_26182_1_br_prediction_bpd_predict_taken :
    T_26182_0_br_prediction_bpd_predict_taken; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4361 = 5'h1 == T_29096 ? T_26182_1_br_prediction_btb_hit : T_26182_0_br_prediction_btb_hit; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4362 = 5'h1 == T_29096 ? T_26182_1_br_prediction_btb_predicted : T_26182_0_br_prediction_btb_predicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4363 = 5'h1 == T_29096 ? T_26182_1_br_prediction_is_br_or_jalr : T_26182_0_br_prediction_is_br_or_jalr; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4364 = 5'h1 == T_29096 ? T_26182_1_stat_brjmp_mispredicted : T_26182_0_stat_brjmp_mispredicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4365 = 5'h1 == T_29096 ? T_26182_1_stat_btb_made_pred : T_26182_0_stat_btb_made_pred; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4366 = 5'h1 == T_29096 ? T_26182_1_stat_btb_mispredicted : T_26182_0_stat_btb_mispredicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4367 = 5'h1 == T_29096 ? T_26182_1_stat_bpd_made_pred : T_26182_0_stat_bpd_made_pred; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4368 = 5'h1 == T_29096 ? T_26182_1_stat_bpd_mispredicted : T_26182_0_stat_bpd_mispredicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4369 = 5'h1 == T_29096 ? T_26182_1_fetch_pc_lob : T_26182_0_fetch_pc_lob; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4370 = 5'h1 == T_29096 ? T_26182_1_imm_packed : T_26182_0_imm_packed; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4371 = 5'h1 == T_29096 ? T_26182_1_csr_addr : T_26182_0_csr_addr; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4372 = 5'h1 == T_29096 ? T_26182_1_rob_idx : T_26182_0_rob_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4373 = 5'h1 == T_29096 ? T_26182_1_ldq_idx : T_26182_0_ldq_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4374 = 5'h1 == T_29096 ? T_26182_1_stq_idx : T_26182_0_stq_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4375 = 5'h1 == T_29096 ? T_26182_1_brob_idx : T_26182_0_brob_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4376 = 5'h1 == T_29096 ? T_26182_1_pdst : T_26182_0_pdst; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4377 = 5'h1 == T_29096 ? T_26182_1_pop1 : T_26182_0_pop1; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4378 = 5'h1 == T_29096 ? T_26182_1_pop2 : T_26182_0_pop2; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4379 = 5'h1 == T_29096 ? T_26182_1_pop3 : T_26182_0_pop3; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4380 = 5'h1 == T_29096 ? T_26182_1_prs1_busy : T_26182_0_prs1_busy; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4381 = 5'h1 == T_29096 ? T_26182_1_prs2_busy : T_26182_0_prs2_busy; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4382 = 5'h1 == T_29096 ? T_26182_1_prs3_busy : T_26182_0_prs3_busy; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4383 = 5'h1 == T_29096 ? T_26182_1_stale_pdst : T_26182_0_stale_pdst; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4384 = 5'h1 == T_29096 ? T_26182_1_exception : T_26182_0_exception; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4385 = 5'h1 == T_29096 ? T_26182_1_exc_cause : T_26182_0_exc_cause; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4386 = 5'h1 == T_29096 ? T_26182_1_bypassable : T_26182_0_bypassable; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4387 = 5'h1 == T_29096 ? T_26182_1_mem_cmd : T_26182_0_mem_cmd; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4388 = 5'h1 == T_29096 ? T_26182_1_mem_typ : T_26182_0_mem_typ; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4389 = 5'h1 == T_29096 ? T_26182_1_is_fence : T_26182_0_is_fence; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4390 = 5'h1 == T_29096 ? T_26182_1_is_fencei : T_26182_0_is_fencei; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4391 = 5'h1 == T_29096 ? T_26182_1_is_store : T_26182_0_is_store; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4392 = 5'h1 == T_29096 ? T_26182_1_is_amo : T_26182_0_is_amo; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4393 = 5'h1 == T_29096 ? T_26182_1_is_load : T_26182_0_is_load; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4394 = 5'h1 == T_29096 ? T_26182_1_is_unique : T_26182_0_is_unique; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4395 = 5'h1 == T_29096 ? T_26182_1_flush_on_commit : T_26182_0_flush_on_commit; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4396 = 5'h1 == T_29096 ? T_26182_1_ldst : T_26182_0_ldst; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4397 = 5'h1 == T_29096 ? T_26182_1_lrs1 : T_26182_0_lrs1; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4398 = 5'h1 == T_29096 ? T_26182_1_lrs2 : T_26182_0_lrs2; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4399 = 5'h1 == T_29096 ? T_26182_1_lrs3 : T_26182_0_lrs3; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4400 = 5'h1 == T_29096 ? T_26182_1_ldst_val : T_26182_0_ldst_val; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4401 = 5'h1 == T_29096 ? T_26182_1_dst_rtype : T_26182_0_dst_rtype; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4402 = 5'h1 == T_29096 ? T_26182_1_lrs1_rtype : T_26182_0_lrs1_rtype; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4403 = 5'h1 == T_29096 ? T_26182_1_lrs2_rtype : T_26182_0_lrs2_rtype; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4404 = 5'h1 == T_29096 ? T_26182_1_frs3_en : T_26182_0_frs3_en; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4405 = 5'h1 == T_29096 ? T_26182_1_fp_val : T_26182_0_fp_val; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4406 = 5'h1 == T_29096 ? T_26182_1_fp_single : T_26182_0_fp_single; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4407 = 5'h1 == T_29096 ? T_26182_1_xcpt_if : T_26182_0_xcpt_if; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4408 = 5'h1 == T_29096 ? T_26182_1_replay_if : T_26182_0_replay_if; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4410 = 5'h1 == T_29096 ? T_26182_1_debug_events_fetch_seq : T_26182_0_debug_events_fetch_seq; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4411 = 5'h2 == T_29096 ? T_26182_2_valid : _GEN_4333; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4412 = 5'h2 == T_29096 ? T_26182_2_iw_state : _GEN_4334; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4413 = 5'h2 == T_29096 ? T_26182_2_uopc : _GEN_4335; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4414 = 5'h2 == T_29096 ? T_26182_2_inst : _GEN_4336; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4415 = 5'h2 == T_29096 ? T_26182_2_pc : _GEN_4337; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4416 = 5'h2 == T_29096 ? T_26182_2_fu_code : _GEN_4338; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4417 = 5'h2 == T_29096 ? T_26182_2_ctrl_br_type : _GEN_4339; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4418 = 5'h2 == T_29096 ? T_26182_2_ctrl_op1_sel : _GEN_4340; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4419 = 5'h2 == T_29096 ? T_26182_2_ctrl_op2_sel : _GEN_4341; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4420 = 5'h2 == T_29096 ? T_26182_2_ctrl_imm_sel : _GEN_4342; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4421 = 5'h2 == T_29096 ? T_26182_2_ctrl_op_fcn : _GEN_4343; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4422 = 5'h2 == T_29096 ? T_26182_2_ctrl_fcn_dw : _GEN_4344; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4423 = 5'h2 == T_29096 ? T_26182_2_ctrl_rf_wen : _GEN_4345; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4424 = 5'h2 == T_29096 ? T_26182_2_ctrl_csr_cmd : _GEN_4346; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4425 = 5'h2 == T_29096 ? T_26182_2_ctrl_is_load : _GEN_4347; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4426 = 5'h2 == T_29096 ? T_26182_2_ctrl_is_sta : _GEN_4348; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4427 = 5'h2 == T_29096 ? T_26182_2_ctrl_is_std : _GEN_4349; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4428 = 5'h2 == T_29096 ? T_26182_2_wakeup_delay : _GEN_4350; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4429 = 5'h2 == T_29096 ? T_26182_2_allocate_brtag : _GEN_4351; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4430 = 5'h2 == T_29096 ? T_26182_2_is_br_or_jmp : _GEN_4352; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4431 = 5'h2 == T_29096 ? T_26182_2_is_jump : _GEN_4353; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4432 = 5'h2 == T_29096 ? T_26182_2_is_jal : _GEN_4354; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4433 = 5'h2 == T_29096 ? T_26182_2_is_ret : _GEN_4355; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4434 = 5'h2 == T_29096 ? T_26182_2_is_call : _GEN_4356; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4435 = 5'h2 == T_29096 ? T_26182_2_br_mask : _GEN_4357; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4436 = 5'h2 == T_29096 ? T_26182_2_br_tag : _GEN_4358; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4437 = 5'h2 == T_29096 ? T_26182_2_br_prediction_bpd_predict_val : _GEN_4359; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4438 = 5'h2 == T_29096 ? T_26182_2_br_prediction_bpd_predict_taken : _GEN_4360; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4439 = 5'h2 == T_29096 ? T_26182_2_br_prediction_btb_hit : _GEN_4361; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4440 = 5'h2 == T_29096 ? T_26182_2_br_prediction_btb_predicted : _GEN_4362; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4441 = 5'h2 == T_29096 ? T_26182_2_br_prediction_is_br_or_jalr : _GEN_4363; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4442 = 5'h2 == T_29096 ? T_26182_2_stat_brjmp_mispredicted : _GEN_4364; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4443 = 5'h2 == T_29096 ? T_26182_2_stat_btb_made_pred : _GEN_4365; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4444 = 5'h2 == T_29096 ? T_26182_2_stat_btb_mispredicted : _GEN_4366; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4445 = 5'h2 == T_29096 ? T_26182_2_stat_bpd_made_pred : _GEN_4367; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4446 = 5'h2 == T_29096 ? T_26182_2_stat_bpd_mispredicted : _GEN_4368; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4447 = 5'h2 == T_29096 ? T_26182_2_fetch_pc_lob : _GEN_4369; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4448 = 5'h2 == T_29096 ? T_26182_2_imm_packed : _GEN_4370; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4449 = 5'h2 == T_29096 ? T_26182_2_csr_addr : _GEN_4371; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4450 = 5'h2 == T_29096 ? T_26182_2_rob_idx : _GEN_4372; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4451 = 5'h2 == T_29096 ? T_26182_2_ldq_idx : _GEN_4373; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4452 = 5'h2 == T_29096 ? T_26182_2_stq_idx : _GEN_4374; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4453 = 5'h2 == T_29096 ? T_26182_2_brob_idx : _GEN_4375; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4454 = 5'h2 == T_29096 ? T_26182_2_pdst : _GEN_4376; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4455 = 5'h2 == T_29096 ? T_26182_2_pop1 : _GEN_4377; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4456 = 5'h2 == T_29096 ? T_26182_2_pop2 : _GEN_4378; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4457 = 5'h2 == T_29096 ? T_26182_2_pop3 : _GEN_4379; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4458 = 5'h2 == T_29096 ? T_26182_2_prs1_busy : _GEN_4380; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4459 = 5'h2 == T_29096 ? T_26182_2_prs2_busy : _GEN_4381; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4460 = 5'h2 == T_29096 ? T_26182_2_prs3_busy : _GEN_4382; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4461 = 5'h2 == T_29096 ? T_26182_2_stale_pdst : _GEN_4383; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4462 = 5'h2 == T_29096 ? T_26182_2_exception : _GEN_4384; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4463 = 5'h2 == T_29096 ? T_26182_2_exc_cause : _GEN_4385; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4464 = 5'h2 == T_29096 ? T_26182_2_bypassable : _GEN_4386; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4465 = 5'h2 == T_29096 ? T_26182_2_mem_cmd : _GEN_4387; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4466 = 5'h2 == T_29096 ? T_26182_2_mem_typ : _GEN_4388; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4467 = 5'h2 == T_29096 ? T_26182_2_is_fence : _GEN_4389; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4468 = 5'h2 == T_29096 ? T_26182_2_is_fencei : _GEN_4390; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4469 = 5'h2 == T_29096 ? T_26182_2_is_store : _GEN_4391; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4470 = 5'h2 == T_29096 ? T_26182_2_is_amo : _GEN_4392; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4471 = 5'h2 == T_29096 ? T_26182_2_is_load : _GEN_4393; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4472 = 5'h2 == T_29096 ? T_26182_2_is_unique : _GEN_4394; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4473 = 5'h2 == T_29096 ? T_26182_2_flush_on_commit : _GEN_4395; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4474 = 5'h2 == T_29096 ? T_26182_2_ldst : _GEN_4396; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4475 = 5'h2 == T_29096 ? T_26182_2_lrs1 : _GEN_4397; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4476 = 5'h2 == T_29096 ? T_26182_2_lrs2 : _GEN_4398; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4477 = 5'h2 == T_29096 ? T_26182_2_lrs3 : _GEN_4399; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4478 = 5'h2 == T_29096 ? T_26182_2_ldst_val : _GEN_4400; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4479 = 5'h2 == T_29096 ? T_26182_2_dst_rtype : _GEN_4401; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4480 = 5'h2 == T_29096 ? T_26182_2_lrs1_rtype : _GEN_4402; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4481 = 5'h2 == T_29096 ? T_26182_2_lrs2_rtype : _GEN_4403; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4482 = 5'h2 == T_29096 ? T_26182_2_frs3_en : _GEN_4404; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4483 = 5'h2 == T_29096 ? T_26182_2_fp_val : _GEN_4405; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4484 = 5'h2 == T_29096 ? T_26182_2_fp_single : _GEN_4406; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4485 = 5'h2 == T_29096 ? T_26182_2_xcpt_if : _GEN_4407; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4486 = 5'h2 == T_29096 ? T_26182_2_replay_if : _GEN_4408; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4488 = 5'h2 == T_29096 ? T_26182_2_debug_events_fetch_seq : _GEN_4410; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4489 = 5'h3 == T_29096 ? T_26182_3_valid : _GEN_4411; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4490 = 5'h3 == T_29096 ? T_26182_3_iw_state : _GEN_4412; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4491 = 5'h3 == T_29096 ? T_26182_3_uopc : _GEN_4413; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4492 = 5'h3 == T_29096 ? T_26182_3_inst : _GEN_4414; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4493 = 5'h3 == T_29096 ? T_26182_3_pc : _GEN_4415; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4494 = 5'h3 == T_29096 ? T_26182_3_fu_code : _GEN_4416; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4495 = 5'h3 == T_29096 ? T_26182_3_ctrl_br_type : _GEN_4417; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4496 = 5'h3 == T_29096 ? T_26182_3_ctrl_op1_sel : _GEN_4418; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4497 = 5'h3 == T_29096 ? T_26182_3_ctrl_op2_sel : _GEN_4419; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4498 = 5'h3 == T_29096 ? T_26182_3_ctrl_imm_sel : _GEN_4420; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4499 = 5'h3 == T_29096 ? T_26182_3_ctrl_op_fcn : _GEN_4421; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4500 = 5'h3 == T_29096 ? T_26182_3_ctrl_fcn_dw : _GEN_4422; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4501 = 5'h3 == T_29096 ? T_26182_3_ctrl_rf_wen : _GEN_4423; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4502 = 5'h3 == T_29096 ? T_26182_3_ctrl_csr_cmd : _GEN_4424; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4503 = 5'h3 == T_29096 ? T_26182_3_ctrl_is_load : _GEN_4425; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4504 = 5'h3 == T_29096 ? T_26182_3_ctrl_is_sta : _GEN_4426; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4505 = 5'h3 == T_29096 ? T_26182_3_ctrl_is_std : _GEN_4427; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4506 = 5'h3 == T_29096 ? T_26182_3_wakeup_delay : _GEN_4428; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4507 = 5'h3 == T_29096 ? T_26182_3_allocate_brtag : _GEN_4429; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4508 = 5'h3 == T_29096 ? T_26182_3_is_br_or_jmp : _GEN_4430; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4509 = 5'h3 == T_29096 ? T_26182_3_is_jump : _GEN_4431; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4510 = 5'h3 == T_29096 ? T_26182_3_is_jal : _GEN_4432; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4511 = 5'h3 == T_29096 ? T_26182_3_is_ret : _GEN_4433; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4512 = 5'h3 == T_29096 ? T_26182_3_is_call : _GEN_4434; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4513 = 5'h3 == T_29096 ? T_26182_3_br_mask : _GEN_4435; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4514 = 5'h3 == T_29096 ? T_26182_3_br_tag : _GEN_4436; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4515 = 5'h3 == T_29096 ? T_26182_3_br_prediction_bpd_predict_val : _GEN_4437; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4516 = 5'h3 == T_29096 ? T_26182_3_br_prediction_bpd_predict_taken : _GEN_4438; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4517 = 5'h3 == T_29096 ? T_26182_3_br_prediction_btb_hit : _GEN_4439; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4518 = 5'h3 == T_29096 ? T_26182_3_br_prediction_btb_predicted : _GEN_4440; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4519 = 5'h3 == T_29096 ? T_26182_3_br_prediction_is_br_or_jalr : _GEN_4441; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4520 = 5'h3 == T_29096 ? T_26182_3_stat_brjmp_mispredicted : _GEN_4442; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4521 = 5'h3 == T_29096 ? T_26182_3_stat_btb_made_pred : _GEN_4443; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4522 = 5'h3 == T_29096 ? T_26182_3_stat_btb_mispredicted : _GEN_4444; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4523 = 5'h3 == T_29096 ? T_26182_3_stat_bpd_made_pred : _GEN_4445; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4524 = 5'h3 == T_29096 ? T_26182_3_stat_bpd_mispredicted : _GEN_4446; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4525 = 5'h3 == T_29096 ? T_26182_3_fetch_pc_lob : _GEN_4447; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4526 = 5'h3 == T_29096 ? T_26182_3_imm_packed : _GEN_4448; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4527 = 5'h3 == T_29096 ? T_26182_3_csr_addr : _GEN_4449; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4528 = 5'h3 == T_29096 ? T_26182_3_rob_idx : _GEN_4450; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4529 = 5'h3 == T_29096 ? T_26182_3_ldq_idx : _GEN_4451; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4530 = 5'h3 == T_29096 ? T_26182_3_stq_idx : _GEN_4452; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4531 = 5'h3 == T_29096 ? T_26182_3_brob_idx : _GEN_4453; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4532 = 5'h3 == T_29096 ? T_26182_3_pdst : _GEN_4454; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4533 = 5'h3 == T_29096 ? T_26182_3_pop1 : _GEN_4455; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4534 = 5'h3 == T_29096 ? T_26182_3_pop2 : _GEN_4456; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4535 = 5'h3 == T_29096 ? T_26182_3_pop3 : _GEN_4457; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4536 = 5'h3 == T_29096 ? T_26182_3_prs1_busy : _GEN_4458; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4537 = 5'h3 == T_29096 ? T_26182_3_prs2_busy : _GEN_4459; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4538 = 5'h3 == T_29096 ? T_26182_3_prs3_busy : _GEN_4460; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4539 = 5'h3 == T_29096 ? T_26182_3_stale_pdst : _GEN_4461; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4540 = 5'h3 == T_29096 ? T_26182_3_exception : _GEN_4462; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4541 = 5'h3 == T_29096 ? T_26182_3_exc_cause : _GEN_4463; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4542 = 5'h3 == T_29096 ? T_26182_3_bypassable : _GEN_4464; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4543 = 5'h3 == T_29096 ? T_26182_3_mem_cmd : _GEN_4465; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4544 = 5'h3 == T_29096 ? T_26182_3_mem_typ : _GEN_4466; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4545 = 5'h3 == T_29096 ? T_26182_3_is_fence : _GEN_4467; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4546 = 5'h3 == T_29096 ? T_26182_3_is_fencei : _GEN_4468; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4547 = 5'h3 == T_29096 ? T_26182_3_is_store : _GEN_4469; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4548 = 5'h3 == T_29096 ? T_26182_3_is_amo : _GEN_4470; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4549 = 5'h3 == T_29096 ? T_26182_3_is_load : _GEN_4471; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4550 = 5'h3 == T_29096 ? T_26182_3_is_unique : _GEN_4472; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4551 = 5'h3 == T_29096 ? T_26182_3_flush_on_commit : _GEN_4473; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4552 = 5'h3 == T_29096 ? T_26182_3_ldst : _GEN_4474; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4553 = 5'h3 == T_29096 ? T_26182_3_lrs1 : _GEN_4475; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4554 = 5'h3 == T_29096 ? T_26182_3_lrs2 : _GEN_4476; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4555 = 5'h3 == T_29096 ? T_26182_3_lrs3 : _GEN_4477; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4556 = 5'h3 == T_29096 ? T_26182_3_ldst_val : _GEN_4478; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4557 = 5'h3 == T_29096 ? T_26182_3_dst_rtype : _GEN_4479; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4558 = 5'h3 == T_29096 ? T_26182_3_lrs1_rtype : _GEN_4480; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4559 = 5'h3 == T_29096 ? T_26182_3_lrs2_rtype : _GEN_4481; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4560 = 5'h3 == T_29096 ? T_26182_3_frs3_en : _GEN_4482; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4561 = 5'h3 == T_29096 ? T_26182_3_fp_val : _GEN_4483; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4562 = 5'h3 == T_29096 ? T_26182_3_fp_single : _GEN_4484; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4563 = 5'h3 == T_29096 ? T_26182_3_xcpt_if : _GEN_4485; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4564 = 5'h3 == T_29096 ? T_26182_3_replay_if : _GEN_4486; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4566 = 5'h3 == T_29096 ? T_26182_3_debug_events_fetch_seq : _GEN_4488; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4567 = 5'h4 == T_29096 ? T_26182_4_valid : _GEN_4489; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4568 = 5'h4 == T_29096 ? T_26182_4_iw_state : _GEN_4490; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4569 = 5'h4 == T_29096 ? T_26182_4_uopc : _GEN_4491; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4570 = 5'h4 == T_29096 ? T_26182_4_inst : _GEN_4492; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4571 = 5'h4 == T_29096 ? T_26182_4_pc : _GEN_4493; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4572 = 5'h4 == T_29096 ? T_26182_4_fu_code : _GEN_4494; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4573 = 5'h4 == T_29096 ? T_26182_4_ctrl_br_type : _GEN_4495; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4574 = 5'h4 == T_29096 ? T_26182_4_ctrl_op1_sel : _GEN_4496; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4575 = 5'h4 == T_29096 ? T_26182_4_ctrl_op2_sel : _GEN_4497; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4576 = 5'h4 == T_29096 ? T_26182_4_ctrl_imm_sel : _GEN_4498; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4577 = 5'h4 == T_29096 ? T_26182_4_ctrl_op_fcn : _GEN_4499; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4578 = 5'h4 == T_29096 ? T_26182_4_ctrl_fcn_dw : _GEN_4500; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4579 = 5'h4 == T_29096 ? T_26182_4_ctrl_rf_wen : _GEN_4501; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4580 = 5'h4 == T_29096 ? T_26182_4_ctrl_csr_cmd : _GEN_4502; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4581 = 5'h4 == T_29096 ? T_26182_4_ctrl_is_load : _GEN_4503; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4582 = 5'h4 == T_29096 ? T_26182_4_ctrl_is_sta : _GEN_4504; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4583 = 5'h4 == T_29096 ? T_26182_4_ctrl_is_std : _GEN_4505; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4584 = 5'h4 == T_29096 ? T_26182_4_wakeup_delay : _GEN_4506; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4585 = 5'h4 == T_29096 ? T_26182_4_allocate_brtag : _GEN_4507; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4586 = 5'h4 == T_29096 ? T_26182_4_is_br_or_jmp : _GEN_4508; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4587 = 5'h4 == T_29096 ? T_26182_4_is_jump : _GEN_4509; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4588 = 5'h4 == T_29096 ? T_26182_4_is_jal : _GEN_4510; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4589 = 5'h4 == T_29096 ? T_26182_4_is_ret : _GEN_4511; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4590 = 5'h4 == T_29096 ? T_26182_4_is_call : _GEN_4512; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4591 = 5'h4 == T_29096 ? T_26182_4_br_mask : _GEN_4513; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4592 = 5'h4 == T_29096 ? T_26182_4_br_tag : _GEN_4514; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4593 = 5'h4 == T_29096 ? T_26182_4_br_prediction_bpd_predict_val : _GEN_4515; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4594 = 5'h4 == T_29096 ? T_26182_4_br_prediction_bpd_predict_taken : _GEN_4516; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4595 = 5'h4 == T_29096 ? T_26182_4_br_prediction_btb_hit : _GEN_4517; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4596 = 5'h4 == T_29096 ? T_26182_4_br_prediction_btb_predicted : _GEN_4518; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4597 = 5'h4 == T_29096 ? T_26182_4_br_prediction_is_br_or_jalr : _GEN_4519; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4598 = 5'h4 == T_29096 ? T_26182_4_stat_brjmp_mispredicted : _GEN_4520; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4599 = 5'h4 == T_29096 ? T_26182_4_stat_btb_made_pred : _GEN_4521; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4600 = 5'h4 == T_29096 ? T_26182_4_stat_btb_mispredicted : _GEN_4522; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4601 = 5'h4 == T_29096 ? T_26182_4_stat_bpd_made_pred : _GEN_4523; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4602 = 5'h4 == T_29096 ? T_26182_4_stat_bpd_mispredicted : _GEN_4524; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4603 = 5'h4 == T_29096 ? T_26182_4_fetch_pc_lob : _GEN_4525; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4604 = 5'h4 == T_29096 ? T_26182_4_imm_packed : _GEN_4526; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4605 = 5'h4 == T_29096 ? T_26182_4_csr_addr : _GEN_4527; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4606 = 5'h4 == T_29096 ? T_26182_4_rob_idx : _GEN_4528; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4607 = 5'h4 == T_29096 ? T_26182_4_ldq_idx : _GEN_4529; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4608 = 5'h4 == T_29096 ? T_26182_4_stq_idx : _GEN_4530; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4609 = 5'h4 == T_29096 ? T_26182_4_brob_idx : _GEN_4531; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4610 = 5'h4 == T_29096 ? T_26182_4_pdst : _GEN_4532; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4611 = 5'h4 == T_29096 ? T_26182_4_pop1 : _GEN_4533; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4612 = 5'h4 == T_29096 ? T_26182_4_pop2 : _GEN_4534; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4613 = 5'h4 == T_29096 ? T_26182_4_pop3 : _GEN_4535; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4614 = 5'h4 == T_29096 ? T_26182_4_prs1_busy : _GEN_4536; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4615 = 5'h4 == T_29096 ? T_26182_4_prs2_busy : _GEN_4537; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4616 = 5'h4 == T_29096 ? T_26182_4_prs3_busy : _GEN_4538; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4617 = 5'h4 == T_29096 ? T_26182_4_stale_pdst : _GEN_4539; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4618 = 5'h4 == T_29096 ? T_26182_4_exception : _GEN_4540; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4619 = 5'h4 == T_29096 ? T_26182_4_exc_cause : _GEN_4541; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4620 = 5'h4 == T_29096 ? T_26182_4_bypassable : _GEN_4542; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4621 = 5'h4 == T_29096 ? T_26182_4_mem_cmd : _GEN_4543; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4622 = 5'h4 == T_29096 ? T_26182_4_mem_typ : _GEN_4544; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4623 = 5'h4 == T_29096 ? T_26182_4_is_fence : _GEN_4545; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4624 = 5'h4 == T_29096 ? T_26182_4_is_fencei : _GEN_4546; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4625 = 5'h4 == T_29096 ? T_26182_4_is_store : _GEN_4547; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4626 = 5'h4 == T_29096 ? T_26182_4_is_amo : _GEN_4548; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4627 = 5'h4 == T_29096 ? T_26182_4_is_load : _GEN_4549; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4628 = 5'h4 == T_29096 ? T_26182_4_is_unique : _GEN_4550; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4629 = 5'h4 == T_29096 ? T_26182_4_flush_on_commit : _GEN_4551; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4630 = 5'h4 == T_29096 ? T_26182_4_ldst : _GEN_4552; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4631 = 5'h4 == T_29096 ? T_26182_4_lrs1 : _GEN_4553; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4632 = 5'h4 == T_29096 ? T_26182_4_lrs2 : _GEN_4554; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4633 = 5'h4 == T_29096 ? T_26182_4_lrs3 : _GEN_4555; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4634 = 5'h4 == T_29096 ? T_26182_4_ldst_val : _GEN_4556; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4635 = 5'h4 == T_29096 ? T_26182_4_dst_rtype : _GEN_4557; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4636 = 5'h4 == T_29096 ? T_26182_4_lrs1_rtype : _GEN_4558; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4637 = 5'h4 == T_29096 ? T_26182_4_lrs2_rtype : _GEN_4559; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4638 = 5'h4 == T_29096 ? T_26182_4_frs3_en : _GEN_4560; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4639 = 5'h4 == T_29096 ? T_26182_4_fp_val : _GEN_4561; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4640 = 5'h4 == T_29096 ? T_26182_4_fp_single : _GEN_4562; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4641 = 5'h4 == T_29096 ? T_26182_4_xcpt_if : _GEN_4563; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4642 = 5'h4 == T_29096 ? T_26182_4_replay_if : _GEN_4564; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4644 = 5'h4 == T_29096 ? T_26182_4_debug_events_fetch_seq : _GEN_4566; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4645 = 5'h5 == T_29096 ? T_26182_5_valid : _GEN_4567; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4646 = 5'h5 == T_29096 ? T_26182_5_iw_state : _GEN_4568; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4647 = 5'h5 == T_29096 ? T_26182_5_uopc : _GEN_4569; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4648 = 5'h5 == T_29096 ? T_26182_5_inst : _GEN_4570; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4649 = 5'h5 == T_29096 ? T_26182_5_pc : _GEN_4571; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4650 = 5'h5 == T_29096 ? T_26182_5_fu_code : _GEN_4572; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4651 = 5'h5 == T_29096 ? T_26182_5_ctrl_br_type : _GEN_4573; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4652 = 5'h5 == T_29096 ? T_26182_5_ctrl_op1_sel : _GEN_4574; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4653 = 5'h5 == T_29096 ? T_26182_5_ctrl_op2_sel : _GEN_4575; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4654 = 5'h5 == T_29096 ? T_26182_5_ctrl_imm_sel : _GEN_4576; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4655 = 5'h5 == T_29096 ? T_26182_5_ctrl_op_fcn : _GEN_4577; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4656 = 5'h5 == T_29096 ? T_26182_5_ctrl_fcn_dw : _GEN_4578; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4657 = 5'h5 == T_29096 ? T_26182_5_ctrl_rf_wen : _GEN_4579; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4658 = 5'h5 == T_29096 ? T_26182_5_ctrl_csr_cmd : _GEN_4580; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4659 = 5'h5 == T_29096 ? T_26182_5_ctrl_is_load : _GEN_4581; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4660 = 5'h5 == T_29096 ? T_26182_5_ctrl_is_sta : _GEN_4582; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4661 = 5'h5 == T_29096 ? T_26182_5_ctrl_is_std : _GEN_4583; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4662 = 5'h5 == T_29096 ? T_26182_5_wakeup_delay : _GEN_4584; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4663 = 5'h5 == T_29096 ? T_26182_5_allocate_brtag : _GEN_4585; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4664 = 5'h5 == T_29096 ? T_26182_5_is_br_or_jmp : _GEN_4586; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4665 = 5'h5 == T_29096 ? T_26182_5_is_jump : _GEN_4587; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4666 = 5'h5 == T_29096 ? T_26182_5_is_jal : _GEN_4588; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4667 = 5'h5 == T_29096 ? T_26182_5_is_ret : _GEN_4589; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4668 = 5'h5 == T_29096 ? T_26182_5_is_call : _GEN_4590; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4669 = 5'h5 == T_29096 ? T_26182_5_br_mask : _GEN_4591; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4670 = 5'h5 == T_29096 ? T_26182_5_br_tag : _GEN_4592; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4671 = 5'h5 == T_29096 ? T_26182_5_br_prediction_bpd_predict_val : _GEN_4593; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4672 = 5'h5 == T_29096 ? T_26182_5_br_prediction_bpd_predict_taken : _GEN_4594; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4673 = 5'h5 == T_29096 ? T_26182_5_br_prediction_btb_hit : _GEN_4595; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4674 = 5'h5 == T_29096 ? T_26182_5_br_prediction_btb_predicted : _GEN_4596; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4675 = 5'h5 == T_29096 ? T_26182_5_br_prediction_is_br_or_jalr : _GEN_4597; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4676 = 5'h5 == T_29096 ? T_26182_5_stat_brjmp_mispredicted : _GEN_4598; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4677 = 5'h5 == T_29096 ? T_26182_5_stat_btb_made_pred : _GEN_4599; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4678 = 5'h5 == T_29096 ? T_26182_5_stat_btb_mispredicted : _GEN_4600; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4679 = 5'h5 == T_29096 ? T_26182_5_stat_bpd_made_pred : _GEN_4601; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4680 = 5'h5 == T_29096 ? T_26182_5_stat_bpd_mispredicted : _GEN_4602; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4681 = 5'h5 == T_29096 ? T_26182_5_fetch_pc_lob : _GEN_4603; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4682 = 5'h5 == T_29096 ? T_26182_5_imm_packed : _GEN_4604; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4683 = 5'h5 == T_29096 ? T_26182_5_csr_addr : _GEN_4605; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4684 = 5'h5 == T_29096 ? T_26182_5_rob_idx : _GEN_4606; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4685 = 5'h5 == T_29096 ? T_26182_5_ldq_idx : _GEN_4607; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4686 = 5'h5 == T_29096 ? T_26182_5_stq_idx : _GEN_4608; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4687 = 5'h5 == T_29096 ? T_26182_5_brob_idx : _GEN_4609; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4688 = 5'h5 == T_29096 ? T_26182_5_pdst : _GEN_4610; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4689 = 5'h5 == T_29096 ? T_26182_5_pop1 : _GEN_4611; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4690 = 5'h5 == T_29096 ? T_26182_5_pop2 : _GEN_4612; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4691 = 5'h5 == T_29096 ? T_26182_5_pop3 : _GEN_4613; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4692 = 5'h5 == T_29096 ? T_26182_5_prs1_busy : _GEN_4614; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4693 = 5'h5 == T_29096 ? T_26182_5_prs2_busy : _GEN_4615; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4694 = 5'h5 == T_29096 ? T_26182_5_prs3_busy : _GEN_4616; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4695 = 5'h5 == T_29096 ? T_26182_5_stale_pdst : _GEN_4617; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4696 = 5'h5 == T_29096 ? T_26182_5_exception : _GEN_4618; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4697 = 5'h5 == T_29096 ? T_26182_5_exc_cause : _GEN_4619; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4698 = 5'h5 == T_29096 ? T_26182_5_bypassable : _GEN_4620; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4699 = 5'h5 == T_29096 ? T_26182_5_mem_cmd : _GEN_4621; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4700 = 5'h5 == T_29096 ? T_26182_5_mem_typ : _GEN_4622; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4701 = 5'h5 == T_29096 ? T_26182_5_is_fence : _GEN_4623; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4702 = 5'h5 == T_29096 ? T_26182_5_is_fencei : _GEN_4624; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4703 = 5'h5 == T_29096 ? T_26182_5_is_store : _GEN_4625; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4704 = 5'h5 == T_29096 ? T_26182_5_is_amo : _GEN_4626; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4705 = 5'h5 == T_29096 ? T_26182_5_is_load : _GEN_4627; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4706 = 5'h5 == T_29096 ? T_26182_5_is_unique : _GEN_4628; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4707 = 5'h5 == T_29096 ? T_26182_5_flush_on_commit : _GEN_4629; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4708 = 5'h5 == T_29096 ? T_26182_5_ldst : _GEN_4630; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4709 = 5'h5 == T_29096 ? T_26182_5_lrs1 : _GEN_4631; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4710 = 5'h5 == T_29096 ? T_26182_5_lrs2 : _GEN_4632; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4711 = 5'h5 == T_29096 ? T_26182_5_lrs3 : _GEN_4633; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4712 = 5'h5 == T_29096 ? T_26182_5_ldst_val : _GEN_4634; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4713 = 5'h5 == T_29096 ? T_26182_5_dst_rtype : _GEN_4635; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4714 = 5'h5 == T_29096 ? T_26182_5_lrs1_rtype : _GEN_4636; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4715 = 5'h5 == T_29096 ? T_26182_5_lrs2_rtype : _GEN_4637; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4716 = 5'h5 == T_29096 ? T_26182_5_frs3_en : _GEN_4638; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4717 = 5'h5 == T_29096 ? T_26182_5_fp_val : _GEN_4639; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4718 = 5'h5 == T_29096 ? T_26182_5_fp_single : _GEN_4640; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4719 = 5'h5 == T_29096 ? T_26182_5_xcpt_if : _GEN_4641; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4720 = 5'h5 == T_29096 ? T_26182_5_replay_if : _GEN_4642; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4722 = 5'h5 == T_29096 ? T_26182_5_debug_events_fetch_seq : _GEN_4644; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4723 = 5'h6 == T_29096 ? T_26182_6_valid : _GEN_4645; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4724 = 5'h6 == T_29096 ? T_26182_6_iw_state : _GEN_4646; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4725 = 5'h6 == T_29096 ? T_26182_6_uopc : _GEN_4647; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4726 = 5'h6 == T_29096 ? T_26182_6_inst : _GEN_4648; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4727 = 5'h6 == T_29096 ? T_26182_6_pc : _GEN_4649; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4728 = 5'h6 == T_29096 ? T_26182_6_fu_code : _GEN_4650; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4729 = 5'h6 == T_29096 ? T_26182_6_ctrl_br_type : _GEN_4651; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4730 = 5'h6 == T_29096 ? T_26182_6_ctrl_op1_sel : _GEN_4652; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4731 = 5'h6 == T_29096 ? T_26182_6_ctrl_op2_sel : _GEN_4653; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4732 = 5'h6 == T_29096 ? T_26182_6_ctrl_imm_sel : _GEN_4654; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4733 = 5'h6 == T_29096 ? T_26182_6_ctrl_op_fcn : _GEN_4655; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4734 = 5'h6 == T_29096 ? T_26182_6_ctrl_fcn_dw : _GEN_4656; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4735 = 5'h6 == T_29096 ? T_26182_6_ctrl_rf_wen : _GEN_4657; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4736 = 5'h6 == T_29096 ? T_26182_6_ctrl_csr_cmd : _GEN_4658; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4737 = 5'h6 == T_29096 ? T_26182_6_ctrl_is_load : _GEN_4659; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4738 = 5'h6 == T_29096 ? T_26182_6_ctrl_is_sta : _GEN_4660; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4739 = 5'h6 == T_29096 ? T_26182_6_ctrl_is_std : _GEN_4661; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4740 = 5'h6 == T_29096 ? T_26182_6_wakeup_delay : _GEN_4662; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4741 = 5'h6 == T_29096 ? T_26182_6_allocate_brtag : _GEN_4663; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4742 = 5'h6 == T_29096 ? T_26182_6_is_br_or_jmp : _GEN_4664; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4743 = 5'h6 == T_29096 ? T_26182_6_is_jump : _GEN_4665; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4744 = 5'h6 == T_29096 ? T_26182_6_is_jal : _GEN_4666; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4745 = 5'h6 == T_29096 ? T_26182_6_is_ret : _GEN_4667; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4746 = 5'h6 == T_29096 ? T_26182_6_is_call : _GEN_4668; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4747 = 5'h6 == T_29096 ? T_26182_6_br_mask : _GEN_4669; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4748 = 5'h6 == T_29096 ? T_26182_6_br_tag : _GEN_4670; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4749 = 5'h6 == T_29096 ? T_26182_6_br_prediction_bpd_predict_val : _GEN_4671; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4750 = 5'h6 == T_29096 ? T_26182_6_br_prediction_bpd_predict_taken : _GEN_4672; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4751 = 5'h6 == T_29096 ? T_26182_6_br_prediction_btb_hit : _GEN_4673; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4752 = 5'h6 == T_29096 ? T_26182_6_br_prediction_btb_predicted : _GEN_4674; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4753 = 5'h6 == T_29096 ? T_26182_6_br_prediction_is_br_or_jalr : _GEN_4675; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4754 = 5'h6 == T_29096 ? T_26182_6_stat_brjmp_mispredicted : _GEN_4676; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4755 = 5'h6 == T_29096 ? T_26182_6_stat_btb_made_pred : _GEN_4677; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4756 = 5'h6 == T_29096 ? T_26182_6_stat_btb_mispredicted : _GEN_4678; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4757 = 5'h6 == T_29096 ? T_26182_6_stat_bpd_made_pred : _GEN_4679; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4758 = 5'h6 == T_29096 ? T_26182_6_stat_bpd_mispredicted : _GEN_4680; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4759 = 5'h6 == T_29096 ? T_26182_6_fetch_pc_lob : _GEN_4681; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4760 = 5'h6 == T_29096 ? T_26182_6_imm_packed : _GEN_4682; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4761 = 5'h6 == T_29096 ? T_26182_6_csr_addr : _GEN_4683; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4762 = 5'h6 == T_29096 ? T_26182_6_rob_idx : _GEN_4684; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4763 = 5'h6 == T_29096 ? T_26182_6_ldq_idx : _GEN_4685; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4764 = 5'h6 == T_29096 ? T_26182_6_stq_idx : _GEN_4686; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4765 = 5'h6 == T_29096 ? T_26182_6_brob_idx : _GEN_4687; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4766 = 5'h6 == T_29096 ? T_26182_6_pdst : _GEN_4688; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4767 = 5'h6 == T_29096 ? T_26182_6_pop1 : _GEN_4689; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4768 = 5'h6 == T_29096 ? T_26182_6_pop2 : _GEN_4690; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4769 = 5'h6 == T_29096 ? T_26182_6_pop3 : _GEN_4691; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4770 = 5'h6 == T_29096 ? T_26182_6_prs1_busy : _GEN_4692; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4771 = 5'h6 == T_29096 ? T_26182_6_prs2_busy : _GEN_4693; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4772 = 5'h6 == T_29096 ? T_26182_6_prs3_busy : _GEN_4694; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4773 = 5'h6 == T_29096 ? T_26182_6_stale_pdst : _GEN_4695; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4774 = 5'h6 == T_29096 ? T_26182_6_exception : _GEN_4696; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4775 = 5'h6 == T_29096 ? T_26182_6_exc_cause : _GEN_4697; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4776 = 5'h6 == T_29096 ? T_26182_6_bypassable : _GEN_4698; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4777 = 5'h6 == T_29096 ? T_26182_6_mem_cmd : _GEN_4699; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4778 = 5'h6 == T_29096 ? T_26182_6_mem_typ : _GEN_4700; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4779 = 5'h6 == T_29096 ? T_26182_6_is_fence : _GEN_4701; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4780 = 5'h6 == T_29096 ? T_26182_6_is_fencei : _GEN_4702; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4781 = 5'h6 == T_29096 ? T_26182_6_is_store : _GEN_4703; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4782 = 5'h6 == T_29096 ? T_26182_6_is_amo : _GEN_4704; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4783 = 5'h6 == T_29096 ? T_26182_6_is_load : _GEN_4705; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4784 = 5'h6 == T_29096 ? T_26182_6_is_unique : _GEN_4706; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4785 = 5'h6 == T_29096 ? T_26182_6_flush_on_commit : _GEN_4707; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4786 = 5'h6 == T_29096 ? T_26182_6_ldst : _GEN_4708; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4787 = 5'h6 == T_29096 ? T_26182_6_lrs1 : _GEN_4709; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4788 = 5'h6 == T_29096 ? T_26182_6_lrs2 : _GEN_4710; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4789 = 5'h6 == T_29096 ? T_26182_6_lrs3 : _GEN_4711; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4790 = 5'h6 == T_29096 ? T_26182_6_ldst_val : _GEN_4712; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4791 = 5'h6 == T_29096 ? T_26182_6_dst_rtype : _GEN_4713; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4792 = 5'h6 == T_29096 ? T_26182_6_lrs1_rtype : _GEN_4714; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4793 = 5'h6 == T_29096 ? T_26182_6_lrs2_rtype : _GEN_4715; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4794 = 5'h6 == T_29096 ? T_26182_6_frs3_en : _GEN_4716; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4795 = 5'h6 == T_29096 ? T_26182_6_fp_val : _GEN_4717; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4796 = 5'h6 == T_29096 ? T_26182_6_fp_single : _GEN_4718; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4797 = 5'h6 == T_29096 ? T_26182_6_xcpt_if : _GEN_4719; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4798 = 5'h6 == T_29096 ? T_26182_6_replay_if : _GEN_4720; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4800 = 5'h6 == T_29096 ? T_26182_6_debug_events_fetch_seq : _GEN_4722; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4801 = 5'h7 == T_29096 ? T_26182_7_valid : _GEN_4723; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4802 = 5'h7 == T_29096 ? T_26182_7_iw_state : _GEN_4724; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4803 = 5'h7 == T_29096 ? T_26182_7_uopc : _GEN_4725; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4804 = 5'h7 == T_29096 ? T_26182_7_inst : _GEN_4726; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4805 = 5'h7 == T_29096 ? T_26182_7_pc : _GEN_4727; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4806 = 5'h7 == T_29096 ? T_26182_7_fu_code : _GEN_4728; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4807 = 5'h7 == T_29096 ? T_26182_7_ctrl_br_type : _GEN_4729; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4808 = 5'h7 == T_29096 ? T_26182_7_ctrl_op1_sel : _GEN_4730; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4809 = 5'h7 == T_29096 ? T_26182_7_ctrl_op2_sel : _GEN_4731; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4810 = 5'h7 == T_29096 ? T_26182_7_ctrl_imm_sel : _GEN_4732; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4811 = 5'h7 == T_29096 ? T_26182_7_ctrl_op_fcn : _GEN_4733; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4812 = 5'h7 == T_29096 ? T_26182_7_ctrl_fcn_dw : _GEN_4734; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4813 = 5'h7 == T_29096 ? T_26182_7_ctrl_rf_wen : _GEN_4735; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4814 = 5'h7 == T_29096 ? T_26182_7_ctrl_csr_cmd : _GEN_4736; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4815 = 5'h7 == T_29096 ? T_26182_7_ctrl_is_load : _GEN_4737; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4816 = 5'h7 == T_29096 ? T_26182_7_ctrl_is_sta : _GEN_4738; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4817 = 5'h7 == T_29096 ? T_26182_7_ctrl_is_std : _GEN_4739; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4818 = 5'h7 == T_29096 ? T_26182_7_wakeup_delay : _GEN_4740; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4819 = 5'h7 == T_29096 ? T_26182_7_allocate_brtag : _GEN_4741; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4820 = 5'h7 == T_29096 ? T_26182_7_is_br_or_jmp : _GEN_4742; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4821 = 5'h7 == T_29096 ? T_26182_7_is_jump : _GEN_4743; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4822 = 5'h7 == T_29096 ? T_26182_7_is_jal : _GEN_4744; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4823 = 5'h7 == T_29096 ? T_26182_7_is_ret : _GEN_4745; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4824 = 5'h7 == T_29096 ? T_26182_7_is_call : _GEN_4746; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4825 = 5'h7 == T_29096 ? T_26182_7_br_mask : _GEN_4747; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4826 = 5'h7 == T_29096 ? T_26182_7_br_tag : _GEN_4748; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4827 = 5'h7 == T_29096 ? T_26182_7_br_prediction_bpd_predict_val : _GEN_4749; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4828 = 5'h7 == T_29096 ? T_26182_7_br_prediction_bpd_predict_taken : _GEN_4750; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4829 = 5'h7 == T_29096 ? T_26182_7_br_prediction_btb_hit : _GEN_4751; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4830 = 5'h7 == T_29096 ? T_26182_7_br_prediction_btb_predicted : _GEN_4752; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4831 = 5'h7 == T_29096 ? T_26182_7_br_prediction_is_br_or_jalr : _GEN_4753; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4832 = 5'h7 == T_29096 ? T_26182_7_stat_brjmp_mispredicted : _GEN_4754; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4833 = 5'h7 == T_29096 ? T_26182_7_stat_btb_made_pred : _GEN_4755; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4834 = 5'h7 == T_29096 ? T_26182_7_stat_btb_mispredicted : _GEN_4756; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4835 = 5'h7 == T_29096 ? T_26182_7_stat_bpd_made_pred : _GEN_4757; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4836 = 5'h7 == T_29096 ? T_26182_7_stat_bpd_mispredicted : _GEN_4758; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4837 = 5'h7 == T_29096 ? T_26182_7_fetch_pc_lob : _GEN_4759; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4838 = 5'h7 == T_29096 ? T_26182_7_imm_packed : _GEN_4760; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4839 = 5'h7 == T_29096 ? T_26182_7_csr_addr : _GEN_4761; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4840 = 5'h7 == T_29096 ? T_26182_7_rob_idx : _GEN_4762; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4841 = 5'h7 == T_29096 ? T_26182_7_ldq_idx : _GEN_4763; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4842 = 5'h7 == T_29096 ? T_26182_7_stq_idx : _GEN_4764; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4843 = 5'h7 == T_29096 ? T_26182_7_brob_idx : _GEN_4765; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4844 = 5'h7 == T_29096 ? T_26182_7_pdst : _GEN_4766; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4845 = 5'h7 == T_29096 ? T_26182_7_pop1 : _GEN_4767; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4846 = 5'h7 == T_29096 ? T_26182_7_pop2 : _GEN_4768; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4847 = 5'h7 == T_29096 ? T_26182_7_pop3 : _GEN_4769; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4848 = 5'h7 == T_29096 ? T_26182_7_prs1_busy : _GEN_4770; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4849 = 5'h7 == T_29096 ? T_26182_7_prs2_busy : _GEN_4771; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4850 = 5'h7 == T_29096 ? T_26182_7_prs3_busy : _GEN_4772; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4851 = 5'h7 == T_29096 ? T_26182_7_stale_pdst : _GEN_4773; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4852 = 5'h7 == T_29096 ? T_26182_7_exception : _GEN_4774; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4853 = 5'h7 == T_29096 ? T_26182_7_exc_cause : _GEN_4775; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4854 = 5'h7 == T_29096 ? T_26182_7_bypassable : _GEN_4776; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4855 = 5'h7 == T_29096 ? T_26182_7_mem_cmd : _GEN_4777; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4856 = 5'h7 == T_29096 ? T_26182_7_mem_typ : _GEN_4778; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4857 = 5'h7 == T_29096 ? T_26182_7_is_fence : _GEN_4779; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4858 = 5'h7 == T_29096 ? T_26182_7_is_fencei : _GEN_4780; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4859 = 5'h7 == T_29096 ? T_26182_7_is_store : _GEN_4781; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4860 = 5'h7 == T_29096 ? T_26182_7_is_amo : _GEN_4782; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4861 = 5'h7 == T_29096 ? T_26182_7_is_load : _GEN_4783; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4862 = 5'h7 == T_29096 ? T_26182_7_is_unique : _GEN_4784; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4863 = 5'h7 == T_29096 ? T_26182_7_flush_on_commit : _GEN_4785; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4864 = 5'h7 == T_29096 ? T_26182_7_ldst : _GEN_4786; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4865 = 5'h7 == T_29096 ? T_26182_7_lrs1 : _GEN_4787; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4866 = 5'h7 == T_29096 ? T_26182_7_lrs2 : _GEN_4788; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4867 = 5'h7 == T_29096 ? T_26182_7_lrs3 : _GEN_4789; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4868 = 5'h7 == T_29096 ? T_26182_7_ldst_val : _GEN_4790; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4869 = 5'h7 == T_29096 ? T_26182_7_dst_rtype : _GEN_4791; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4870 = 5'h7 == T_29096 ? T_26182_7_lrs1_rtype : _GEN_4792; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4871 = 5'h7 == T_29096 ? T_26182_7_lrs2_rtype : _GEN_4793; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4872 = 5'h7 == T_29096 ? T_26182_7_frs3_en : _GEN_4794; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4873 = 5'h7 == T_29096 ? T_26182_7_fp_val : _GEN_4795; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4874 = 5'h7 == T_29096 ? T_26182_7_fp_single : _GEN_4796; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4875 = 5'h7 == T_29096 ? T_26182_7_xcpt_if : _GEN_4797; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4876 = 5'h7 == T_29096 ? T_26182_7_replay_if : _GEN_4798; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4878 = 5'h7 == T_29096 ? T_26182_7_debug_events_fetch_seq : _GEN_4800; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4879 = 5'h8 == T_29096 ? T_26182_8_valid : _GEN_4801; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4880 = 5'h8 == T_29096 ? T_26182_8_iw_state : _GEN_4802; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4881 = 5'h8 == T_29096 ? T_26182_8_uopc : _GEN_4803; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4882 = 5'h8 == T_29096 ? T_26182_8_inst : _GEN_4804; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4883 = 5'h8 == T_29096 ? T_26182_8_pc : _GEN_4805; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4884 = 5'h8 == T_29096 ? T_26182_8_fu_code : _GEN_4806; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4885 = 5'h8 == T_29096 ? T_26182_8_ctrl_br_type : _GEN_4807; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4886 = 5'h8 == T_29096 ? T_26182_8_ctrl_op1_sel : _GEN_4808; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4887 = 5'h8 == T_29096 ? T_26182_8_ctrl_op2_sel : _GEN_4809; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4888 = 5'h8 == T_29096 ? T_26182_8_ctrl_imm_sel : _GEN_4810; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4889 = 5'h8 == T_29096 ? T_26182_8_ctrl_op_fcn : _GEN_4811; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4890 = 5'h8 == T_29096 ? T_26182_8_ctrl_fcn_dw : _GEN_4812; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4891 = 5'h8 == T_29096 ? T_26182_8_ctrl_rf_wen : _GEN_4813; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4892 = 5'h8 == T_29096 ? T_26182_8_ctrl_csr_cmd : _GEN_4814; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4893 = 5'h8 == T_29096 ? T_26182_8_ctrl_is_load : _GEN_4815; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4894 = 5'h8 == T_29096 ? T_26182_8_ctrl_is_sta : _GEN_4816; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4895 = 5'h8 == T_29096 ? T_26182_8_ctrl_is_std : _GEN_4817; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4896 = 5'h8 == T_29096 ? T_26182_8_wakeup_delay : _GEN_4818; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4897 = 5'h8 == T_29096 ? T_26182_8_allocate_brtag : _GEN_4819; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4898 = 5'h8 == T_29096 ? T_26182_8_is_br_or_jmp : _GEN_4820; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4899 = 5'h8 == T_29096 ? T_26182_8_is_jump : _GEN_4821; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4900 = 5'h8 == T_29096 ? T_26182_8_is_jal : _GEN_4822; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4901 = 5'h8 == T_29096 ? T_26182_8_is_ret : _GEN_4823; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4902 = 5'h8 == T_29096 ? T_26182_8_is_call : _GEN_4824; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4903 = 5'h8 == T_29096 ? T_26182_8_br_mask : _GEN_4825; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4904 = 5'h8 == T_29096 ? T_26182_8_br_tag : _GEN_4826; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4905 = 5'h8 == T_29096 ? T_26182_8_br_prediction_bpd_predict_val : _GEN_4827; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4906 = 5'h8 == T_29096 ? T_26182_8_br_prediction_bpd_predict_taken : _GEN_4828; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4907 = 5'h8 == T_29096 ? T_26182_8_br_prediction_btb_hit : _GEN_4829; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4908 = 5'h8 == T_29096 ? T_26182_8_br_prediction_btb_predicted : _GEN_4830; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4909 = 5'h8 == T_29096 ? T_26182_8_br_prediction_is_br_or_jalr : _GEN_4831; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4910 = 5'h8 == T_29096 ? T_26182_8_stat_brjmp_mispredicted : _GEN_4832; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4911 = 5'h8 == T_29096 ? T_26182_8_stat_btb_made_pred : _GEN_4833; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4912 = 5'h8 == T_29096 ? T_26182_8_stat_btb_mispredicted : _GEN_4834; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4913 = 5'h8 == T_29096 ? T_26182_8_stat_bpd_made_pred : _GEN_4835; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4914 = 5'h8 == T_29096 ? T_26182_8_stat_bpd_mispredicted : _GEN_4836; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4915 = 5'h8 == T_29096 ? T_26182_8_fetch_pc_lob : _GEN_4837; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4916 = 5'h8 == T_29096 ? T_26182_8_imm_packed : _GEN_4838; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4917 = 5'h8 == T_29096 ? T_26182_8_csr_addr : _GEN_4839; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4918 = 5'h8 == T_29096 ? T_26182_8_rob_idx : _GEN_4840; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4919 = 5'h8 == T_29096 ? T_26182_8_ldq_idx : _GEN_4841; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4920 = 5'h8 == T_29096 ? T_26182_8_stq_idx : _GEN_4842; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4921 = 5'h8 == T_29096 ? T_26182_8_brob_idx : _GEN_4843; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4922 = 5'h8 == T_29096 ? T_26182_8_pdst : _GEN_4844; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4923 = 5'h8 == T_29096 ? T_26182_8_pop1 : _GEN_4845; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4924 = 5'h8 == T_29096 ? T_26182_8_pop2 : _GEN_4846; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4925 = 5'h8 == T_29096 ? T_26182_8_pop3 : _GEN_4847; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4926 = 5'h8 == T_29096 ? T_26182_8_prs1_busy : _GEN_4848; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4927 = 5'h8 == T_29096 ? T_26182_8_prs2_busy : _GEN_4849; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4928 = 5'h8 == T_29096 ? T_26182_8_prs3_busy : _GEN_4850; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_4929 = 5'h8 == T_29096 ? T_26182_8_stale_pdst : _GEN_4851; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4930 = 5'h8 == T_29096 ? T_26182_8_exception : _GEN_4852; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_4931 = 5'h8 == T_29096 ? T_26182_8_exc_cause : _GEN_4853; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4932 = 5'h8 == T_29096 ? T_26182_8_bypassable : _GEN_4854; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4933 = 5'h8 == T_29096 ? T_26182_8_mem_cmd : _GEN_4855; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4934 = 5'h8 == T_29096 ? T_26182_8_mem_typ : _GEN_4856; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4935 = 5'h8 == T_29096 ? T_26182_8_is_fence : _GEN_4857; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4936 = 5'h8 == T_29096 ? T_26182_8_is_fencei : _GEN_4858; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4937 = 5'h8 == T_29096 ? T_26182_8_is_store : _GEN_4859; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4938 = 5'h8 == T_29096 ? T_26182_8_is_amo : _GEN_4860; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4939 = 5'h8 == T_29096 ? T_26182_8_is_load : _GEN_4861; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4940 = 5'h8 == T_29096 ? T_26182_8_is_unique : _GEN_4862; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4941 = 5'h8 == T_29096 ? T_26182_8_flush_on_commit : _GEN_4863; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4942 = 5'h8 == T_29096 ? T_26182_8_ldst : _GEN_4864; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4943 = 5'h8 == T_29096 ? T_26182_8_lrs1 : _GEN_4865; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4944 = 5'h8 == T_29096 ? T_26182_8_lrs2 : _GEN_4866; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4945 = 5'h8 == T_29096 ? T_26182_8_lrs3 : _GEN_4867; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4946 = 5'h8 == T_29096 ? T_26182_8_ldst_val : _GEN_4868; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4947 = 5'h8 == T_29096 ? T_26182_8_dst_rtype : _GEN_4869; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4948 = 5'h8 == T_29096 ? T_26182_8_lrs1_rtype : _GEN_4870; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4949 = 5'h8 == T_29096 ? T_26182_8_lrs2_rtype : _GEN_4871; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4950 = 5'h8 == T_29096 ? T_26182_8_frs3_en : _GEN_4872; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4951 = 5'h8 == T_29096 ? T_26182_8_fp_val : _GEN_4873; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4952 = 5'h8 == T_29096 ? T_26182_8_fp_single : _GEN_4874; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4953 = 5'h8 == T_29096 ? T_26182_8_xcpt_if : _GEN_4875; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4954 = 5'h8 == T_29096 ? T_26182_8_replay_if : _GEN_4876; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4956 = 5'h8 == T_29096 ? T_26182_8_debug_events_fetch_seq : _GEN_4878; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4957 = 5'h9 == T_29096 ? T_26182_9_valid : _GEN_4879; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4958 = 5'h9 == T_29096 ? T_26182_9_iw_state : _GEN_4880; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_4959 = 5'h9 == T_29096 ? T_26182_9_uopc : _GEN_4881; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_4960 = 5'h9 == T_29096 ? T_26182_9_inst : _GEN_4882; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_4961 = 5'h9 == T_29096 ? T_26182_9_pc : _GEN_4883; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4962 = 5'h9 == T_29096 ? T_26182_9_fu_code : _GEN_4884; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4963 = 5'h9 == T_29096 ? T_26182_9_ctrl_br_type : _GEN_4885; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4964 = 5'h9 == T_29096 ? T_26182_9_ctrl_op1_sel : _GEN_4886; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4965 = 5'h9 == T_29096 ? T_26182_9_ctrl_op2_sel : _GEN_4887; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4966 = 5'h9 == T_29096 ? T_26182_9_ctrl_imm_sel : _GEN_4888; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4967 = 5'h9 == T_29096 ? T_26182_9_ctrl_op_fcn : _GEN_4889; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4968 = 5'h9 == T_29096 ? T_26182_9_ctrl_fcn_dw : _GEN_4890; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4969 = 5'h9 == T_29096 ? T_26182_9_ctrl_rf_wen : _GEN_4891; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4970 = 5'h9 == T_29096 ? T_26182_9_ctrl_csr_cmd : _GEN_4892; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4971 = 5'h9 == T_29096 ? T_26182_9_ctrl_is_load : _GEN_4893; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4972 = 5'h9 == T_29096 ? T_26182_9_ctrl_is_sta : _GEN_4894; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4973 = 5'h9 == T_29096 ? T_26182_9_ctrl_is_std : _GEN_4895; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_4974 = 5'h9 == T_29096 ? T_26182_9_wakeup_delay : _GEN_4896; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4975 = 5'h9 == T_29096 ? T_26182_9_allocate_brtag : _GEN_4897; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4976 = 5'h9 == T_29096 ? T_26182_9_is_br_or_jmp : _GEN_4898; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4977 = 5'h9 == T_29096 ? T_26182_9_is_jump : _GEN_4899; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4978 = 5'h9 == T_29096 ? T_26182_9_is_jal : _GEN_4900; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4979 = 5'h9 == T_29096 ? T_26182_9_is_ret : _GEN_4901; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4980 = 5'h9 == T_29096 ? T_26182_9_is_call : _GEN_4902; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_4981 = 5'h9 == T_29096 ? T_26182_9_br_mask : _GEN_4903; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4982 = 5'h9 == T_29096 ? T_26182_9_br_tag : _GEN_4904; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4983 = 5'h9 == T_29096 ? T_26182_9_br_prediction_bpd_predict_val : _GEN_4905; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4984 = 5'h9 == T_29096 ? T_26182_9_br_prediction_bpd_predict_taken : _GEN_4906; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4985 = 5'h9 == T_29096 ? T_26182_9_br_prediction_btb_hit : _GEN_4907; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4986 = 5'h9 == T_29096 ? T_26182_9_br_prediction_btb_predicted : _GEN_4908; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4987 = 5'h9 == T_29096 ? T_26182_9_br_prediction_is_br_or_jalr : _GEN_4909; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4988 = 5'h9 == T_29096 ? T_26182_9_stat_brjmp_mispredicted : _GEN_4910; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4989 = 5'h9 == T_29096 ? T_26182_9_stat_btb_made_pred : _GEN_4911; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4990 = 5'h9 == T_29096 ? T_26182_9_stat_btb_mispredicted : _GEN_4912; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4991 = 5'h9 == T_29096 ? T_26182_9_stat_bpd_made_pred : _GEN_4913; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_4992 = 5'h9 == T_29096 ? T_26182_9_stat_bpd_mispredicted : _GEN_4914; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_4993 = 5'h9 == T_29096 ? T_26182_9_fetch_pc_lob : _GEN_4915; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_4994 = 5'h9 == T_29096 ? T_26182_9_imm_packed : _GEN_4916; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_4995 = 5'h9 == T_29096 ? T_26182_9_csr_addr : _GEN_4917; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_4996 = 5'h9 == T_29096 ? T_26182_9_rob_idx : _GEN_4918; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4997 = 5'h9 == T_29096 ? T_26182_9_ldq_idx : _GEN_4919; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_4998 = 5'h9 == T_29096 ? T_26182_9_stq_idx : _GEN_4920; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_4999 = 5'h9 == T_29096 ? T_26182_9_brob_idx : _GEN_4921; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5000 = 5'h9 == T_29096 ? T_26182_9_pdst : _GEN_4922; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5001 = 5'h9 == T_29096 ? T_26182_9_pop1 : _GEN_4923; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5002 = 5'h9 == T_29096 ? T_26182_9_pop2 : _GEN_4924; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5003 = 5'h9 == T_29096 ? T_26182_9_pop3 : _GEN_4925; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5004 = 5'h9 == T_29096 ? T_26182_9_prs1_busy : _GEN_4926; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5005 = 5'h9 == T_29096 ? T_26182_9_prs2_busy : _GEN_4927; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5006 = 5'h9 == T_29096 ? T_26182_9_prs3_busy : _GEN_4928; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5007 = 5'h9 == T_29096 ? T_26182_9_stale_pdst : _GEN_4929; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5008 = 5'h9 == T_29096 ? T_26182_9_exception : _GEN_4930; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5009 = 5'h9 == T_29096 ? T_26182_9_exc_cause : _GEN_4931; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5010 = 5'h9 == T_29096 ? T_26182_9_bypassable : _GEN_4932; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5011 = 5'h9 == T_29096 ? T_26182_9_mem_cmd : _GEN_4933; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5012 = 5'h9 == T_29096 ? T_26182_9_mem_typ : _GEN_4934; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5013 = 5'h9 == T_29096 ? T_26182_9_is_fence : _GEN_4935; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5014 = 5'h9 == T_29096 ? T_26182_9_is_fencei : _GEN_4936; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5015 = 5'h9 == T_29096 ? T_26182_9_is_store : _GEN_4937; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5016 = 5'h9 == T_29096 ? T_26182_9_is_amo : _GEN_4938; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5017 = 5'h9 == T_29096 ? T_26182_9_is_load : _GEN_4939; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5018 = 5'h9 == T_29096 ? T_26182_9_is_unique : _GEN_4940; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5019 = 5'h9 == T_29096 ? T_26182_9_flush_on_commit : _GEN_4941; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5020 = 5'h9 == T_29096 ? T_26182_9_ldst : _GEN_4942; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5021 = 5'h9 == T_29096 ? T_26182_9_lrs1 : _GEN_4943; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5022 = 5'h9 == T_29096 ? T_26182_9_lrs2 : _GEN_4944; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5023 = 5'h9 == T_29096 ? T_26182_9_lrs3 : _GEN_4945; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5024 = 5'h9 == T_29096 ? T_26182_9_ldst_val : _GEN_4946; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5025 = 5'h9 == T_29096 ? T_26182_9_dst_rtype : _GEN_4947; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5026 = 5'h9 == T_29096 ? T_26182_9_lrs1_rtype : _GEN_4948; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5027 = 5'h9 == T_29096 ? T_26182_9_lrs2_rtype : _GEN_4949; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5028 = 5'h9 == T_29096 ? T_26182_9_frs3_en : _GEN_4950; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5029 = 5'h9 == T_29096 ? T_26182_9_fp_val : _GEN_4951; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5030 = 5'h9 == T_29096 ? T_26182_9_fp_single : _GEN_4952; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5031 = 5'h9 == T_29096 ? T_26182_9_xcpt_if : _GEN_4953; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5032 = 5'h9 == T_29096 ? T_26182_9_replay_if : _GEN_4954; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5034 = 5'h9 == T_29096 ? T_26182_9_debug_events_fetch_seq : _GEN_4956; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5035 = 5'ha == T_29096 ? T_26182_10_valid : _GEN_4957; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5036 = 5'ha == T_29096 ? T_26182_10_iw_state : _GEN_4958; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5037 = 5'ha == T_29096 ? T_26182_10_uopc : _GEN_4959; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5038 = 5'ha == T_29096 ? T_26182_10_inst : _GEN_4960; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5039 = 5'ha == T_29096 ? T_26182_10_pc : _GEN_4961; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5040 = 5'ha == T_29096 ? T_26182_10_fu_code : _GEN_4962; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5041 = 5'ha == T_29096 ? T_26182_10_ctrl_br_type : _GEN_4963; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5042 = 5'ha == T_29096 ? T_26182_10_ctrl_op1_sel : _GEN_4964; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5043 = 5'ha == T_29096 ? T_26182_10_ctrl_op2_sel : _GEN_4965; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5044 = 5'ha == T_29096 ? T_26182_10_ctrl_imm_sel : _GEN_4966; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5045 = 5'ha == T_29096 ? T_26182_10_ctrl_op_fcn : _GEN_4967; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5046 = 5'ha == T_29096 ? T_26182_10_ctrl_fcn_dw : _GEN_4968; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5047 = 5'ha == T_29096 ? T_26182_10_ctrl_rf_wen : _GEN_4969; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5048 = 5'ha == T_29096 ? T_26182_10_ctrl_csr_cmd : _GEN_4970; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5049 = 5'ha == T_29096 ? T_26182_10_ctrl_is_load : _GEN_4971; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5050 = 5'ha == T_29096 ? T_26182_10_ctrl_is_sta : _GEN_4972; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5051 = 5'ha == T_29096 ? T_26182_10_ctrl_is_std : _GEN_4973; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5052 = 5'ha == T_29096 ? T_26182_10_wakeup_delay : _GEN_4974; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5053 = 5'ha == T_29096 ? T_26182_10_allocate_brtag : _GEN_4975; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5054 = 5'ha == T_29096 ? T_26182_10_is_br_or_jmp : _GEN_4976; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5055 = 5'ha == T_29096 ? T_26182_10_is_jump : _GEN_4977; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5056 = 5'ha == T_29096 ? T_26182_10_is_jal : _GEN_4978; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5057 = 5'ha == T_29096 ? T_26182_10_is_ret : _GEN_4979; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5058 = 5'ha == T_29096 ? T_26182_10_is_call : _GEN_4980; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5059 = 5'ha == T_29096 ? T_26182_10_br_mask : _GEN_4981; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5060 = 5'ha == T_29096 ? T_26182_10_br_tag : _GEN_4982; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5061 = 5'ha == T_29096 ? T_26182_10_br_prediction_bpd_predict_val : _GEN_4983; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5062 = 5'ha == T_29096 ? T_26182_10_br_prediction_bpd_predict_taken : _GEN_4984; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5063 = 5'ha == T_29096 ? T_26182_10_br_prediction_btb_hit : _GEN_4985; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5064 = 5'ha == T_29096 ? T_26182_10_br_prediction_btb_predicted : _GEN_4986; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5065 = 5'ha == T_29096 ? T_26182_10_br_prediction_is_br_or_jalr : _GEN_4987; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5066 = 5'ha == T_29096 ? T_26182_10_stat_brjmp_mispredicted : _GEN_4988; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5067 = 5'ha == T_29096 ? T_26182_10_stat_btb_made_pred : _GEN_4989; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5068 = 5'ha == T_29096 ? T_26182_10_stat_btb_mispredicted : _GEN_4990; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5069 = 5'ha == T_29096 ? T_26182_10_stat_bpd_made_pred : _GEN_4991; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5070 = 5'ha == T_29096 ? T_26182_10_stat_bpd_mispredicted : _GEN_4992; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5071 = 5'ha == T_29096 ? T_26182_10_fetch_pc_lob : _GEN_4993; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5072 = 5'ha == T_29096 ? T_26182_10_imm_packed : _GEN_4994; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5073 = 5'ha == T_29096 ? T_26182_10_csr_addr : _GEN_4995; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5074 = 5'ha == T_29096 ? T_26182_10_rob_idx : _GEN_4996; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5075 = 5'ha == T_29096 ? T_26182_10_ldq_idx : _GEN_4997; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5076 = 5'ha == T_29096 ? T_26182_10_stq_idx : _GEN_4998; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5077 = 5'ha == T_29096 ? T_26182_10_brob_idx : _GEN_4999; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5078 = 5'ha == T_29096 ? T_26182_10_pdst : _GEN_5000; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5079 = 5'ha == T_29096 ? T_26182_10_pop1 : _GEN_5001; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5080 = 5'ha == T_29096 ? T_26182_10_pop2 : _GEN_5002; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5081 = 5'ha == T_29096 ? T_26182_10_pop3 : _GEN_5003; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5082 = 5'ha == T_29096 ? T_26182_10_prs1_busy : _GEN_5004; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5083 = 5'ha == T_29096 ? T_26182_10_prs2_busy : _GEN_5005; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5084 = 5'ha == T_29096 ? T_26182_10_prs3_busy : _GEN_5006; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5085 = 5'ha == T_29096 ? T_26182_10_stale_pdst : _GEN_5007; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5086 = 5'ha == T_29096 ? T_26182_10_exception : _GEN_5008; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5087 = 5'ha == T_29096 ? T_26182_10_exc_cause : _GEN_5009; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5088 = 5'ha == T_29096 ? T_26182_10_bypassable : _GEN_5010; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5089 = 5'ha == T_29096 ? T_26182_10_mem_cmd : _GEN_5011; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5090 = 5'ha == T_29096 ? T_26182_10_mem_typ : _GEN_5012; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5091 = 5'ha == T_29096 ? T_26182_10_is_fence : _GEN_5013; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5092 = 5'ha == T_29096 ? T_26182_10_is_fencei : _GEN_5014; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5093 = 5'ha == T_29096 ? T_26182_10_is_store : _GEN_5015; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5094 = 5'ha == T_29096 ? T_26182_10_is_amo : _GEN_5016; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5095 = 5'ha == T_29096 ? T_26182_10_is_load : _GEN_5017; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5096 = 5'ha == T_29096 ? T_26182_10_is_unique : _GEN_5018; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5097 = 5'ha == T_29096 ? T_26182_10_flush_on_commit : _GEN_5019; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5098 = 5'ha == T_29096 ? T_26182_10_ldst : _GEN_5020; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5099 = 5'ha == T_29096 ? T_26182_10_lrs1 : _GEN_5021; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5100 = 5'ha == T_29096 ? T_26182_10_lrs2 : _GEN_5022; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5101 = 5'ha == T_29096 ? T_26182_10_lrs3 : _GEN_5023; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5102 = 5'ha == T_29096 ? T_26182_10_ldst_val : _GEN_5024; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5103 = 5'ha == T_29096 ? T_26182_10_dst_rtype : _GEN_5025; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5104 = 5'ha == T_29096 ? T_26182_10_lrs1_rtype : _GEN_5026; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5105 = 5'ha == T_29096 ? T_26182_10_lrs2_rtype : _GEN_5027; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5106 = 5'ha == T_29096 ? T_26182_10_frs3_en : _GEN_5028; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5107 = 5'ha == T_29096 ? T_26182_10_fp_val : _GEN_5029; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5108 = 5'ha == T_29096 ? T_26182_10_fp_single : _GEN_5030; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5109 = 5'ha == T_29096 ? T_26182_10_xcpt_if : _GEN_5031; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5110 = 5'ha == T_29096 ? T_26182_10_replay_if : _GEN_5032; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5112 = 5'ha == T_29096 ? T_26182_10_debug_events_fetch_seq : _GEN_5034; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5113 = 5'hb == T_29096 ? T_26182_11_valid : _GEN_5035; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5114 = 5'hb == T_29096 ? T_26182_11_iw_state : _GEN_5036; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5115 = 5'hb == T_29096 ? T_26182_11_uopc : _GEN_5037; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5116 = 5'hb == T_29096 ? T_26182_11_inst : _GEN_5038; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5117 = 5'hb == T_29096 ? T_26182_11_pc : _GEN_5039; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5118 = 5'hb == T_29096 ? T_26182_11_fu_code : _GEN_5040; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5119 = 5'hb == T_29096 ? T_26182_11_ctrl_br_type : _GEN_5041; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5120 = 5'hb == T_29096 ? T_26182_11_ctrl_op1_sel : _GEN_5042; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5121 = 5'hb == T_29096 ? T_26182_11_ctrl_op2_sel : _GEN_5043; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5122 = 5'hb == T_29096 ? T_26182_11_ctrl_imm_sel : _GEN_5044; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5123 = 5'hb == T_29096 ? T_26182_11_ctrl_op_fcn : _GEN_5045; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5124 = 5'hb == T_29096 ? T_26182_11_ctrl_fcn_dw : _GEN_5046; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5125 = 5'hb == T_29096 ? T_26182_11_ctrl_rf_wen : _GEN_5047; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5126 = 5'hb == T_29096 ? T_26182_11_ctrl_csr_cmd : _GEN_5048; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5127 = 5'hb == T_29096 ? T_26182_11_ctrl_is_load : _GEN_5049; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5128 = 5'hb == T_29096 ? T_26182_11_ctrl_is_sta : _GEN_5050; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5129 = 5'hb == T_29096 ? T_26182_11_ctrl_is_std : _GEN_5051; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5130 = 5'hb == T_29096 ? T_26182_11_wakeup_delay : _GEN_5052; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5131 = 5'hb == T_29096 ? T_26182_11_allocate_brtag : _GEN_5053; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5132 = 5'hb == T_29096 ? T_26182_11_is_br_or_jmp : _GEN_5054; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5133 = 5'hb == T_29096 ? T_26182_11_is_jump : _GEN_5055; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5134 = 5'hb == T_29096 ? T_26182_11_is_jal : _GEN_5056; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5135 = 5'hb == T_29096 ? T_26182_11_is_ret : _GEN_5057; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5136 = 5'hb == T_29096 ? T_26182_11_is_call : _GEN_5058; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5137 = 5'hb == T_29096 ? T_26182_11_br_mask : _GEN_5059; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5138 = 5'hb == T_29096 ? T_26182_11_br_tag : _GEN_5060; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5139 = 5'hb == T_29096 ? T_26182_11_br_prediction_bpd_predict_val : _GEN_5061; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5140 = 5'hb == T_29096 ? T_26182_11_br_prediction_bpd_predict_taken : _GEN_5062; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5141 = 5'hb == T_29096 ? T_26182_11_br_prediction_btb_hit : _GEN_5063; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5142 = 5'hb == T_29096 ? T_26182_11_br_prediction_btb_predicted : _GEN_5064; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5143 = 5'hb == T_29096 ? T_26182_11_br_prediction_is_br_or_jalr : _GEN_5065; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5144 = 5'hb == T_29096 ? T_26182_11_stat_brjmp_mispredicted : _GEN_5066; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5145 = 5'hb == T_29096 ? T_26182_11_stat_btb_made_pred : _GEN_5067; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5146 = 5'hb == T_29096 ? T_26182_11_stat_btb_mispredicted : _GEN_5068; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5147 = 5'hb == T_29096 ? T_26182_11_stat_bpd_made_pred : _GEN_5069; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5148 = 5'hb == T_29096 ? T_26182_11_stat_bpd_mispredicted : _GEN_5070; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5149 = 5'hb == T_29096 ? T_26182_11_fetch_pc_lob : _GEN_5071; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5150 = 5'hb == T_29096 ? T_26182_11_imm_packed : _GEN_5072; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5151 = 5'hb == T_29096 ? T_26182_11_csr_addr : _GEN_5073; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5152 = 5'hb == T_29096 ? T_26182_11_rob_idx : _GEN_5074; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5153 = 5'hb == T_29096 ? T_26182_11_ldq_idx : _GEN_5075; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5154 = 5'hb == T_29096 ? T_26182_11_stq_idx : _GEN_5076; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5155 = 5'hb == T_29096 ? T_26182_11_brob_idx : _GEN_5077; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5156 = 5'hb == T_29096 ? T_26182_11_pdst : _GEN_5078; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5157 = 5'hb == T_29096 ? T_26182_11_pop1 : _GEN_5079; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5158 = 5'hb == T_29096 ? T_26182_11_pop2 : _GEN_5080; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5159 = 5'hb == T_29096 ? T_26182_11_pop3 : _GEN_5081; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5160 = 5'hb == T_29096 ? T_26182_11_prs1_busy : _GEN_5082; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5161 = 5'hb == T_29096 ? T_26182_11_prs2_busy : _GEN_5083; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5162 = 5'hb == T_29096 ? T_26182_11_prs3_busy : _GEN_5084; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5163 = 5'hb == T_29096 ? T_26182_11_stale_pdst : _GEN_5085; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5164 = 5'hb == T_29096 ? T_26182_11_exception : _GEN_5086; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5165 = 5'hb == T_29096 ? T_26182_11_exc_cause : _GEN_5087; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5166 = 5'hb == T_29096 ? T_26182_11_bypassable : _GEN_5088; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5167 = 5'hb == T_29096 ? T_26182_11_mem_cmd : _GEN_5089; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5168 = 5'hb == T_29096 ? T_26182_11_mem_typ : _GEN_5090; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5169 = 5'hb == T_29096 ? T_26182_11_is_fence : _GEN_5091; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5170 = 5'hb == T_29096 ? T_26182_11_is_fencei : _GEN_5092; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5171 = 5'hb == T_29096 ? T_26182_11_is_store : _GEN_5093; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5172 = 5'hb == T_29096 ? T_26182_11_is_amo : _GEN_5094; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5173 = 5'hb == T_29096 ? T_26182_11_is_load : _GEN_5095; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5174 = 5'hb == T_29096 ? T_26182_11_is_unique : _GEN_5096; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5175 = 5'hb == T_29096 ? T_26182_11_flush_on_commit : _GEN_5097; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5176 = 5'hb == T_29096 ? T_26182_11_ldst : _GEN_5098; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5177 = 5'hb == T_29096 ? T_26182_11_lrs1 : _GEN_5099; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5178 = 5'hb == T_29096 ? T_26182_11_lrs2 : _GEN_5100; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5179 = 5'hb == T_29096 ? T_26182_11_lrs3 : _GEN_5101; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5180 = 5'hb == T_29096 ? T_26182_11_ldst_val : _GEN_5102; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5181 = 5'hb == T_29096 ? T_26182_11_dst_rtype : _GEN_5103; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5182 = 5'hb == T_29096 ? T_26182_11_lrs1_rtype : _GEN_5104; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5183 = 5'hb == T_29096 ? T_26182_11_lrs2_rtype : _GEN_5105; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5184 = 5'hb == T_29096 ? T_26182_11_frs3_en : _GEN_5106; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5185 = 5'hb == T_29096 ? T_26182_11_fp_val : _GEN_5107; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5186 = 5'hb == T_29096 ? T_26182_11_fp_single : _GEN_5108; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5187 = 5'hb == T_29096 ? T_26182_11_xcpt_if : _GEN_5109; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5188 = 5'hb == T_29096 ? T_26182_11_replay_if : _GEN_5110; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5190 = 5'hb == T_29096 ? T_26182_11_debug_events_fetch_seq : _GEN_5112; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5191 = 5'hc == T_29096 ? T_26182_12_valid : _GEN_5113; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5192 = 5'hc == T_29096 ? T_26182_12_iw_state : _GEN_5114; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5193 = 5'hc == T_29096 ? T_26182_12_uopc : _GEN_5115; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5194 = 5'hc == T_29096 ? T_26182_12_inst : _GEN_5116; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5195 = 5'hc == T_29096 ? T_26182_12_pc : _GEN_5117; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5196 = 5'hc == T_29096 ? T_26182_12_fu_code : _GEN_5118; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5197 = 5'hc == T_29096 ? T_26182_12_ctrl_br_type : _GEN_5119; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5198 = 5'hc == T_29096 ? T_26182_12_ctrl_op1_sel : _GEN_5120; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5199 = 5'hc == T_29096 ? T_26182_12_ctrl_op2_sel : _GEN_5121; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5200 = 5'hc == T_29096 ? T_26182_12_ctrl_imm_sel : _GEN_5122; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5201 = 5'hc == T_29096 ? T_26182_12_ctrl_op_fcn : _GEN_5123; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5202 = 5'hc == T_29096 ? T_26182_12_ctrl_fcn_dw : _GEN_5124; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5203 = 5'hc == T_29096 ? T_26182_12_ctrl_rf_wen : _GEN_5125; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5204 = 5'hc == T_29096 ? T_26182_12_ctrl_csr_cmd : _GEN_5126; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5205 = 5'hc == T_29096 ? T_26182_12_ctrl_is_load : _GEN_5127; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5206 = 5'hc == T_29096 ? T_26182_12_ctrl_is_sta : _GEN_5128; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5207 = 5'hc == T_29096 ? T_26182_12_ctrl_is_std : _GEN_5129; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5208 = 5'hc == T_29096 ? T_26182_12_wakeup_delay : _GEN_5130; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5209 = 5'hc == T_29096 ? T_26182_12_allocate_brtag : _GEN_5131; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5210 = 5'hc == T_29096 ? T_26182_12_is_br_or_jmp : _GEN_5132; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5211 = 5'hc == T_29096 ? T_26182_12_is_jump : _GEN_5133; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5212 = 5'hc == T_29096 ? T_26182_12_is_jal : _GEN_5134; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5213 = 5'hc == T_29096 ? T_26182_12_is_ret : _GEN_5135; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5214 = 5'hc == T_29096 ? T_26182_12_is_call : _GEN_5136; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5215 = 5'hc == T_29096 ? T_26182_12_br_mask : _GEN_5137; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5216 = 5'hc == T_29096 ? T_26182_12_br_tag : _GEN_5138; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5217 = 5'hc == T_29096 ? T_26182_12_br_prediction_bpd_predict_val : _GEN_5139; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5218 = 5'hc == T_29096 ? T_26182_12_br_prediction_bpd_predict_taken : _GEN_5140; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5219 = 5'hc == T_29096 ? T_26182_12_br_prediction_btb_hit : _GEN_5141; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5220 = 5'hc == T_29096 ? T_26182_12_br_prediction_btb_predicted : _GEN_5142; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5221 = 5'hc == T_29096 ? T_26182_12_br_prediction_is_br_or_jalr : _GEN_5143; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5222 = 5'hc == T_29096 ? T_26182_12_stat_brjmp_mispredicted : _GEN_5144; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5223 = 5'hc == T_29096 ? T_26182_12_stat_btb_made_pred : _GEN_5145; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5224 = 5'hc == T_29096 ? T_26182_12_stat_btb_mispredicted : _GEN_5146; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5225 = 5'hc == T_29096 ? T_26182_12_stat_bpd_made_pred : _GEN_5147; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5226 = 5'hc == T_29096 ? T_26182_12_stat_bpd_mispredicted : _GEN_5148; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5227 = 5'hc == T_29096 ? T_26182_12_fetch_pc_lob : _GEN_5149; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5228 = 5'hc == T_29096 ? T_26182_12_imm_packed : _GEN_5150; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5229 = 5'hc == T_29096 ? T_26182_12_csr_addr : _GEN_5151; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5230 = 5'hc == T_29096 ? T_26182_12_rob_idx : _GEN_5152; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5231 = 5'hc == T_29096 ? T_26182_12_ldq_idx : _GEN_5153; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5232 = 5'hc == T_29096 ? T_26182_12_stq_idx : _GEN_5154; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5233 = 5'hc == T_29096 ? T_26182_12_brob_idx : _GEN_5155; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5234 = 5'hc == T_29096 ? T_26182_12_pdst : _GEN_5156; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5235 = 5'hc == T_29096 ? T_26182_12_pop1 : _GEN_5157; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5236 = 5'hc == T_29096 ? T_26182_12_pop2 : _GEN_5158; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5237 = 5'hc == T_29096 ? T_26182_12_pop3 : _GEN_5159; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5238 = 5'hc == T_29096 ? T_26182_12_prs1_busy : _GEN_5160; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5239 = 5'hc == T_29096 ? T_26182_12_prs2_busy : _GEN_5161; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5240 = 5'hc == T_29096 ? T_26182_12_prs3_busy : _GEN_5162; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5241 = 5'hc == T_29096 ? T_26182_12_stale_pdst : _GEN_5163; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5242 = 5'hc == T_29096 ? T_26182_12_exception : _GEN_5164; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5243 = 5'hc == T_29096 ? T_26182_12_exc_cause : _GEN_5165; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5244 = 5'hc == T_29096 ? T_26182_12_bypassable : _GEN_5166; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5245 = 5'hc == T_29096 ? T_26182_12_mem_cmd : _GEN_5167; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5246 = 5'hc == T_29096 ? T_26182_12_mem_typ : _GEN_5168; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5247 = 5'hc == T_29096 ? T_26182_12_is_fence : _GEN_5169; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5248 = 5'hc == T_29096 ? T_26182_12_is_fencei : _GEN_5170; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5249 = 5'hc == T_29096 ? T_26182_12_is_store : _GEN_5171; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5250 = 5'hc == T_29096 ? T_26182_12_is_amo : _GEN_5172; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5251 = 5'hc == T_29096 ? T_26182_12_is_load : _GEN_5173; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5252 = 5'hc == T_29096 ? T_26182_12_is_unique : _GEN_5174; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5253 = 5'hc == T_29096 ? T_26182_12_flush_on_commit : _GEN_5175; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5254 = 5'hc == T_29096 ? T_26182_12_ldst : _GEN_5176; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5255 = 5'hc == T_29096 ? T_26182_12_lrs1 : _GEN_5177; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5256 = 5'hc == T_29096 ? T_26182_12_lrs2 : _GEN_5178; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5257 = 5'hc == T_29096 ? T_26182_12_lrs3 : _GEN_5179; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5258 = 5'hc == T_29096 ? T_26182_12_ldst_val : _GEN_5180; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5259 = 5'hc == T_29096 ? T_26182_12_dst_rtype : _GEN_5181; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5260 = 5'hc == T_29096 ? T_26182_12_lrs1_rtype : _GEN_5182; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5261 = 5'hc == T_29096 ? T_26182_12_lrs2_rtype : _GEN_5183; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5262 = 5'hc == T_29096 ? T_26182_12_frs3_en : _GEN_5184; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5263 = 5'hc == T_29096 ? T_26182_12_fp_val : _GEN_5185; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5264 = 5'hc == T_29096 ? T_26182_12_fp_single : _GEN_5186; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5265 = 5'hc == T_29096 ? T_26182_12_xcpt_if : _GEN_5187; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5266 = 5'hc == T_29096 ? T_26182_12_replay_if : _GEN_5188; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5268 = 5'hc == T_29096 ? T_26182_12_debug_events_fetch_seq : _GEN_5190; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5269 = 5'hd == T_29096 ? T_26182_13_valid : _GEN_5191; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5270 = 5'hd == T_29096 ? T_26182_13_iw_state : _GEN_5192; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5271 = 5'hd == T_29096 ? T_26182_13_uopc : _GEN_5193; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5272 = 5'hd == T_29096 ? T_26182_13_inst : _GEN_5194; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5273 = 5'hd == T_29096 ? T_26182_13_pc : _GEN_5195; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5274 = 5'hd == T_29096 ? T_26182_13_fu_code : _GEN_5196; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5275 = 5'hd == T_29096 ? T_26182_13_ctrl_br_type : _GEN_5197; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5276 = 5'hd == T_29096 ? T_26182_13_ctrl_op1_sel : _GEN_5198; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5277 = 5'hd == T_29096 ? T_26182_13_ctrl_op2_sel : _GEN_5199; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5278 = 5'hd == T_29096 ? T_26182_13_ctrl_imm_sel : _GEN_5200; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5279 = 5'hd == T_29096 ? T_26182_13_ctrl_op_fcn : _GEN_5201; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5280 = 5'hd == T_29096 ? T_26182_13_ctrl_fcn_dw : _GEN_5202; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5281 = 5'hd == T_29096 ? T_26182_13_ctrl_rf_wen : _GEN_5203; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5282 = 5'hd == T_29096 ? T_26182_13_ctrl_csr_cmd : _GEN_5204; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5283 = 5'hd == T_29096 ? T_26182_13_ctrl_is_load : _GEN_5205; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5284 = 5'hd == T_29096 ? T_26182_13_ctrl_is_sta : _GEN_5206; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5285 = 5'hd == T_29096 ? T_26182_13_ctrl_is_std : _GEN_5207; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5286 = 5'hd == T_29096 ? T_26182_13_wakeup_delay : _GEN_5208; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5287 = 5'hd == T_29096 ? T_26182_13_allocate_brtag : _GEN_5209; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5288 = 5'hd == T_29096 ? T_26182_13_is_br_or_jmp : _GEN_5210; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5289 = 5'hd == T_29096 ? T_26182_13_is_jump : _GEN_5211; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5290 = 5'hd == T_29096 ? T_26182_13_is_jal : _GEN_5212; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5291 = 5'hd == T_29096 ? T_26182_13_is_ret : _GEN_5213; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5292 = 5'hd == T_29096 ? T_26182_13_is_call : _GEN_5214; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5293 = 5'hd == T_29096 ? T_26182_13_br_mask : _GEN_5215; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5294 = 5'hd == T_29096 ? T_26182_13_br_tag : _GEN_5216; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5295 = 5'hd == T_29096 ? T_26182_13_br_prediction_bpd_predict_val : _GEN_5217; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5296 = 5'hd == T_29096 ? T_26182_13_br_prediction_bpd_predict_taken : _GEN_5218; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5297 = 5'hd == T_29096 ? T_26182_13_br_prediction_btb_hit : _GEN_5219; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5298 = 5'hd == T_29096 ? T_26182_13_br_prediction_btb_predicted : _GEN_5220; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5299 = 5'hd == T_29096 ? T_26182_13_br_prediction_is_br_or_jalr : _GEN_5221; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5300 = 5'hd == T_29096 ? T_26182_13_stat_brjmp_mispredicted : _GEN_5222; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5301 = 5'hd == T_29096 ? T_26182_13_stat_btb_made_pred : _GEN_5223; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5302 = 5'hd == T_29096 ? T_26182_13_stat_btb_mispredicted : _GEN_5224; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5303 = 5'hd == T_29096 ? T_26182_13_stat_bpd_made_pred : _GEN_5225; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5304 = 5'hd == T_29096 ? T_26182_13_stat_bpd_mispredicted : _GEN_5226; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5305 = 5'hd == T_29096 ? T_26182_13_fetch_pc_lob : _GEN_5227; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5306 = 5'hd == T_29096 ? T_26182_13_imm_packed : _GEN_5228; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5307 = 5'hd == T_29096 ? T_26182_13_csr_addr : _GEN_5229; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5308 = 5'hd == T_29096 ? T_26182_13_rob_idx : _GEN_5230; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5309 = 5'hd == T_29096 ? T_26182_13_ldq_idx : _GEN_5231; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5310 = 5'hd == T_29096 ? T_26182_13_stq_idx : _GEN_5232; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5311 = 5'hd == T_29096 ? T_26182_13_brob_idx : _GEN_5233; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5312 = 5'hd == T_29096 ? T_26182_13_pdst : _GEN_5234; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5313 = 5'hd == T_29096 ? T_26182_13_pop1 : _GEN_5235; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5314 = 5'hd == T_29096 ? T_26182_13_pop2 : _GEN_5236; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5315 = 5'hd == T_29096 ? T_26182_13_pop3 : _GEN_5237; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5316 = 5'hd == T_29096 ? T_26182_13_prs1_busy : _GEN_5238; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5317 = 5'hd == T_29096 ? T_26182_13_prs2_busy : _GEN_5239; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5318 = 5'hd == T_29096 ? T_26182_13_prs3_busy : _GEN_5240; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5319 = 5'hd == T_29096 ? T_26182_13_stale_pdst : _GEN_5241; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5320 = 5'hd == T_29096 ? T_26182_13_exception : _GEN_5242; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5321 = 5'hd == T_29096 ? T_26182_13_exc_cause : _GEN_5243; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5322 = 5'hd == T_29096 ? T_26182_13_bypassable : _GEN_5244; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5323 = 5'hd == T_29096 ? T_26182_13_mem_cmd : _GEN_5245; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5324 = 5'hd == T_29096 ? T_26182_13_mem_typ : _GEN_5246; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5325 = 5'hd == T_29096 ? T_26182_13_is_fence : _GEN_5247; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5326 = 5'hd == T_29096 ? T_26182_13_is_fencei : _GEN_5248; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5327 = 5'hd == T_29096 ? T_26182_13_is_store : _GEN_5249; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5328 = 5'hd == T_29096 ? T_26182_13_is_amo : _GEN_5250; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5329 = 5'hd == T_29096 ? T_26182_13_is_load : _GEN_5251; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5330 = 5'hd == T_29096 ? T_26182_13_is_unique : _GEN_5252; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5331 = 5'hd == T_29096 ? T_26182_13_flush_on_commit : _GEN_5253; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5332 = 5'hd == T_29096 ? T_26182_13_ldst : _GEN_5254; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5333 = 5'hd == T_29096 ? T_26182_13_lrs1 : _GEN_5255; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5334 = 5'hd == T_29096 ? T_26182_13_lrs2 : _GEN_5256; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5335 = 5'hd == T_29096 ? T_26182_13_lrs3 : _GEN_5257; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5336 = 5'hd == T_29096 ? T_26182_13_ldst_val : _GEN_5258; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5337 = 5'hd == T_29096 ? T_26182_13_dst_rtype : _GEN_5259; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5338 = 5'hd == T_29096 ? T_26182_13_lrs1_rtype : _GEN_5260; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5339 = 5'hd == T_29096 ? T_26182_13_lrs2_rtype : _GEN_5261; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5340 = 5'hd == T_29096 ? T_26182_13_frs3_en : _GEN_5262; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5341 = 5'hd == T_29096 ? T_26182_13_fp_val : _GEN_5263; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5342 = 5'hd == T_29096 ? T_26182_13_fp_single : _GEN_5264; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5343 = 5'hd == T_29096 ? T_26182_13_xcpt_if : _GEN_5265; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5344 = 5'hd == T_29096 ? T_26182_13_replay_if : _GEN_5266; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5346 = 5'hd == T_29096 ? T_26182_13_debug_events_fetch_seq : _GEN_5268; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5347 = 5'he == T_29096 ? T_26182_14_valid : _GEN_5269; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5348 = 5'he == T_29096 ? T_26182_14_iw_state : _GEN_5270; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5349 = 5'he == T_29096 ? T_26182_14_uopc : _GEN_5271; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5350 = 5'he == T_29096 ? T_26182_14_inst : _GEN_5272; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5351 = 5'he == T_29096 ? T_26182_14_pc : _GEN_5273; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5352 = 5'he == T_29096 ? T_26182_14_fu_code : _GEN_5274; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5353 = 5'he == T_29096 ? T_26182_14_ctrl_br_type : _GEN_5275; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5354 = 5'he == T_29096 ? T_26182_14_ctrl_op1_sel : _GEN_5276; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5355 = 5'he == T_29096 ? T_26182_14_ctrl_op2_sel : _GEN_5277; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5356 = 5'he == T_29096 ? T_26182_14_ctrl_imm_sel : _GEN_5278; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5357 = 5'he == T_29096 ? T_26182_14_ctrl_op_fcn : _GEN_5279; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5358 = 5'he == T_29096 ? T_26182_14_ctrl_fcn_dw : _GEN_5280; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5359 = 5'he == T_29096 ? T_26182_14_ctrl_rf_wen : _GEN_5281; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5360 = 5'he == T_29096 ? T_26182_14_ctrl_csr_cmd : _GEN_5282; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5361 = 5'he == T_29096 ? T_26182_14_ctrl_is_load : _GEN_5283; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5362 = 5'he == T_29096 ? T_26182_14_ctrl_is_sta : _GEN_5284; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5363 = 5'he == T_29096 ? T_26182_14_ctrl_is_std : _GEN_5285; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5364 = 5'he == T_29096 ? T_26182_14_wakeup_delay : _GEN_5286; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5365 = 5'he == T_29096 ? T_26182_14_allocate_brtag : _GEN_5287; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5366 = 5'he == T_29096 ? T_26182_14_is_br_or_jmp : _GEN_5288; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5367 = 5'he == T_29096 ? T_26182_14_is_jump : _GEN_5289; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5368 = 5'he == T_29096 ? T_26182_14_is_jal : _GEN_5290; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5369 = 5'he == T_29096 ? T_26182_14_is_ret : _GEN_5291; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5370 = 5'he == T_29096 ? T_26182_14_is_call : _GEN_5292; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5371 = 5'he == T_29096 ? T_26182_14_br_mask : _GEN_5293; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5372 = 5'he == T_29096 ? T_26182_14_br_tag : _GEN_5294; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5373 = 5'he == T_29096 ? T_26182_14_br_prediction_bpd_predict_val : _GEN_5295; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5374 = 5'he == T_29096 ? T_26182_14_br_prediction_bpd_predict_taken : _GEN_5296; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5375 = 5'he == T_29096 ? T_26182_14_br_prediction_btb_hit : _GEN_5297; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5376 = 5'he == T_29096 ? T_26182_14_br_prediction_btb_predicted : _GEN_5298; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5377 = 5'he == T_29096 ? T_26182_14_br_prediction_is_br_or_jalr : _GEN_5299; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5378 = 5'he == T_29096 ? T_26182_14_stat_brjmp_mispredicted : _GEN_5300; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5379 = 5'he == T_29096 ? T_26182_14_stat_btb_made_pred : _GEN_5301; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5380 = 5'he == T_29096 ? T_26182_14_stat_btb_mispredicted : _GEN_5302; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5381 = 5'he == T_29096 ? T_26182_14_stat_bpd_made_pred : _GEN_5303; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5382 = 5'he == T_29096 ? T_26182_14_stat_bpd_mispredicted : _GEN_5304; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5383 = 5'he == T_29096 ? T_26182_14_fetch_pc_lob : _GEN_5305; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5384 = 5'he == T_29096 ? T_26182_14_imm_packed : _GEN_5306; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5385 = 5'he == T_29096 ? T_26182_14_csr_addr : _GEN_5307; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5386 = 5'he == T_29096 ? T_26182_14_rob_idx : _GEN_5308; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5387 = 5'he == T_29096 ? T_26182_14_ldq_idx : _GEN_5309; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5388 = 5'he == T_29096 ? T_26182_14_stq_idx : _GEN_5310; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5389 = 5'he == T_29096 ? T_26182_14_brob_idx : _GEN_5311; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5390 = 5'he == T_29096 ? T_26182_14_pdst : _GEN_5312; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5391 = 5'he == T_29096 ? T_26182_14_pop1 : _GEN_5313; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5392 = 5'he == T_29096 ? T_26182_14_pop2 : _GEN_5314; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5393 = 5'he == T_29096 ? T_26182_14_pop3 : _GEN_5315; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5394 = 5'he == T_29096 ? T_26182_14_prs1_busy : _GEN_5316; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5395 = 5'he == T_29096 ? T_26182_14_prs2_busy : _GEN_5317; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5396 = 5'he == T_29096 ? T_26182_14_prs3_busy : _GEN_5318; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5397 = 5'he == T_29096 ? T_26182_14_stale_pdst : _GEN_5319; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5398 = 5'he == T_29096 ? T_26182_14_exception : _GEN_5320; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5399 = 5'he == T_29096 ? T_26182_14_exc_cause : _GEN_5321; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5400 = 5'he == T_29096 ? T_26182_14_bypassable : _GEN_5322; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5401 = 5'he == T_29096 ? T_26182_14_mem_cmd : _GEN_5323; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5402 = 5'he == T_29096 ? T_26182_14_mem_typ : _GEN_5324; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5403 = 5'he == T_29096 ? T_26182_14_is_fence : _GEN_5325; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5404 = 5'he == T_29096 ? T_26182_14_is_fencei : _GEN_5326; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5405 = 5'he == T_29096 ? T_26182_14_is_store : _GEN_5327; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5406 = 5'he == T_29096 ? T_26182_14_is_amo : _GEN_5328; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5407 = 5'he == T_29096 ? T_26182_14_is_load : _GEN_5329; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5408 = 5'he == T_29096 ? T_26182_14_is_unique : _GEN_5330; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5409 = 5'he == T_29096 ? T_26182_14_flush_on_commit : _GEN_5331; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5410 = 5'he == T_29096 ? T_26182_14_ldst : _GEN_5332; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5411 = 5'he == T_29096 ? T_26182_14_lrs1 : _GEN_5333; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5412 = 5'he == T_29096 ? T_26182_14_lrs2 : _GEN_5334; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5413 = 5'he == T_29096 ? T_26182_14_lrs3 : _GEN_5335; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5414 = 5'he == T_29096 ? T_26182_14_ldst_val : _GEN_5336; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5415 = 5'he == T_29096 ? T_26182_14_dst_rtype : _GEN_5337; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5416 = 5'he == T_29096 ? T_26182_14_lrs1_rtype : _GEN_5338; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5417 = 5'he == T_29096 ? T_26182_14_lrs2_rtype : _GEN_5339; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5418 = 5'he == T_29096 ? T_26182_14_frs3_en : _GEN_5340; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5419 = 5'he == T_29096 ? T_26182_14_fp_val : _GEN_5341; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5420 = 5'he == T_29096 ? T_26182_14_fp_single : _GEN_5342; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5421 = 5'he == T_29096 ? T_26182_14_xcpt_if : _GEN_5343; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5422 = 5'he == T_29096 ? T_26182_14_replay_if : _GEN_5344; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5424 = 5'he == T_29096 ? T_26182_14_debug_events_fetch_seq : _GEN_5346; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5425 = 5'hf == T_29096 ? T_26182_15_valid : _GEN_5347; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5426 = 5'hf == T_29096 ? T_26182_15_iw_state : _GEN_5348; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5427 = 5'hf == T_29096 ? T_26182_15_uopc : _GEN_5349; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5428 = 5'hf == T_29096 ? T_26182_15_inst : _GEN_5350; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5429 = 5'hf == T_29096 ? T_26182_15_pc : _GEN_5351; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5430 = 5'hf == T_29096 ? T_26182_15_fu_code : _GEN_5352; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5431 = 5'hf == T_29096 ? T_26182_15_ctrl_br_type : _GEN_5353; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5432 = 5'hf == T_29096 ? T_26182_15_ctrl_op1_sel : _GEN_5354; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5433 = 5'hf == T_29096 ? T_26182_15_ctrl_op2_sel : _GEN_5355; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5434 = 5'hf == T_29096 ? T_26182_15_ctrl_imm_sel : _GEN_5356; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5435 = 5'hf == T_29096 ? T_26182_15_ctrl_op_fcn : _GEN_5357; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5436 = 5'hf == T_29096 ? T_26182_15_ctrl_fcn_dw : _GEN_5358; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5437 = 5'hf == T_29096 ? T_26182_15_ctrl_rf_wen : _GEN_5359; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5438 = 5'hf == T_29096 ? T_26182_15_ctrl_csr_cmd : _GEN_5360; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5439 = 5'hf == T_29096 ? T_26182_15_ctrl_is_load : _GEN_5361; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5440 = 5'hf == T_29096 ? T_26182_15_ctrl_is_sta : _GEN_5362; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5441 = 5'hf == T_29096 ? T_26182_15_ctrl_is_std : _GEN_5363; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5442 = 5'hf == T_29096 ? T_26182_15_wakeup_delay : _GEN_5364; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5443 = 5'hf == T_29096 ? T_26182_15_allocate_brtag : _GEN_5365; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5444 = 5'hf == T_29096 ? T_26182_15_is_br_or_jmp : _GEN_5366; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5445 = 5'hf == T_29096 ? T_26182_15_is_jump : _GEN_5367; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5446 = 5'hf == T_29096 ? T_26182_15_is_jal : _GEN_5368; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5447 = 5'hf == T_29096 ? T_26182_15_is_ret : _GEN_5369; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5448 = 5'hf == T_29096 ? T_26182_15_is_call : _GEN_5370; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5449 = 5'hf == T_29096 ? T_26182_15_br_mask : _GEN_5371; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5450 = 5'hf == T_29096 ? T_26182_15_br_tag : _GEN_5372; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5451 = 5'hf == T_29096 ? T_26182_15_br_prediction_bpd_predict_val : _GEN_5373; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5452 = 5'hf == T_29096 ? T_26182_15_br_prediction_bpd_predict_taken : _GEN_5374; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5453 = 5'hf == T_29096 ? T_26182_15_br_prediction_btb_hit : _GEN_5375; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5454 = 5'hf == T_29096 ? T_26182_15_br_prediction_btb_predicted : _GEN_5376; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5455 = 5'hf == T_29096 ? T_26182_15_br_prediction_is_br_or_jalr : _GEN_5377; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5456 = 5'hf == T_29096 ? T_26182_15_stat_brjmp_mispredicted : _GEN_5378; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5457 = 5'hf == T_29096 ? T_26182_15_stat_btb_made_pred : _GEN_5379; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5458 = 5'hf == T_29096 ? T_26182_15_stat_btb_mispredicted : _GEN_5380; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5459 = 5'hf == T_29096 ? T_26182_15_stat_bpd_made_pred : _GEN_5381; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5460 = 5'hf == T_29096 ? T_26182_15_stat_bpd_mispredicted : _GEN_5382; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5461 = 5'hf == T_29096 ? T_26182_15_fetch_pc_lob : _GEN_5383; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5462 = 5'hf == T_29096 ? T_26182_15_imm_packed : _GEN_5384; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5463 = 5'hf == T_29096 ? T_26182_15_csr_addr : _GEN_5385; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5464 = 5'hf == T_29096 ? T_26182_15_rob_idx : _GEN_5386; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5465 = 5'hf == T_29096 ? T_26182_15_ldq_idx : _GEN_5387; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5466 = 5'hf == T_29096 ? T_26182_15_stq_idx : _GEN_5388; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5467 = 5'hf == T_29096 ? T_26182_15_brob_idx : _GEN_5389; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5468 = 5'hf == T_29096 ? T_26182_15_pdst : _GEN_5390; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5469 = 5'hf == T_29096 ? T_26182_15_pop1 : _GEN_5391; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5470 = 5'hf == T_29096 ? T_26182_15_pop2 : _GEN_5392; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5471 = 5'hf == T_29096 ? T_26182_15_pop3 : _GEN_5393; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5472 = 5'hf == T_29096 ? T_26182_15_prs1_busy : _GEN_5394; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5473 = 5'hf == T_29096 ? T_26182_15_prs2_busy : _GEN_5395; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5474 = 5'hf == T_29096 ? T_26182_15_prs3_busy : _GEN_5396; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5475 = 5'hf == T_29096 ? T_26182_15_stale_pdst : _GEN_5397; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5476 = 5'hf == T_29096 ? T_26182_15_exception : _GEN_5398; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5477 = 5'hf == T_29096 ? T_26182_15_exc_cause : _GEN_5399; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5478 = 5'hf == T_29096 ? T_26182_15_bypassable : _GEN_5400; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5479 = 5'hf == T_29096 ? T_26182_15_mem_cmd : _GEN_5401; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5480 = 5'hf == T_29096 ? T_26182_15_mem_typ : _GEN_5402; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5481 = 5'hf == T_29096 ? T_26182_15_is_fence : _GEN_5403; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5482 = 5'hf == T_29096 ? T_26182_15_is_fencei : _GEN_5404; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5483 = 5'hf == T_29096 ? T_26182_15_is_store : _GEN_5405; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5484 = 5'hf == T_29096 ? T_26182_15_is_amo : _GEN_5406; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5485 = 5'hf == T_29096 ? T_26182_15_is_load : _GEN_5407; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5486 = 5'hf == T_29096 ? T_26182_15_is_unique : _GEN_5408; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5487 = 5'hf == T_29096 ? T_26182_15_flush_on_commit : _GEN_5409; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5488 = 5'hf == T_29096 ? T_26182_15_ldst : _GEN_5410; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5489 = 5'hf == T_29096 ? T_26182_15_lrs1 : _GEN_5411; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5490 = 5'hf == T_29096 ? T_26182_15_lrs2 : _GEN_5412; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5491 = 5'hf == T_29096 ? T_26182_15_lrs3 : _GEN_5413; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5492 = 5'hf == T_29096 ? T_26182_15_ldst_val : _GEN_5414; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5493 = 5'hf == T_29096 ? T_26182_15_dst_rtype : _GEN_5415; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5494 = 5'hf == T_29096 ? T_26182_15_lrs1_rtype : _GEN_5416; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5495 = 5'hf == T_29096 ? T_26182_15_lrs2_rtype : _GEN_5417; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5496 = 5'hf == T_29096 ? T_26182_15_frs3_en : _GEN_5418; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5497 = 5'hf == T_29096 ? T_26182_15_fp_val : _GEN_5419; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5498 = 5'hf == T_29096 ? T_26182_15_fp_single : _GEN_5420; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5499 = 5'hf == T_29096 ? T_26182_15_xcpt_if : _GEN_5421; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5500 = 5'hf == T_29096 ? T_26182_15_replay_if : _GEN_5422; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5502 = 5'hf == T_29096 ? T_26182_15_debug_events_fetch_seq : _GEN_5424; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5503 = 5'h10 == T_29096 ? T_26182_16_valid : _GEN_5425; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5504 = 5'h10 == T_29096 ? T_26182_16_iw_state : _GEN_5426; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5505 = 5'h10 == T_29096 ? T_26182_16_uopc : _GEN_5427; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5506 = 5'h10 == T_29096 ? T_26182_16_inst : _GEN_5428; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5507 = 5'h10 == T_29096 ? T_26182_16_pc : _GEN_5429; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5508 = 5'h10 == T_29096 ? T_26182_16_fu_code : _GEN_5430; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5509 = 5'h10 == T_29096 ? T_26182_16_ctrl_br_type : _GEN_5431; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5510 = 5'h10 == T_29096 ? T_26182_16_ctrl_op1_sel : _GEN_5432; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5511 = 5'h10 == T_29096 ? T_26182_16_ctrl_op2_sel : _GEN_5433; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5512 = 5'h10 == T_29096 ? T_26182_16_ctrl_imm_sel : _GEN_5434; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5513 = 5'h10 == T_29096 ? T_26182_16_ctrl_op_fcn : _GEN_5435; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5514 = 5'h10 == T_29096 ? T_26182_16_ctrl_fcn_dw : _GEN_5436; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5515 = 5'h10 == T_29096 ? T_26182_16_ctrl_rf_wen : _GEN_5437; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5516 = 5'h10 == T_29096 ? T_26182_16_ctrl_csr_cmd : _GEN_5438; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5517 = 5'h10 == T_29096 ? T_26182_16_ctrl_is_load : _GEN_5439; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5518 = 5'h10 == T_29096 ? T_26182_16_ctrl_is_sta : _GEN_5440; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5519 = 5'h10 == T_29096 ? T_26182_16_ctrl_is_std : _GEN_5441; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5520 = 5'h10 == T_29096 ? T_26182_16_wakeup_delay : _GEN_5442; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5521 = 5'h10 == T_29096 ? T_26182_16_allocate_brtag : _GEN_5443; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5522 = 5'h10 == T_29096 ? T_26182_16_is_br_or_jmp : _GEN_5444; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5523 = 5'h10 == T_29096 ? T_26182_16_is_jump : _GEN_5445; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5524 = 5'h10 == T_29096 ? T_26182_16_is_jal : _GEN_5446; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5525 = 5'h10 == T_29096 ? T_26182_16_is_ret : _GEN_5447; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5526 = 5'h10 == T_29096 ? T_26182_16_is_call : _GEN_5448; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5527 = 5'h10 == T_29096 ? T_26182_16_br_mask : _GEN_5449; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5528 = 5'h10 == T_29096 ? T_26182_16_br_tag : _GEN_5450; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5529 = 5'h10 == T_29096 ? T_26182_16_br_prediction_bpd_predict_val : _GEN_5451; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5530 = 5'h10 == T_29096 ? T_26182_16_br_prediction_bpd_predict_taken : _GEN_5452; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5531 = 5'h10 == T_29096 ? T_26182_16_br_prediction_btb_hit : _GEN_5453; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5532 = 5'h10 == T_29096 ? T_26182_16_br_prediction_btb_predicted : _GEN_5454; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5533 = 5'h10 == T_29096 ? T_26182_16_br_prediction_is_br_or_jalr : _GEN_5455; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5534 = 5'h10 == T_29096 ? T_26182_16_stat_brjmp_mispredicted : _GEN_5456; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5535 = 5'h10 == T_29096 ? T_26182_16_stat_btb_made_pred : _GEN_5457; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5536 = 5'h10 == T_29096 ? T_26182_16_stat_btb_mispredicted : _GEN_5458; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5537 = 5'h10 == T_29096 ? T_26182_16_stat_bpd_made_pred : _GEN_5459; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5538 = 5'h10 == T_29096 ? T_26182_16_stat_bpd_mispredicted : _GEN_5460; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5539 = 5'h10 == T_29096 ? T_26182_16_fetch_pc_lob : _GEN_5461; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5540 = 5'h10 == T_29096 ? T_26182_16_imm_packed : _GEN_5462; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5541 = 5'h10 == T_29096 ? T_26182_16_csr_addr : _GEN_5463; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5542 = 5'h10 == T_29096 ? T_26182_16_rob_idx : _GEN_5464; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5543 = 5'h10 == T_29096 ? T_26182_16_ldq_idx : _GEN_5465; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5544 = 5'h10 == T_29096 ? T_26182_16_stq_idx : _GEN_5466; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5545 = 5'h10 == T_29096 ? T_26182_16_brob_idx : _GEN_5467; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5546 = 5'h10 == T_29096 ? T_26182_16_pdst : _GEN_5468; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5547 = 5'h10 == T_29096 ? T_26182_16_pop1 : _GEN_5469; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5548 = 5'h10 == T_29096 ? T_26182_16_pop2 : _GEN_5470; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5549 = 5'h10 == T_29096 ? T_26182_16_pop3 : _GEN_5471; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5550 = 5'h10 == T_29096 ? T_26182_16_prs1_busy : _GEN_5472; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5551 = 5'h10 == T_29096 ? T_26182_16_prs2_busy : _GEN_5473; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5552 = 5'h10 == T_29096 ? T_26182_16_prs3_busy : _GEN_5474; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5553 = 5'h10 == T_29096 ? T_26182_16_stale_pdst : _GEN_5475; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5554 = 5'h10 == T_29096 ? T_26182_16_exception : _GEN_5476; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5555 = 5'h10 == T_29096 ? T_26182_16_exc_cause : _GEN_5477; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5556 = 5'h10 == T_29096 ? T_26182_16_bypassable : _GEN_5478; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5557 = 5'h10 == T_29096 ? T_26182_16_mem_cmd : _GEN_5479; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5558 = 5'h10 == T_29096 ? T_26182_16_mem_typ : _GEN_5480; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5559 = 5'h10 == T_29096 ? T_26182_16_is_fence : _GEN_5481; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5560 = 5'h10 == T_29096 ? T_26182_16_is_fencei : _GEN_5482; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5561 = 5'h10 == T_29096 ? T_26182_16_is_store : _GEN_5483; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5562 = 5'h10 == T_29096 ? T_26182_16_is_amo : _GEN_5484; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5563 = 5'h10 == T_29096 ? T_26182_16_is_load : _GEN_5485; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5564 = 5'h10 == T_29096 ? T_26182_16_is_unique : _GEN_5486; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5565 = 5'h10 == T_29096 ? T_26182_16_flush_on_commit : _GEN_5487; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5566 = 5'h10 == T_29096 ? T_26182_16_ldst : _GEN_5488; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5567 = 5'h10 == T_29096 ? T_26182_16_lrs1 : _GEN_5489; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5568 = 5'h10 == T_29096 ? T_26182_16_lrs2 : _GEN_5490; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5569 = 5'h10 == T_29096 ? T_26182_16_lrs3 : _GEN_5491; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5570 = 5'h10 == T_29096 ? T_26182_16_ldst_val : _GEN_5492; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5571 = 5'h10 == T_29096 ? T_26182_16_dst_rtype : _GEN_5493; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5572 = 5'h10 == T_29096 ? T_26182_16_lrs1_rtype : _GEN_5494; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5573 = 5'h10 == T_29096 ? T_26182_16_lrs2_rtype : _GEN_5495; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5574 = 5'h10 == T_29096 ? T_26182_16_frs3_en : _GEN_5496; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5575 = 5'h10 == T_29096 ? T_26182_16_fp_val : _GEN_5497; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5576 = 5'h10 == T_29096 ? T_26182_16_fp_single : _GEN_5498; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5577 = 5'h10 == T_29096 ? T_26182_16_xcpt_if : _GEN_5499; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5578 = 5'h10 == T_29096 ? T_26182_16_replay_if : _GEN_5500; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5580 = 5'h10 == T_29096 ? T_26182_16_debug_events_fetch_seq : _GEN_5502; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5581 = 5'h11 == T_29096 ? T_26182_17_valid : _GEN_5503; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5582 = 5'h11 == T_29096 ? T_26182_17_iw_state : _GEN_5504; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5583 = 5'h11 == T_29096 ? T_26182_17_uopc : _GEN_5505; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5584 = 5'h11 == T_29096 ? T_26182_17_inst : _GEN_5506; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5585 = 5'h11 == T_29096 ? T_26182_17_pc : _GEN_5507; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5586 = 5'h11 == T_29096 ? T_26182_17_fu_code : _GEN_5508; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5587 = 5'h11 == T_29096 ? T_26182_17_ctrl_br_type : _GEN_5509; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5588 = 5'h11 == T_29096 ? T_26182_17_ctrl_op1_sel : _GEN_5510; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5589 = 5'h11 == T_29096 ? T_26182_17_ctrl_op2_sel : _GEN_5511; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5590 = 5'h11 == T_29096 ? T_26182_17_ctrl_imm_sel : _GEN_5512; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5591 = 5'h11 == T_29096 ? T_26182_17_ctrl_op_fcn : _GEN_5513; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5592 = 5'h11 == T_29096 ? T_26182_17_ctrl_fcn_dw : _GEN_5514; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5593 = 5'h11 == T_29096 ? T_26182_17_ctrl_rf_wen : _GEN_5515; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5594 = 5'h11 == T_29096 ? T_26182_17_ctrl_csr_cmd : _GEN_5516; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5595 = 5'h11 == T_29096 ? T_26182_17_ctrl_is_load : _GEN_5517; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5596 = 5'h11 == T_29096 ? T_26182_17_ctrl_is_sta : _GEN_5518; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5597 = 5'h11 == T_29096 ? T_26182_17_ctrl_is_std : _GEN_5519; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5598 = 5'h11 == T_29096 ? T_26182_17_wakeup_delay : _GEN_5520; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5599 = 5'h11 == T_29096 ? T_26182_17_allocate_brtag : _GEN_5521; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5600 = 5'h11 == T_29096 ? T_26182_17_is_br_or_jmp : _GEN_5522; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5601 = 5'h11 == T_29096 ? T_26182_17_is_jump : _GEN_5523; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5602 = 5'h11 == T_29096 ? T_26182_17_is_jal : _GEN_5524; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5603 = 5'h11 == T_29096 ? T_26182_17_is_ret : _GEN_5525; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5604 = 5'h11 == T_29096 ? T_26182_17_is_call : _GEN_5526; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5605 = 5'h11 == T_29096 ? T_26182_17_br_mask : _GEN_5527; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5606 = 5'h11 == T_29096 ? T_26182_17_br_tag : _GEN_5528; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5607 = 5'h11 == T_29096 ? T_26182_17_br_prediction_bpd_predict_val : _GEN_5529; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5608 = 5'h11 == T_29096 ? T_26182_17_br_prediction_bpd_predict_taken : _GEN_5530; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5609 = 5'h11 == T_29096 ? T_26182_17_br_prediction_btb_hit : _GEN_5531; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5610 = 5'h11 == T_29096 ? T_26182_17_br_prediction_btb_predicted : _GEN_5532; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5611 = 5'h11 == T_29096 ? T_26182_17_br_prediction_is_br_or_jalr : _GEN_5533; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5612 = 5'h11 == T_29096 ? T_26182_17_stat_brjmp_mispredicted : _GEN_5534; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5613 = 5'h11 == T_29096 ? T_26182_17_stat_btb_made_pred : _GEN_5535; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5614 = 5'h11 == T_29096 ? T_26182_17_stat_btb_mispredicted : _GEN_5536; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5615 = 5'h11 == T_29096 ? T_26182_17_stat_bpd_made_pred : _GEN_5537; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5616 = 5'h11 == T_29096 ? T_26182_17_stat_bpd_mispredicted : _GEN_5538; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5617 = 5'h11 == T_29096 ? T_26182_17_fetch_pc_lob : _GEN_5539; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5618 = 5'h11 == T_29096 ? T_26182_17_imm_packed : _GEN_5540; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5619 = 5'h11 == T_29096 ? T_26182_17_csr_addr : _GEN_5541; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5620 = 5'h11 == T_29096 ? T_26182_17_rob_idx : _GEN_5542; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5621 = 5'h11 == T_29096 ? T_26182_17_ldq_idx : _GEN_5543; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5622 = 5'h11 == T_29096 ? T_26182_17_stq_idx : _GEN_5544; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5623 = 5'h11 == T_29096 ? T_26182_17_brob_idx : _GEN_5545; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5624 = 5'h11 == T_29096 ? T_26182_17_pdst : _GEN_5546; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5625 = 5'h11 == T_29096 ? T_26182_17_pop1 : _GEN_5547; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5626 = 5'h11 == T_29096 ? T_26182_17_pop2 : _GEN_5548; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5627 = 5'h11 == T_29096 ? T_26182_17_pop3 : _GEN_5549; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5628 = 5'h11 == T_29096 ? T_26182_17_prs1_busy : _GEN_5550; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5629 = 5'h11 == T_29096 ? T_26182_17_prs2_busy : _GEN_5551; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5630 = 5'h11 == T_29096 ? T_26182_17_prs3_busy : _GEN_5552; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5631 = 5'h11 == T_29096 ? T_26182_17_stale_pdst : _GEN_5553; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5632 = 5'h11 == T_29096 ? T_26182_17_exception : _GEN_5554; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5633 = 5'h11 == T_29096 ? T_26182_17_exc_cause : _GEN_5555; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5634 = 5'h11 == T_29096 ? T_26182_17_bypassable : _GEN_5556; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5635 = 5'h11 == T_29096 ? T_26182_17_mem_cmd : _GEN_5557; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5636 = 5'h11 == T_29096 ? T_26182_17_mem_typ : _GEN_5558; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5637 = 5'h11 == T_29096 ? T_26182_17_is_fence : _GEN_5559; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5638 = 5'h11 == T_29096 ? T_26182_17_is_fencei : _GEN_5560; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5639 = 5'h11 == T_29096 ? T_26182_17_is_store : _GEN_5561; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5640 = 5'h11 == T_29096 ? T_26182_17_is_amo : _GEN_5562; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5641 = 5'h11 == T_29096 ? T_26182_17_is_load : _GEN_5563; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5642 = 5'h11 == T_29096 ? T_26182_17_is_unique : _GEN_5564; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5643 = 5'h11 == T_29096 ? T_26182_17_flush_on_commit : _GEN_5565; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5644 = 5'h11 == T_29096 ? T_26182_17_ldst : _GEN_5566; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5645 = 5'h11 == T_29096 ? T_26182_17_lrs1 : _GEN_5567; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5646 = 5'h11 == T_29096 ? T_26182_17_lrs2 : _GEN_5568; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5647 = 5'h11 == T_29096 ? T_26182_17_lrs3 : _GEN_5569; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5648 = 5'h11 == T_29096 ? T_26182_17_ldst_val : _GEN_5570; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5649 = 5'h11 == T_29096 ? T_26182_17_dst_rtype : _GEN_5571; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5650 = 5'h11 == T_29096 ? T_26182_17_lrs1_rtype : _GEN_5572; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5651 = 5'h11 == T_29096 ? T_26182_17_lrs2_rtype : _GEN_5573; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5652 = 5'h11 == T_29096 ? T_26182_17_frs3_en : _GEN_5574; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5653 = 5'h11 == T_29096 ? T_26182_17_fp_val : _GEN_5575; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5654 = 5'h11 == T_29096 ? T_26182_17_fp_single : _GEN_5576; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5655 = 5'h11 == T_29096 ? T_26182_17_xcpt_if : _GEN_5577; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5656 = 5'h11 == T_29096 ? T_26182_17_replay_if : _GEN_5578; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5658 = 5'h11 == T_29096 ? T_26182_17_debug_events_fetch_seq : _GEN_5580; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5659 = 5'h12 == T_29096 ? T_26182_18_valid : _GEN_5581; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5660 = 5'h12 == T_29096 ? T_26182_18_iw_state : _GEN_5582; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5661 = 5'h12 == T_29096 ? T_26182_18_uopc : _GEN_5583; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5662 = 5'h12 == T_29096 ? T_26182_18_inst : _GEN_5584; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5663 = 5'h12 == T_29096 ? T_26182_18_pc : _GEN_5585; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5664 = 5'h12 == T_29096 ? T_26182_18_fu_code : _GEN_5586; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5665 = 5'h12 == T_29096 ? T_26182_18_ctrl_br_type : _GEN_5587; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5666 = 5'h12 == T_29096 ? T_26182_18_ctrl_op1_sel : _GEN_5588; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5667 = 5'h12 == T_29096 ? T_26182_18_ctrl_op2_sel : _GEN_5589; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5668 = 5'h12 == T_29096 ? T_26182_18_ctrl_imm_sel : _GEN_5590; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5669 = 5'h12 == T_29096 ? T_26182_18_ctrl_op_fcn : _GEN_5591; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5670 = 5'h12 == T_29096 ? T_26182_18_ctrl_fcn_dw : _GEN_5592; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5671 = 5'h12 == T_29096 ? T_26182_18_ctrl_rf_wen : _GEN_5593; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5672 = 5'h12 == T_29096 ? T_26182_18_ctrl_csr_cmd : _GEN_5594; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5673 = 5'h12 == T_29096 ? T_26182_18_ctrl_is_load : _GEN_5595; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5674 = 5'h12 == T_29096 ? T_26182_18_ctrl_is_sta : _GEN_5596; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5675 = 5'h12 == T_29096 ? T_26182_18_ctrl_is_std : _GEN_5597; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5676 = 5'h12 == T_29096 ? T_26182_18_wakeup_delay : _GEN_5598; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5677 = 5'h12 == T_29096 ? T_26182_18_allocate_brtag : _GEN_5599; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5678 = 5'h12 == T_29096 ? T_26182_18_is_br_or_jmp : _GEN_5600; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5679 = 5'h12 == T_29096 ? T_26182_18_is_jump : _GEN_5601; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5680 = 5'h12 == T_29096 ? T_26182_18_is_jal : _GEN_5602; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5681 = 5'h12 == T_29096 ? T_26182_18_is_ret : _GEN_5603; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5682 = 5'h12 == T_29096 ? T_26182_18_is_call : _GEN_5604; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5683 = 5'h12 == T_29096 ? T_26182_18_br_mask : _GEN_5605; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5684 = 5'h12 == T_29096 ? T_26182_18_br_tag : _GEN_5606; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5685 = 5'h12 == T_29096 ? T_26182_18_br_prediction_bpd_predict_val : _GEN_5607; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5686 = 5'h12 == T_29096 ? T_26182_18_br_prediction_bpd_predict_taken : _GEN_5608; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5687 = 5'h12 == T_29096 ? T_26182_18_br_prediction_btb_hit : _GEN_5609; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5688 = 5'h12 == T_29096 ? T_26182_18_br_prediction_btb_predicted : _GEN_5610; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5689 = 5'h12 == T_29096 ? T_26182_18_br_prediction_is_br_or_jalr : _GEN_5611; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5690 = 5'h12 == T_29096 ? T_26182_18_stat_brjmp_mispredicted : _GEN_5612; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5691 = 5'h12 == T_29096 ? T_26182_18_stat_btb_made_pred : _GEN_5613; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5692 = 5'h12 == T_29096 ? T_26182_18_stat_btb_mispredicted : _GEN_5614; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5693 = 5'h12 == T_29096 ? T_26182_18_stat_bpd_made_pred : _GEN_5615; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5694 = 5'h12 == T_29096 ? T_26182_18_stat_bpd_mispredicted : _GEN_5616; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5695 = 5'h12 == T_29096 ? T_26182_18_fetch_pc_lob : _GEN_5617; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5696 = 5'h12 == T_29096 ? T_26182_18_imm_packed : _GEN_5618; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5697 = 5'h12 == T_29096 ? T_26182_18_csr_addr : _GEN_5619; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5698 = 5'h12 == T_29096 ? T_26182_18_rob_idx : _GEN_5620; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5699 = 5'h12 == T_29096 ? T_26182_18_ldq_idx : _GEN_5621; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5700 = 5'h12 == T_29096 ? T_26182_18_stq_idx : _GEN_5622; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5701 = 5'h12 == T_29096 ? T_26182_18_brob_idx : _GEN_5623; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5702 = 5'h12 == T_29096 ? T_26182_18_pdst : _GEN_5624; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5703 = 5'h12 == T_29096 ? T_26182_18_pop1 : _GEN_5625; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5704 = 5'h12 == T_29096 ? T_26182_18_pop2 : _GEN_5626; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5705 = 5'h12 == T_29096 ? T_26182_18_pop3 : _GEN_5627; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5706 = 5'h12 == T_29096 ? T_26182_18_prs1_busy : _GEN_5628; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5707 = 5'h12 == T_29096 ? T_26182_18_prs2_busy : _GEN_5629; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5708 = 5'h12 == T_29096 ? T_26182_18_prs3_busy : _GEN_5630; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5709 = 5'h12 == T_29096 ? T_26182_18_stale_pdst : _GEN_5631; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5710 = 5'h12 == T_29096 ? T_26182_18_exception : _GEN_5632; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5711 = 5'h12 == T_29096 ? T_26182_18_exc_cause : _GEN_5633; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5712 = 5'h12 == T_29096 ? T_26182_18_bypassable : _GEN_5634; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5713 = 5'h12 == T_29096 ? T_26182_18_mem_cmd : _GEN_5635; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5714 = 5'h12 == T_29096 ? T_26182_18_mem_typ : _GEN_5636; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5715 = 5'h12 == T_29096 ? T_26182_18_is_fence : _GEN_5637; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5716 = 5'h12 == T_29096 ? T_26182_18_is_fencei : _GEN_5638; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5717 = 5'h12 == T_29096 ? T_26182_18_is_store : _GEN_5639; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5718 = 5'h12 == T_29096 ? T_26182_18_is_amo : _GEN_5640; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5719 = 5'h12 == T_29096 ? T_26182_18_is_load : _GEN_5641; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5720 = 5'h12 == T_29096 ? T_26182_18_is_unique : _GEN_5642; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5721 = 5'h12 == T_29096 ? T_26182_18_flush_on_commit : _GEN_5643; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5722 = 5'h12 == T_29096 ? T_26182_18_ldst : _GEN_5644; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5723 = 5'h12 == T_29096 ? T_26182_18_lrs1 : _GEN_5645; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5724 = 5'h12 == T_29096 ? T_26182_18_lrs2 : _GEN_5646; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5725 = 5'h12 == T_29096 ? T_26182_18_lrs3 : _GEN_5647; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5726 = 5'h12 == T_29096 ? T_26182_18_ldst_val : _GEN_5648; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5727 = 5'h12 == T_29096 ? T_26182_18_dst_rtype : _GEN_5649; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5728 = 5'h12 == T_29096 ? T_26182_18_lrs1_rtype : _GEN_5650; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5729 = 5'h12 == T_29096 ? T_26182_18_lrs2_rtype : _GEN_5651; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5730 = 5'h12 == T_29096 ? T_26182_18_frs3_en : _GEN_5652; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5731 = 5'h12 == T_29096 ? T_26182_18_fp_val : _GEN_5653; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5732 = 5'h12 == T_29096 ? T_26182_18_fp_single : _GEN_5654; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5733 = 5'h12 == T_29096 ? T_26182_18_xcpt_if : _GEN_5655; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5734 = 5'h12 == T_29096 ? T_26182_18_replay_if : _GEN_5656; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5736 = 5'h12 == T_29096 ? T_26182_18_debug_events_fetch_seq : _GEN_5658; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5737 = 5'h13 == T_29096 ? T_26182_19_valid : _GEN_5659; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5738 = 5'h13 == T_29096 ? T_26182_19_iw_state : _GEN_5660; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5739 = 5'h13 == T_29096 ? T_26182_19_uopc : _GEN_5661; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5740 = 5'h13 == T_29096 ? T_26182_19_inst : _GEN_5662; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5741 = 5'h13 == T_29096 ? T_26182_19_pc : _GEN_5663; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5742 = 5'h13 == T_29096 ? T_26182_19_fu_code : _GEN_5664; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5743 = 5'h13 == T_29096 ? T_26182_19_ctrl_br_type : _GEN_5665; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5744 = 5'h13 == T_29096 ? T_26182_19_ctrl_op1_sel : _GEN_5666; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5745 = 5'h13 == T_29096 ? T_26182_19_ctrl_op2_sel : _GEN_5667; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5746 = 5'h13 == T_29096 ? T_26182_19_ctrl_imm_sel : _GEN_5668; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5747 = 5'h13 == T_29096 ? T_26182_19_ctrl_op_fcn : _GEN_5669; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5748 = 5'h13 == T_29096 ? T_26182_19_ctrl_fcn_dw : _GEN_5670; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5749 = 5'h13 == T_29096 ? T_26182_19_ctrl_rf_wen : _GEN_5671; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5750 = 5'h13 == T_29096 ? T_26182_19_ctrl_csr_cmd : _GEN_5672; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5751 = 5'h13 == T_29096 ? T_26182_19_ctrl_is_load : _GEN_5673; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5752 = 5'h13 == T_29096 ? T_26182_19_ctrl_is_sta : _GEN_5674; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5753 = 5'h13 == T_29096 ? T_26182_19_ctrl_is_std : _GEN_5675; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5754 = 5'h13 == T_29096 ? T_26182_19_wakeup_delay : _GEN_5676; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5755 = 5'h13 == T_29096 ? T_26182_19_allocate_brtag : _GEN_5677; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5756 = 5'h13 == T_29096 ? T_26182_19_is_br_or_jmp : _GEN_5678; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5757 = 5'h13 == T_29096 ? T_26182_19_is_jump : _GEN_5679; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5758 = 5'h13 == T_29096 ? T_26182_19_is_jal : _GEN_5680; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5759 = 5'h13 == T_29096 ? T_26182_19_is_ret : _GEN_5681; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5760 = 5'h13 == T_29096 ? T_26182_19_is_call : _GEN_5682; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5761 = 5'h13 == T_29096 ? T_26182_19_br_mask : _GEN_5683; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5762 = 5'h13 == T_29096 ? T_26182_19_br_tag : _GEN_5684; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5763 = 5'h13 == T_29096 ? T_26182_19_br_prediction_bpd_predict_val : _GEN_5685; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5764 = 5'h13 == T_29096 ? T_26182_19_br_prediction_bpd_predict_taken : _GEN_5686; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5765 = 5'h13 == T_29096 ? T_26182_19_br_prediction_btb_hit : _GEN_5687; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5766 = 5'h13 == T_29096 ? T_26182_19_br_prediction_btb_predicted : _GEN_5688; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5767 = 5'h13 == T_29096 ? T_26182_19_br_prediction_is_br_or_jalr : _GEN_5689; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5768 = 5'h13 == T_29096 ? T_26182_19_stat_brjmp_mispredicted : _GEN_5690; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5769 = 5'h13 == T_29096 ? T_26182_19_stat_btb_made_pred : _GEN_5691; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5770 = 5'h13 == T_29096 ? T_26182_19_stat_btb_mispredicted : _GEN_5692; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5771 = 5'h13 == T_29096 ? T_26182_19_stat_bpd_made_pred : _GEN_5693; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5772 = 5'h13 == T_29096 ? T_26182_19_stat_bpd_mispredicted : _GEN_5694; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5773 = 5'h13 == T_29096 ? T_26182_19_fetch_pc_lob : _GEN_5695; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5774 = 5'h13 == T_29096 ? T_26182_19_imm_packed : _GEN_5696; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5775 = 5'h13 == T_29096 ? T_26182_19_csr_addr : _GEN_5697; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5776 = 5'h13 == T_29096 ? T_26182_19_rob_idx : _GEN_5698; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5777 = 5'h13 == T_29096 ? T_26182_19_ldq_idx : _GEN_5699; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5778 = 5'h13 == T_29096 ? T_26182_19_stq_idx : _GEN_5700; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5779 = 5'h13 == T_29096 ? T_26182_19_brob_idx : _GEN_5701; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5780 = 5'h13 == T_29096 ? T_26182_19_pdst : _GEN_5702; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5781 = 5'h13 == T_29096 ? T_26182_19_pop1 : _GEN_5703; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5782 = 5'h13 == T_29096 ? T_26182_19_pop2 : _GEN_5704; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5783 = 5'h13 == T_29096 ? T_26182_19_pop3 : _GEN_5705; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5784 = 5'h13 == T_29096 ? T_26182_19_prs1_busy : _GEN_5706; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5785 = 5'h13 == T_29096 ? T_26182_19_prs2_busy : _GEN_5707; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5786 = 5'h13 == T_29096 ? T_26182_19_prs3_busy : _GEN_5708; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5787 = 5'h13 == T_29096 ? T_26182_19_stale_pdst : _GEN_5709; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5788 = 5'h13 == T_29096 ? T_26182_19_exception : _GEN_5710; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5789 = 5'h13 == T_29096 ? T_26182_19_exc_cause : _GEN_5711; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5790 = 5'h13 == T_29096 ? T_26182_19_bypassable : _GEN_5712; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5791 = 5'h13 == T_29096 ? T_26182_19_mem_cmd : _GEN_5713; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5792 = 5'h13 == T_29096 ? T_26182_19_mem_typ : _GEN_5714; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5793 = 5'h13 == T_29096 ? T_26182_19_is_fence : _GEN_5715; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5794 = 5'h13 == T_29096 ? T_26182_19_is_fencei : _GEN_5716; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5795 = 5'h13 == T_29096 ? T_26182_19_is_store : _GEN_5717; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5796 = 5'h13 == T_29096 ? T_26182_19_is_amo : _GEN_5718; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5797 = 5'h13 == T_29096 ? T_26182_19_is_load : _GEN_5719; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5798 = 5'h13 == T_29096 ? T_26182_19_is_unique : _GEN_5720; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5799 = 5'h13 == T_29096 ? T_26182_19_flush_on_commit : _GEN_5721; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5800 = 5'h13 == T_29096 ? T_26182_19_ldst : _GEN_5722; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5801 = 5'h13 == T_29096 ? T_26182_19_lrs1 : _GEN_5723; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5802 = 5'h13 == T_29096 ? T_26182_19_lrs2 : _GEN_5724; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5803 = 5'h13 == T_29096 ? T_26182_19_lrs3 : _GEN_5725; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5804 = 5'h13 == T_29096 ? T_26182_19_ldst_val : _GEN_5726; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5805 = 5'h13 == T_29096 ? T_26182_19_dst_rtype : _GEN_5727; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5806 = 5'h13 == T_29096 ? T_26182_19_lrs1_rtype : _GEN_5728; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5807 = 5'h13 == T_29096 ? T_26182_19_lrs2_rtype : _GEN_5729; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5808 = 5'h13 == T_29096 ? T_26182_19_frs3_en : _GEN_5730; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5809 = 5'h13 == T_29096 ? T_26182_19_fp_val : _GEN_5731; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5810 = 5'h13 == T_29096 ? T_26182_19_fp_single : _GEN_5732; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5811 = 5'h13 == T_29096 ? T_26182_19_xcpt_if : _GEN_5733; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5812 = 5'h13 == T_29096 ? T_26182_19_replay_if : _GEN_5734; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5814 = 5'h13 == T_29096 ? T_26182_19_debug_events_fetch_seq : _GEN_5736; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5815 = 5'h14 == T_29096 ? T_26182_20_valid : _GEN_5737; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5816 = 5'h14 == T_29096 ? T_26182_20_iw_state : _GEN_5738; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5817 = 5'h14 == T_29096 ? T_26182_20_uopc : _GEN_5739; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5818 = 5'h14 == T_29096 ? T_26182_20_inst : _GEN_5740; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5819 = 5'h14 == T_29096 ? T_26182_20_pc : _GEN_5741; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5820 = 5'h14 == T_29096 ? T_26182_20_fu_code : _GEN_5742; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5821 = 5'h14 == T_29096 ? T_26182_20_ctrl_br_type : _GEN_5743; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5822 = 5'h14 == T_29096 ? T_26182_20_ctrl_op1_sel : _GEN_5744; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5823 = 5'h14 == T_29096 ? T_26182_20_ctrl_op2_sel : _GEN_5745; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5824 = 5'h14 == T_29096 ? T_26182_20_ctrl_imm_sel : _GEN_5746; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5825 = 5'h14 == T_29096 ? T_26182_20_ctrl_op_fcn : _GEN_5747; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5826 = 5'h14 == T_29096 ? T_26182_20_ctrl_fcn_dw : _GEN_5748; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5827 = 5'h14 == T_29096 ? T_26182_20_ctrl_rf_wen : _GEN_5749; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5828 = 5'h14 == T_29096 ? T_26182_20_ctrl_csr_cmd : _GEN_5750; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5829 = 5'h14 == T_29096 ? T_26182_20_ctrl_is_load : _GEN_5751; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5830 = 5'h14 == T_29096 ? T_26182_20_ctrl_is_sta : _GEN_5752; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5831 = 5'h14 == T_29096 ? T_26182_20_ctrl_is_std : _GEN_5753; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5832 = 5'h14 == T_29096 ? T_26182_20_wakeup_delay : _GEN_5754; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5833 = 5'h14 == T_29096 ? T_26182_20_allocate_brtag : _GEN_5755; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5834 = 5'h14 == T_29096 ? T_26182_20_is_br_or_jmp : _GEN_5756; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5835 = 5'h14 == T_29096 ? T_26182_20_is_jump : _GEN_5757; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5836 = 5'h14 == T_29096 ? T_26182_20_is_jal : _GEN_5758; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5837 = 5'h14 == T_29096 ? T_26182_20_is_ret : _GEN_5759; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5838 = 5'h14 == T_29096 ? T_26182_20_is_call : _GEN_5760; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5839 = 5'h14 == T_29096 ? T_26182_20_br_mask : _GEN_5761; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5840 = 5'h14 == T_29096 ? T_26182_20_br_tag : _GEN_5762; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5841 = 5'h14 == T_29096 ? T_26182_20_br_prediction_bpd_predict_val : _GEN_5763; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5842 = 5'h14 == T_29096 ? T_26182_20_br_prediction_bpd_predict_taken : _GEN_5764; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5843 = 5'h14 == T_29096 ? T_26182_20_br_prediction_btb_hit : _GEN_5765; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5844 = 5'h14 == T_29096 ? T_26182_20_br_prediction_btb_predicted : _GEN_5766; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5845 = 5'h14 == T_29096 ? T_26182_20_br_prediction_is_br_or_jalr : _GEN_5767; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5846 = 5'h14 == T_29096 ? T_26182_20_stat_brjmp_mispredicted : _GEN_5768; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5847 = 5'h14 == T_29096 ? T_26182_20_stat_btb_made_pred : _GEN_5769; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5848 = 5'h14 == T_29096 ? T_26182_20_stat_btb_mispredicted : _GEN_5770; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5849 = 5'h14 == T_29096 ? T_26182_20_stat_bpd_made_pred : _GEN_5771; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5850 = 5'h14 == T_29096 ? T_26182_20_stat_bpd_mispredicted : _GEN_5772; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5851 = 5'h14 == T_29096 ? T_26182_20_fetch_pc_lob : _GEN_5773; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5852 = 5'h14 == T_29096 ? T_26182_20_imm_packed : _GEN_5774; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5853 = 5'h14 == T_29096 ? T_26182_20_csr_addr : _GEN_5775; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5854 = 5'h14 == T_29096 ? T_26182_20_rob_idx : _GEN_5776; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5855 = 5'h14 == T_29096 ? T_26182_20_ldq_idx : _GEN_5777; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5856 = 5'h14 == T_29096 ? T_26182_20_stq_idx : _GEN_5778; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5857 = 5'h14 == T_29096 ? T_26182_20_brob_idx : _GEN_5779; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5858 = 5'h14 == T_29096 ? T_26182_20_pdst : _GEN_5780; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5859 = 5'h14 == T_29096 ? T_26182_20_pop1 : _GEN_5781; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5860 = 5'h14 == T_29096 ? T_26182_20_pop2 : _GEN_5782; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5861 = 5'h14 == T_29096 ? T_26182_20_pop3 : _GEN_5783; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5862 = 5'h14 == T_29096 ? T_26182_20_prs1_busy : _GEN_5784; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5863 = 5'h14 == T_29096 ? T_26182_20_prs2_busy : _GEN_5785; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5864 = 5'h14 == T_29096 ? T_26182_20_prs3_busy : _GEN_5786; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5865 = 5'h14 == T_29096 ? T_26182_20_stale_pdst : _GEN_5787; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5866 = 5'h14 == T_29096 ? T_26182_20_exception : _GEN_5788; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5867 = 5'h14 == T_29096 ? T_26182_20_exc_cause : _GEN_5789; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5868 = 5'h14 == T_29096 ? T_26182_20_bypassable : _GEN_5790; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5869 = 5'h14 == T_29096 ? T_26182_20_mem_cmd : _GEN_5791; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5870 = 5'h14 == T_29096 ? T_26182_20_mem_typ : _GEN_5792; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5871 = 5'h14 == T_29096 ? T_26182_20_is_fence : _GEN_5793; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5872 = 5'h14 == T_29096 ? T_26182_20_is_fencei : _GEN_5794; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5873 = 5'h14 == T_29096 ? T_26182_20_is_store : _GEN_5795; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5874 = 5'h14 == T_29096 ? T_26182_20_is_amo : _GEN_5796; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5875 = 5'h14 == T_29096 ? T_26182_20_is_load : _GEN_5797; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5876 = 5'h14 == T_29096 ? T_26182_20_is_unique : _GEN_5798; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5877 = 5'h14 == T_29096 ? T_26182_20_flush_on_commit : _GEN_5799; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5878 = 5'h14 == T_29096 ? T_26182_20_ldst : _GEN_5800; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5879 = 5'h14 == T_29096 ? T_26182_20_lrs1 : _GEN_5801; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5880 = 5'h14 == T_29096 ? T_26182_20_lrs2 : _GEN_5802; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5881 = 5'h14 == T_29096 ? T_26182_20_lrs3 : _GEN_5803; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5882 = 5'h14 == T_29096 ? T_26182_20_ldst_val : _GEN_5804; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5883 = 5'h14 == T_29096 ? T_26182_20_dst_rtype : _GEN_5805; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5884 = 5'h14 == T_29096 ? T_26182_20_lrs1_rtype : _GEN_5806; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5885 = 5'h14 == T_29096 ? T_26182_20_lrs2_rtype : _GEN_5807; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5886 = 5'h14 == T_29096 ? T_26182_20_frs3_en : _GEN_5808; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5887 = 5'h14 == T_29096 ? T_26182_20_fp_val : _GEN_5809; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5888 = 5'h14 == T_29096 ? T_26182_20_fp_single : _GEN_5810; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5889 = 5'h14 == T_29096 ? T_26182_20_xcpt_if : _GEN_5811; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5890 = 5'h14 == T_29096 ? T_26182_20_replay_if : _GEN_5812; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5892 = 5'h14 == T_29096 ? T_26182_20_debug_events_fetch_seq : _GEN_5814; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5893 = 5'h15 == T_29096 ? T_26182_21_valid : _GEN_5815; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5894 = 5'h15 == T_29096 ? T_26182_21_iw_state : _GEN_5816; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5895 = 5'h15 == T_29096 ? T_26182_21_uopc : _GEN_5817; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5896 = 5'h15 == T_29096 ? T_26182_21_inst : _GEN_5818; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5897 = 5'h15 == T_29096 ? T_26182_21_pc : _GEN_5819; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5898 = 5'h15 == T_29096 ? T_26182_21_fu_code : _GEN_5820; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5899 = 5'h15 == T_29096 ? T_26182_21_ctrl_br_type : _GEN_5821; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5900 = 5'h15 == T_29096 ? T_26182_21_ctrl_op1_sel : _GEN_5822; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5901 = 5'h15 == T_29096 ? T_26182_21_ctrl_op2_sel : _GEN_5823; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5902 = 5'h15 == T_29096 ? T_26182_21_ctrl_imm_sel : _GEN_5824; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5903 = 5'h15 == T_29096 ? T_26182_21_ctrl_op_fcn : _GEN_5825; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5904 = 5'h15 == T_29096 ? T_26182_21_ctrl_fcn_dw : _GEN_5826; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5905 = 5'h15 == T_29096 ? T_26182_21_ctrl_rf_wen : _GEN_5827; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5906 = 5'h15 == T_29096 ? T_26182_21_ctrl_csr_cmd : _GEN_5828; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5907 = 5'h15 == T_29096 ? T_26182_21_ctrl_is_load : _GEN_5829; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5908 = 5'h15 == T_29096 ? T_26182_21_ctrl_is_sta : _GEN_5830; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5909 = 5'h15 == T_29096 ? T_26182_21_ctrl_is_std : _GEN_5831; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5910 = 5'h15 == T_29096 ? T_26182_21_wakeup_delay : _GEN_5832; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5911 = 5'h15 == T_29096 ? T_26182_21_allocate_brtag : _GEN_5833; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5912 = 5'h15 == T_29096 ? T_26182_21_is_br_or_jmp : _GEN_5834; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5913 = 5'h15 == T_29096 ? T_26182_21_is_jump : _GEN_5835; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5914 = 5'h15 == T_29096 ? T_26182_21_is_jal : _GEN_5836; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5915 = 5'h15 == T_29096 ? T_26182_21_is_ret : _GEN_5837; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5916 = 5'h15 == T_29096 ? T_26182_21_is_call : _GEN_5838; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5917 = 5'h15 == T_29096 ? T_26182_21_br_mask : _GEN_5839; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5918 = 5'h15 == T_29096 ? T_26182_21_br_tag : _GEN_5840; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5919 = 5'h15 == T_29096 ? T_26182_21_br_prediction_bpd_predict_val : _GEN_5841; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5920 = 5'h15 == T_29096 ? T_26182_21_br_prediction_bpd_predict_taken : _GEN_5842; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5921 = 5'h15 == T_29096 ? T_26182_21_br_prediction_btb_hit : _GEN_5843; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5922 = 5'h15 == T_29096 ? T_26182_21_br_prediction_btb_predicted : _GEN_5844; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5923 = 5'h15 == T_29096 ? T_26182_21_br_prediction_is_br_or_jalr : _GEN_5845; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5924 = 5'h15 == T_29096 ? T_26182_21_stat_brjmp_mispredicted : _GEN_5846; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5925 = 5'h15 == T_29096 ? T_26182_21_stat_btb_made_pred : _GEN_5847; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5926 = 5'h15 == T_29096 ? T_26182_21_stat_btb_mispredicted : _GEN_5848; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5927 = 5'h15 == T_29096 ? T_26182_21_stat_bpd_made_pred : _GEN_5849; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5928 = 5'h15 == T_29096 ? T_26182_21_stat_bpd_mispredicted : _GEN_5850; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5929 = 5'h15 == T_29096 ? T_26182_21_fetch_pc_lob : _GEN_5851; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_5930 = 5'h15 == T_29096 ? T_26182_21_imm_packed : _GEN_5852; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_5931 = 5'h15 == T_29096 ? T_26182_21_csr_addr : _GEN_5853; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5932 = 5'h15 == T_29096 ? T_26182_21_rob_idx : _GEN_5854; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5933 = 5'h15 == T_29096 ? T_26182_21_ldq_idx : _GEN_5855; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5934 = 5'h15 == T_29096 ? T_26182_21_stq_idx : _GEN_5856; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_5935 = 5'h15 == T_29096 ? T_26182_21_brob_idx : _GEN_5857; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5936 = 5'h15 == T_29096 ? T_26182_21_pdst : _GEN_5858; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5937 = 5'h15 == T_29096 ? T_26182_21_pop1 : _GEN_5859; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5938 = 5'h15 == T_29096 ? T_26182_21_pop2 : _GEN_5860; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5939 = 5'h15 == T_29096 ? T_26182_21_pop3 : _GEN_5861; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5940 = 5'h15 == T_29096 ? T_26182_21_prs1_busy : _GEN_5862; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5941 = 5'h15 == T_29096 ? T_26182_21_prs2_busy : _GEN_5863; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5942 = 5'h15 == T_29096 ? T_26182_21_prs3_busy : _GEN_5864; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_5943 = 5'h15 == T_29096 ? T_26182_21_stale_pdst : _GEN_5865; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5944 = 5'h15 == T_29096 ? T_26182_21_exception : _GEN_5866; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_5945 = 5'h15 == T_29096 ? T_26182_21_exc_cause : _GEN_5867; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5946 = 5'h15 == T_29096 ? T_26182_21_bypassable : _GEN_5868; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5947 = 5'h15 == T_29096 ? T_26182_21_mem_cmd : _GEN_5869; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5948 = 5'h15 == T_29096 ? T_26182_21_mem_typ : _GEN_5870; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5949 = 5'h15 == T_29096 ? T_26182_21_is_fence : _GEN_5871; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5950 = 5'h15 == T_29096 ? T_26182_21_is_fencei : _GEN_5872; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5951 = 5'h15 == T_29096 ? T_26182_21_is_store : _GEN_5873; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5952 = 5'h15 == T_29096 ? T_26182_21_is_amo : _GEN_5874; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5953 = 5'h15 == T_29096 ? T_26182_21_is_load : _GEN_5875; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5954 = 5'h15 == T_29096 ? T_26182_21_is_unique : _GEN_5876; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5955 = 5'h15 == T_29096 ? T_26182_21_flush_on_commit : _GEN_5877; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5956 = 5'h15 == T_29096 ? T_26182_21_ldst : _GEN_5878; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5957 = 5'h15 == T_29096 ? T_26182_21_lrs1 : _GEN_5879; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5958 = 5'h15 == T_29096 ? T_26182_21_lrs2 : _GEN_5880; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_5959 = 5'h15 == T_29096 ? T_26182_21_lrs3 : _GEN_5881; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5960 = 5'h15 == T_29096 ? T_26182_21_ldst_val : _GEN_5882; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5961 = 5'h15 == T_29096 ? T_26182_21_dst_rtype : _GEN_5883; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5962 = 5'h15 == T_29096 ? T_26182_21_lrs1_rtype : _GEN_5884; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5963 = 5'h15 == T_29096 ? T_26182_21_lrs2_rtype : _GEN_5885; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5964 = 5'h15 == T_29096 ? T_26182_21_frs3_en : _GEN_5886; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5965 = 5'h15 == T_29096 ? T_26182_21_fp_val : _GEN_5887; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5966 = 5'h15 == T_29096 ? T_26182_21_fp_single : _GEN_5888; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5967 = 5'h15 == T_29096 ? T_26182_21_xcpt_if : _GEN_5889; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5968 = 5'h15 == T_29096 ? T_26182_21_replay_if : _GEN_5890; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5970 = 5'h15 == T_29096 ? T_26182_21_debug_events_fetch_seq : _GEN_5892; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5971 = 5'h16 == T_29096 ? T_26182_22_valid : _GEN_5893; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5972 = 5'h16 == T_29096 ? T_26182_22_iw_state : _GEN_5894; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_5973 = 5'h16 == T_29096 ? T_26182_22_uopc : _GEN_5895; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_5974 = 5'h16 == T_29096 ? T_26182_22_inst : _GEN_5896; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_5975 = 5'h16 == T_29096 ? T_26182_22_pc : _GEN_5897; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5976 = 5'h16 == T_29096 ? T_26182_22_fu_code : _GEN_5898; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5977 = 5'h16 == T_29096 ? T_26182_22_ctrl_br_type : _GEN_5899; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5978 = 5'h16 == T_29096 ? T_26182_22_ctrl_op1_sel : _GEN_5900; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5979 = 5'h16 == T_29096 ? T_26182_22_ctrl_op2_sel : _GEN_5901; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5980 = 5'h16 == T_29096 ? T_26182_22_ctrl_imm_sel : _GEN_5902; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_5981 = 5'h16 == T_29096 ? T_26182_22_ctrl_op_fcn : _GEN_5903; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5982 = 5'h16 == T_29096 ? T_26182_22_ctrl_fcn_dw : _GEN_5904; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5983 = 5'h16 == T_29096 ? T_26182_22_ctrl_rf_wen : _GEN_5905; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5984 = 5'h16 == T_29096 ? T_26182_22_ctrl_csr_cmd : _GEN_5906; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5985 = 5'h16 == T_29096 ? T_26182_22_ctrl_is_load : _GEN_5907; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5986 = 5'h16 == T_29096 ? T_26182_22_ctrl_is_sta : _GEN_5908; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5987 = 5'h16 == T_29096 ? T_26182_22_ctrl_is_std : _GEN_5909; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_5988 = 5'h16 == T_29096 ? T_26182_22_wakeup_delay : _GEN_5910; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5989 = 5'h16 == T_29096 ? T_26182_22_allocate_brtag : _GEN_5911; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5990 = 5'h16 == T_29096 ? T_26182_22_is_br_or_jmp : _GEN_5912; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5991 = 5'h16 == T_29096 ? T_26182_22_is_jump : _GEN_5913; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5992 = 5'h16 == T_29096 ? T_26182_22_is_jal : _GEN_5914; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5993 = 5'h16 == T_29096 ? T_26182_22_is_ret : _GEN_5915; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5994 = 5'h16 == T_29096 ? T_26182_22_is_call : _GEN_5916; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_5995 = 5'h16 == T_29096 ? T_26182_22_br_mask : _GEN_5917; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_5996 = 5'h16 == T_29096 ? T_26182_22_br_tag : _GEN_5918; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5997 = 5'h16 == T_29096 ? T_26182_22_br_prediction_bpd_predict_val : _GEN_5919; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5998 = 5'h16 == T_29096 ? T_26182_22_br_prediction_bpd_predict_taken : _GEN_5920; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_5999 = 5'h16 == T_29096 ? T_26182_22_br_prediction_btb_hit : _GEN_5921; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6000 = 5'h16 == T_29096 ? T_26182_22_br_prediction_btb_predicted : _GEN_5922; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6001 = 5'h16 == T_29096 ? T_26182_22_br_prediction_is_br_or_jalr : _GEN_5923; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6002 = 5'h16 == T_29096 ? T_26182_22_stat_brjmp_mispredicted : _GEN_5924; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6003 = 5'h16 == T_29096 ? T_26182_22_stat_btb_made_pred : _GEN_5925; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6004 = 5'h16 == T_29096 ? T_26182_22_stat_btb_mispredicted : _GEN_5926; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6005 = 5'h16 == T_29096 ? T_26182_22_stat_bpd_made_pred : _GEN_5927; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6006 = 5'h16 == T_29096 ? T_26182_22_stat_bpd_mispredicted : _GEN_5928; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_6007 = 5'h16 == T_29096 ? T_26182_22_fetch_pc_lob : _GEN_5929; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_6008 = 5'h16 == T_29096 ? T_26182_22_imm_packed : _GEN_5930; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_6009 = 5'h16 == T_29096 ? T_26182_22_csr_addr : _GEN_5931; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_6010 = 5'h16 == T_29096 ? T_26182_22_rob_idx : _GEN_5932; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_6011 = 5'h16 == T_29096 ? T_26182_22_ldq_idx : _GEN_5933; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_6012 = 5'h16 == T_29096 ? T_26182_22_stq_idx : _GEN_5934; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_6013 = 5'h16 == T_29096 ? T_26182_22_brob_idx : _GEN_5935; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_6014 = 5'h16 == T_29096 ? T_26182_22_pdst : _GEN_5936; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_6015 = 5'h16 == T_29096 ? T_26182_22_pop1 : _GEN_5937; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_6016 = 5'h16 == T_29096 ? T_26182_22_pop2 : _GEN_5938; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_6017 = 5'h16 == T_29096 ? T_26182_22_pop3 : _GEN_5939; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6018 = 5'h16 == T_29096 ? T_26182_22_prs1_busy : _GEN_5940; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6019 = 5'h16 == T_29096 ? T_26182_22_prs2_busy : _GEN_5941; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6020 = 5'h16 == T_29096 ? T_26182_22_prs3_busy : _GEN_5942; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_6021 = 5'h16 == T_29096 ? T_26182_22_stale_pdst : _GEN_5943; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6022 = 5'h16 == T_29096 ? T_26182_22_exception : _GEN_5944; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_6023 = 5'h16 == T_29096 ? T_26182_22_exc_cause : _GEN_5945; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6024 = 5'h16 == T_29096 ? T_26182_22_bypassable : _GEN_5946; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_6025 = 5'h16 == T_29096 ? T_26182_22_mem_cmd : _GEN_5947; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_6026 = 5'h16 == T_29096 ? T_26182_22_mem_typ : _GEN_5948; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6027 = 5'h16 == T_29096 ? T_26182_22_is_fence : _GEN_5949; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6028 = 5'h16 == T_29096 ? T_26182_22_is_fencei : _GEN_5950; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6029 = 5'h16 == T_29096 ? T_26182_22_is_store : _GEN_5951; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6030 = 5'h16 == T_29096 ? T_26182_22_is_amo : _GEN_5952; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6031 = 5'h16 == T_29096 ? T_26182_22_is_load : _GEN_5953; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6032 = 5'h16 == T_29096 ? T_26182_22_is_unique : _GEN_5954; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6033 = 5'h16 == T_29096 ? T_26182_22_flush_on_commit : _GEN_5955; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_6034 = 5'h16 == T_29096 ? T_26182_22_ldst : _GEN_5956; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_6035 = 5'h16 == T_29096 ? T_26182_22_lrs1 : _GEN_5957; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_6036 = 5'h16 == T_29096 ? T_26182_22_lrs2 : _GEN_5958; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_6037 = 5'h16 == T_29096 ? T_26182_22_lrs3 : _GEN_5959; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6038 = 5'h16 == T_29096 ? T_26182_22_ldst_val : _GEN_5960; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_6039 = 5'h16 == T_29096 ? T_26182_22_dst_rtype : _GEN_5961; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_6040 = 5'h16 == T_29096 ? T_26182_22_lrs1_rtype : _GEN_5962; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_6041 = 5'h16 == T_29096 ? T_26182_22_lrs2_rtype : _GEN_5963; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6042 = 5'h16 == T_29096 ? T_26182_22_frs3_en : _GEN_5964; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6043 = 5'h16 == T_29096 ? T_26182_22_fp_val : _GEN_5965; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6044 = 5'h16 == T_29096 ? T_26182_22_fp_single : _GEN_5966; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6045 = 5'h16 == T_29096 ? T_26182_22_xcpt_if : _GEN_5967; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_6046 = 5'h16 == T_29096 ? T_26182_22_replay_if : _GEN_5968; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_6048 = 5'h16 == T_29096 ? T_26182_22_debug_events_fetch_seq : _GEN_5970; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_6117 = 5'h17 == T_29096 ? T_26182_23_dst_rtype : _GEN_6039; // @[rob.scala 453:59 rob.scala 453:59]
  wire  T_29185 = _GEN_6117 == 2'h0; // @[rob.scala 453:59]
  wire  T_29271 = _GEN_6117 == 2'h1; // @[rob.scala 453:100]
  wire  T_29272 = T_29185 | T_29271; // @[rob.scala 453:70]
  wire  _GEN_6127 = 5'h0 == T_29096 ? 1'h0 : _GEN_1953; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6128 = 5'h1 == T_29096 ? 1'h0 : _GEN_1954; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6129 = 5'h2 == T_29096 ? 1'h0 : _GEN_1955; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6130 = 5'h3 == T_29096 ? 1'h0 : _GEN_1956; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6131 = 5'h4 == T_29096 ? 1'h0 : _GEN_1957; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6132 = 5'h5 == T_29096 ? 1'h0 : _GEN_1958; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6133 = 5'h6 == T_29096 ? 1'h0 : _GEN_1959; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6134 = 5'h7 == T_29096 ? 1'h0 : _GEN_1960; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6135 = 5'h8 == T_29096 ? 1'h0 : _GEN_1961; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6136 = 5'h9 == T_29096 ? 1'h0 : _GEN_1962; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6137 = 5'ha == T_29096 ? 1'h0 : _GEN_1963; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6138 = 5'hb == T_29096 ? 1'h0 : _GEN_1964; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6139 = 5'hc == T_29096 ? 1'h0 : _GEN_1965; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6140 = 5'hd == T_29096 ? 1'h0 : _GEN_1966; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6141 = 5'he == T_29096 ? 1'h0 : _GEN_1967; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6142 = 5'hf == T_29096 ? 1'h0 : _GEN_1968; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6143 = 5'h10 == T_29096 ? 1'h0 : _GEN_1969; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6144 = 5'h11 == T_29096 ? 1'h0 : _GEN_1970; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6145 = 5'h12 == T_29096 ? 1'h0 : _GEN_1971; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6146 = 5'h13 == T_29096 ? 1'h0 : _GEN_1972; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6147 = 5'h14 == T_29096 ? 1'h0 : _GEN_1973; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6148 = 5'h15 == T_29096 ? 1'h0 : _GEN_1974; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6149 = 5'h16 == T_29096 ? 1'h0 : _GEN_1975; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6150 = 5'h17 == T_29096 ? 1'h0 : _GEN_1976; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_6151 = T_29097 ? _GEN_6127 : _GEN_1953; // @[rob.scala 458:7]
  wire  _GEN_6152 = T_29097 ? _GEN_6128 : _GEN_1954; // @[rob.scala 458:7]
  wire  _GEN_6153 = T_29097 ? _GEN_6129 : _GEN_1955; // @[rob.scala 458:7]
  wire  _GEN_6154 = T_29097 ? _GEN_6130 : _GEN_1956; // @[rob.scala 458:7]
  wire  _GEN_6155 = T_29097 ? _GEN_6131 : _GEN_1957; // @[rob.scala 458:7]
  wire  _GEN_6156 = T_29097 ? _GEN_6132 : _GEN_1958; // @[rob.scala 458:7]
  wire  _GEN_6157 = T_29097 ? _GEN_6133 : _GEN_1959; // @[rob.scala 458:7]
  wire  _GEN_6158 = T_29097 ? _GEN_6134 : _GEN_1960; // @[rob.scala 458:7]
  wire  _GEN_6159 = T_29097 ? _GEN_6135 : _GEN_1961; // @[rob.scala 458:7]
  wire  _GEN_6160 = T_29097 ? _GEN_6136 : _GEN_1962; // @[rob.scala 458:7]
  wire  _GEN_6161 = T_29097 ? _GEN_6137 : _GEN_1963; // @[rob.scala 458:7]
  wire  _GEN_6162 = T_29097 ? _GEN_6138 : _GEN_1964; // @[rob.scala 458:7]
  wire  _GEN_6163 = T_29097 ? _GEN_6139 : _GEN_1965; // @[rob.scala 458:7]
  wire  _GEN_6164 = T_29097 ? _GEN_6140 : _GEN_1966; // @[rob.scala 458:7]
  wire  _GEN_6165 = T_29097 ? _GEN_6141 : _GEN_1967; // @[rob.scala 458:7]
  wire  _GEN_6166 = T_29097 ? _GEN_6142 : _GEN_1968; // @[rob.scala 458:7]
  wire  _GEN_6167 = T_29097 ? _GEN_6143 : _GEN_1969; // @[rob.scala 458:7]
  wire  _GEN_6168 = T_29097 ? _GEN_6144 : _GEN_1970; // @[rob.scala 458:7]
  wire  _GEN_6169 = T_29097 ? _GEN_6145 : _GEN_1971; // @[rob.scala 458:7]
  wire  _GEN_6170 = T_29097 ? _GEN_6146 : _GEN_1972; // @[rob.scala 458:7]
  wire  _GEN_6171 = T_29097 ? _GEN_6147 : _GEN_1973; // @[rob.scala 458:7]
  wire  _GEN_6172 = T_29097 ? _GEN_6148 : _GEN_1974; // @[rob.scala 458:7]
  wire  _GEN_6173 = T_29097 ? _GEN_6149 : _GEN_1975; // @[rob.scala 458:7]
  wire  _GEN_6174 = T_29097 ? _GEN_6150 : _GEN_1976; // @[rob.scala 458:7]
  wire [7:0] T_29365 = io_brinfo_mask & T_26182_0_br_mask; // @[util.scala 45:52]
  wire  T_29367 = T_29365 != 8'h0; // @[util.scala 45:60]
  wire  T_29368 = T_23706_0 & T_29367; // @[rob.scala 481:39]
  wire  T_29369 = io_brinfo_valid & io_brinfo_mispredict; // @[rob.scala 484:32]
  wire  T_29370 = T_29369 & T_29368; // @[rob.scala 484:56]
  wire  _GEN_6180 = T_29370 ? 1'h0 : _GEN_6151; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6181 = T_29370 ? 32'h4033 : _GEN_3904; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_29459 = ~io_brinfo_mispredict; // @[rob.scala 489:40]
  wire  T_29460 = io_brinfo_valid & T_29459; // @[rob.scala 489:37]
  wire  T_29461 = T_29460 & T_29368; // @[rob.scala 489:62]
  wire  T_29463 = ~T_29370; // @[rob.scala 485:10]
  wire  T_29464 = T_29463 & T_29461; // @[rob.scala 490:10]
  wire [7:0] T_29465 = ~io_brinfo_mask; // @[rob.scala 492:46]
  wire [7:0] T_29466 = T_26182_0_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_29467 = io_brinfo_mask & T_26182_1_br_mask; // @[util.scala 45:52]
  wire  T_29469 = T_29467 != 8'h0; // @[util.scala 45:60]
  wire  T_29470 = T_23706_1 & T_29469; // @[rob.scala 481:39]
  wire  T_29472 = T_29369 & T_29470; // @[rob.scala 484:56]
  wire  _GEN_6183 = T_29472 ? 1'h0 : _GEN_6152; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6184 = T_29472 ? 32'h4033 : _GEN_3905; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_29563 = T_29460 & T_29470; // @[rob.scala 489:62]
  wire  T_29565 = ~T_29472; // @[rob.scala 485:10]
  wire  T_29566 = T_29565 & T_29563; // @[rob.scala 490:10]
  wire [7:0] T_29568 = T_26182_1_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_29569 = io_brinfo_mask & T_26182_2_br_mask; // @[util.scala 45:52]
  wire  T_29571 = T_29569 != 8'h0; // @[util.scala 45:60]
  wire  T_29572 = T_23706_2 & T_29571; // @[rob.scala 481:39]
  wire  T_29574 = T_29369 & T_29572; // @[rob.scala 484:56]
  wire  _GEN_6186 = T_29574 ? 1'h0 : _GEN_6153; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6187 = T_29574 ? 32'h4033 : _GEN_3906; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_29665 = T_29460 & T_29572; // @[rob.scala 489:62]
  wire  T_29667 = ~T_29574; // @[rob.scala 485:10]
  wire  T_29668 = T_29667 & T_29665; // @[rob.scala 490:10]
  wire [7:0] T_29670 = T_26182_2_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_29671 = io_brinfo_mask & T_26182_3_br_mask; // @[util.scala 45:52]
  wire  T_29673 = T_29671 != 8'h0; // @[util.scala 45:60]
  wire  T_29674 = T_23706_3 & T_29673; // @[rob.scala 481:39]
  wire  T_29676 = T_29369 & T_29674; // @[rob.scala 484:56]
  wire  _GEN_6189 = T_29676 ? 1'h0 : _GEN_6154; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6190 = T_29676 ? 32'h4033 : _GEN_3907; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_29767 = T_29460 & T_29674; // @[rob.scala 489:62]
  wire  T_29769 = ~T_29676; // @[rob.scala 485:10]
  wire  T_29770 = T_29769 & T_29767; // @[rob.scala 490:10]
  wire [7:0] T_29772 = T_26182_3_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_29773 = io_brinfo_mask & T_26182_4_br_mask; // @[util.scala 45:52]
  wire  T_29775 = T_29773 != 8'h0; // @[util.scala 45:60]
  wire  T_29776 = T_23706_4 & T_29775; // @[rob.scala 481:39]
  wire  T_29778 = T_29369 & T_29776; // @[rob.scala 484:56]
  wire  _GEN_6192 = T_29778 ? 1'h0 : _GEN_6155; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6193 = T_29778 ? 32'h4033 : _GEN_3908; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_29869 = T_29460 & T_29776; // @[rob.scala 489:62]
  wire  T_29871 = ~T_29778; // @[rob.scala 485:10]
  wire  T_29872 = T_29871 & T_29869; // @[rob.scala 490:10]
  wire [7:0] T_29874 = T_26182_4_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_29875 = io_brinfo_mask & T_26182_5_br_mask; // @[util.scala 45:52]
  wire  T_29877 = T_29875 != 8'h0; // @[util.scala 45:60]
  wire  T_29878 = T_23706_5 & T_29877; // @[rob.scala 481:39]
  wire  T_29880 = T_29369 & T_29878; // @[rob.scala 484:56]
  wire  _GEN_6195 = T_29880 ? 1'h0 : _GEN_6156; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6196 = T_29880 ? 32'h4033 : _GEN_3909; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_29971 = T_29460 & T_29878; // @[rob.scala 489:62]
  wire  T_29973 = ~T_29880; // @[rob.scala 485:10]
  wire  T_29974 = T_29973 & T_29971; // @[rob.scala 490:10]
  wire [7:0] T_29976 = T_26182_5_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_29977 = io_brinfo_mask & T_26182_6_br_mask; // @[util.scala 45:52]
  wire  T_29979 = T_29977 != 8'h0; // @[util.scala 45:60]
  wire  T_29980 = T_23706_6 & T_29979; // @[rob.scala 481:39]
  wire  T_29982 = T_29369 & T_29980; // @[rob.scala 484:56]
  wire  _GEN_6198 = T_29982 ? 1'h0 : _GEN_6157; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6199 = T_29982 ? 32'h4033 : _GEN_3910; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30073 = T_29460 & T_29980; // @[rob.scala 489:62]
  wire  T_30075 = ~T_29982; // @[rob.scala 485:10]
  wire  T_30076 = T_30075 & T_30073; // @[rob.scala 490:10]
  wire [7:0] T_30078 = T_26182_6_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30079 = io_brinfo_mask & T_26182_7_br_mask; // @[util.scala 45:52]
  wire  T_30081 = T_30079 != 8'h0; // @[util.scala 45:60]
  wire  T_30082 = T_23706_7 & T_30081; // @[rob.scala 481:39]
  wire  T_30084 = T_29369 & T_30082; // @[rob.scala 484:56]
  wire  _GEN_6201 = T_30084 ? 1'h0 : _GEN_6158; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6202 = T_30084 ? 32'h4033 : _GEN_3911; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30175 = T_29460 & T_30082; // @[rob.scala 489:62]
  wire  T_30177 = ~T_30084; // @[rob.scala 485:10]
  wire  T_30178 = T_30177 & T_30175; // @[rob.scala 490:10]
  wire [7:0] T_30180 = T_26182_7_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30181 = io_brinfo_mask & T_26182_8_br_mask; // @[util.scala 45:52]
  wire  T_30183 = T_30181 != 8'h0; // @[util.scala 45:60]
  wire  T_30184 = T_23706_8 & T_30183; // @[rob.scala 481:39]
  wire  T_30186 = T_29369 & T_30184; // @[rob.scala 484:56]
  wire  _GEN_6204 = T_30186 ? 1'h0 : _GEN_6159; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6205 = T_30186 ? 32'h4033 : _GEN_3912; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30277 = T_29460 & T_30184; // @[rob.scala 489:62]
  wire  T_30279 = ~T_30186; // @[rob.scala 485:10]
  wire  T_30280 = T_30279 & T_30277; // @[rob.scala 490:10]
  wire [7:0] T_30282 = T_26182_8_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30283 = io_brinfo_mask & T_26182_9_br_mask; // @[util.scala 45:52]
  wire  T_30285 = T_30283 != 8'h0; // @[util.scala 45:60]
  wire  T_30286 = T_23706_9 & T_30285; // @[rob.scala 481:39]
  wire  T_30288 = T_29369 & T_30286; // @[rob.scala 484:56]
  wire  _GEN_6207 = T_30288 ? 1'h0 : _GEN_6160; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6208 = T_30288 ? 32'h4033 : _GEN_3913; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30379 = T_29460 & T_30286; // @[rob.scala 489:62]
  wire  T_30381 = ~T_30288; // @[rob.scala 485:10]
  wire  T_30382 = T_30381 & T_30379; // @[rob.scala 490:10]
  wire [7:0] T_30384 = T_26182_9_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30385 = io_brinfo_mask & T_26182_10_br_mask; // @[util.scala 45:52]
  wire  T_30387 = T_30385 != 8'h0; // @[util.scala 45:60]
  wire  T_30388 = T_23706_10 & T_30387; // @[rob.scala 481:39]
  wire  T_30390 = T_29369 & T_30388; // @[rob.scala 484:56]
  wire  _GEN_6210 = T_30390 ? 1'h0 : _GEN_6161; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6211 = T_30390 ? 32'h4033 : _GEN_3914; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30481 = T_29460 & T_30388; // @[rob.scala 489:62]
  wire  T_30483 = ~T_30390; // @[rob.scala 485:10]
  wire  T_30484 = T_30483 & T_30481; // @[rob.scala 490:10]
  wire [7:0] T_30486 = T_26182_10_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30487 = io_brinfo_mask & T_26182_11_br_mask; // @[util.scala 45:52]
  wire  T_30489 = T_30487 != 8'h0; // @[util.scala 45:60]
  wire  T_30490 = T_23706_11 & T_30489; // @[rob.scala 481:39]
  wire  T_30492 = T_29369 & T_30490; // @[rob.scala 484:56]
  wire  _GEN_6213 = T_30492 ? 1'h0 : _GEN_6162; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6214 = T_30492 ? 32'h4033 : _GEN_3915; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30583 = T_29460 & T_30490; // @[rob.scala 489:62]
  wire  T_30585 = ~T_30492; // @[rob.scala 485:10]
  wire  T_30586 = T_30585 & T_30583; // @[rob.scala 490:10]
  wire [7:0] T_30588 = T_26182_11_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30589 = io_brinfo_mask & T_26182_12_br_mask; // @[util.scala 45:52]
  wire  T_30591 = T_30589 != 8'h0; // @[util.scala 45:60]
  wire  T_30592 = T_23706_12 & T_30591; // @[rob.scala 481:39]
  wire  T_30594 = T_29369 & T_30592; // @[rob.scala 484:56]
  wire  _GEN_6216 = T_30594 ? 1'h0 : _GEN_6163; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6217 = T_30594 ? 32'h4033 : _GEN_3916; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30685 = T_29460 & T_30592; // @[rob.scala 489:62]
  wire  T_30687 = ~T_30594; // @[rob.scala 485:10]
  wire  T_30688 = T_30687 & T_30685; // @[rob.scala 490:10]
  wire [7:0] T_30690 = T_26182_12_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30691 = io_brinfo_mask & T_26182_13_br_mask; // @[util.scala 45:52]
  wire  T_30693 = T_30691 != 8'h0; // @[util.scala 45:60]
  wire  T_30694 = T_23706_13 & T_30693; // @[rob.scala 481:39]
  wire  T_30696 = T_29369 & T_30694; // @[rob.scala 484:56]
  wire  _GEN_6219 = T_30696 ? 1'h0 : _GEN_6164; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6220 = T_30696 ? 32'h4033 : _GEN_3917; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30787 = T_29460 & T_30694; // @[rob.scala 489:62]
  wire  T_30789 = ~T_30696; // @[rob.scala 485:10]
  wire  T_30790 = T_30789 & T_30787; // @[rob.scala 490:10]
  wire [7:0] T_30792 = T_26182_13_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30793 = io_brinfo_mask & T_26182_14_br_mask; // @[util.scala 45:52]
  wire  T_30795 = T_30793 != 8'h0; // @[util.scala 45:60]
  wire  T_30796 = T_23706_14 & T_30795; // @[rob.scala 481:39]
  wire  T_30798 = T_29369 & T_30796; // @[rob.scala 484:56]
  wire  _GEN_6222 = T_30798 ? 1'h0 : _GEN_6165; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6223 = T_30798 ? 32'h4033 : _GEN_3918; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30889 = T_29460 & T_30796; // @[rob.scala 489:62]
  wire  T_30891 = ~T_30798; // @[rob.scala 485:10]
  wire  T_30892 = T_30891 & T_30889; // @[rob.scala 490:10]
  wire [7:0] T_30894 = T_26182_14_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30895 = io_brinfo_mask & T_26182_15_br_mask; // @[util.scala 45:52]
  wire  T_30897 = T_30895 != 8'h0; // @[util.scala 45:60]
  wire  T_30898 = T_23706_15 & T_30897; // @[rob.scala 481:39]
  wire  T_30900 = T_29369 & T_30898; // @[rob.scala 484:56]
  wire  _GEN_6225 = T_30900 ? 1'h0 : _GEN_6166; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6226 = T_30900 ? 32'h4033 : _GEN_3919; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_30991 = T_29460 & T_30898; // @[rob.scala 489:62]
  wire  T_30993 = ~T_30900; // @[rob.scala 485:10]
  wire  T_30994 = T_30993 & T_30991; // @[rob.scala 490:10]
  wire [7:0] T_30996 = T_26182_15_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_30997 = io_brinfo_mask & T_26182_16_br_mask; // @[util.scala 45:52]
  wire  T_30999 = T_30997 != 8'h0; // @[util.scala 45:60]
  wire  T_31000 = T_23706_16 & T_30999; // @[rob.scala 481:39]
  wire  T_31002 = T_29369 & T_31000; // @[rob.scala 484:56]
  wire  _GEN_6228 = T_31002 ? 1'h0 : _GEN_6167; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6229 = T_31002 ? 32'h4033 : _GEN_3920; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31093 = T_29460 & T_31000; // @[rob.scala 489:62]
  wire  T_31095 = ~T_31002; // @[rob.scala 485:10]
  wire  T_31096 = T_31095 & T_31093; // @[rob.scala 490:10]
  wire [7:0] T_31098 = T_26182_16_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31099 = io_brinfo_mask & T_26182_17_br_mask; // @[util.scala 45:52]
  wire  T_31101 = T_31099 != 8'h0; // @[util.scala 45:60]
  wire  T_31102 = T_23706_17 & T_31101; // @[rob.scala 481:39]
  wire  T_31104 = T_29369 & T_31102; // @[rob.scala 484:56]
  wire  _GEN_6231 = T_31104 ? 1'h0 : _GEN_6168; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6232 = T_31104 ? 32'h4033 : _GEN_3921; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31195 = T_29460 & T_31102; // @[rob.scala 489:62]
  wire  T_31197 = ~T_31104; // @[rob.scala 485:10]
  wire  T_31198 = T_31197 & T_31195; // @[rob.scala 490:10]
  wire [7:0] T_31200 = T_26182_17_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31201 = io_brinfo_mask & T_26182_18_br_mask; // @[util.scala 45:52]
  wire  T_31203 = T_31201 != 8'h0; // @[util.scala 45:60]
  wire  T_31204 = T_23706_18 & T_31203; // @[rob.scala 481:39]
  wire  T_31206 = T_29369 & T_31204; // @[rob.scala 484:56]
  wire  _GEN_6234 = T_31206 ? 1'h0 : _GEN_6169; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6235 = T_31206 ? 32'h4033 : _GEN_3922; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31297 = T_29460 & T_31204; // @[rob.scala 489:62]
  wire  T_31299 = ~T_31206; // @[rob.scala 485:10]
  wire  T_31300 = T_31299 & T_31297; // @[rob.scala 490:10]
  wire [7:0] T_31302 = T_26182_18_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31303 = io_brinfo_mask & T_26182_19_br_mask; // @[util.scala 45:52]
  wire  T_31305 = T_31303 != 8'h0; // @[util.scala 45:60]
  wire  T_31306 = T_23706_19 & T_31305; // @[rob.scala 481:39]
  wire  T_31308 = T_29369 & T_31306; // @[rob.scala 484:56]
  wire  _GEN_6237 = T_31308 ? 1'h0 : _GEN_6170; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6238 = T_31308 ? 32'h4033 : _GEN_3923; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31399 = T_29460 & T_31306; // @[rob.scala 489:62]
  wire  T_31401 = ~T_31308; // @[rob.scala 485:10]
  wire  T_31402 = T_31401 & T_31399; // @[rob.scala 490:10]
  wire [7:0] T_31404 = T_26182_19_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31405 = io_brinfo_mask & T_26182_20_br_mask; // @[util.scala 45:52]
  wire  T_31407 = T_31405 != 8'h0; // @[util.scala 45:60]
  wire  T_31408 = T_23706_20 & T_31407; // @[rob.scala 481:39]
  wire  T_31410 = T_29369 & T_31408; // @[rob.scala 484:56]
  wire  _GEN_6240 = T_31410 ? 1'h0 : _GEN_6171; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6241 = T_31410 ? 32'h4033 : _GEN_3924; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31501 = T_29460 & T_31408; // @[rob.scala 489:62]
  wire  T_31503 = ~T_31410; // @[rob.scala 485:10]
  wire  T_31504 = T_31503 & T_31501; // @[rob.scala 490:10]
  wire [7:0] T_31506 = T_26182_20_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31507 = io_brinfo_mask & T_26182_21_br_mask; // @[util.scala 45:52]
  wire  T_31509 = T_31507 != 8'h0; // @[util.scala 45:60]
  wire  T_31510 = T_23706_21 & T_31509; // @[rob.scala 481:39]
  wire  T_31512 = T_29369 & T_31510; // @[rob.scala 484:56]
  wire  _GEN_6243 = T_31512 ? 1'h0 : _GEN_6172; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6244 = T_31512 ? 32'h4033 : _GEN_3925; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31603 = T_29460 & T_31510; // @[rob.scala 489:62]
  wire  T_31605 = ~T_31512; // @[rob.scala 485:10]
  wire  T_31606 = T_31605 & T_31603; // @[rob.scala 490:10]
  wire [7:0] T_31608 = T_26182_21_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31609 = io_brinfo_mask & T_26182_22_br_mask; // @[util.scala 45:52]
  wire  T_31611 = T_31609 != 8'h0; // @[util.scala 45:60]
  wire  T_31612 = T_23706_22 & T_31611; // @[rob.scala 481:39]
  wire  T_31614 = T_29369 & T_31612; // @[rob.scala 484:56]
  wire  _GEN_6246 = T_31614 ? 1'h0 : _GEN_6173; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6247 = T_31614 ? 32'h4033 : _GEN_3926; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31705 = T_29460 & T_31612; // @[rob.scala 489:62]
  wire  T_31707 = ~T_31614; // @[rob.scala 485:10]
  wire  T_31708 = T_31707 & T_31705; // @[rob.scala 490:10]
  wire [7:0] T_31710 = T_26182_22_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_31711 = io_brinfo_mask & T_26182_23_br_mask; // @[util.scala 45:52]
  wire  T_31713 = T_31711 != 8'h0; // @[util.scala 45:60]
  wire  T_31714 = T_23706_23 & T_31713; // @[rob.scala 481:39]
  wire  T_31716 = T_29369 & T_31714; // @[rob.scala 484:56]
  wire  _GEN_6249 = T_31716 ? 1'h0 : _GEN_6174; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_6250 = T_31716 ? 32'h4033 : _GEN_3927; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_31807 = T_29460 & T_31714; // @[rob.scala 489:62]
  wire  T_31809 = ~T_31716; // @[rob.scala 485:10]
  wire  T_31810 = T_31809 & T_31807; // @[rob.scala 490:10]
  wire [7:0] T_31812 = T_26182_23_br_mask & T_29465; // @[rob.scala 492:44]
  wire  _GEN_6436 = 5'h1 == rob_head ? T_26182_1_is_store : T_26182_0_is_store; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6438 = 5'h1 == rob_head ? T_26182_1_is_load : T_26182_0_is_load; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6454 = 5'h1 == rob_head ? T_26182_1_debug_wdata : T_26182_0_debug_wdata; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6514 = 5'h2 == rob_head ? T_26182_2_is_store : _GEN_6436; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6516 = 5'h2 == rob_head ? T_26182_2_is_load : _GEN_6438; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6532 = 5'h2 == rob_head ? T_26182_2_debug_wdata : _GEN_6454; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6592 = 5'h3 == rob_head ? T_26182_3_is_store : _GEN_6514; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6594 = 5'h3 == rob_head ? T_26182_3_is_load : _GEN_6516; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6610 = 5'h3 == rob_head ? T_26182_3_debug_wdata : _GEN_6532; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6670 = 5'h4 == rob_head ? T_26182_4_is_store : _GEN_6592; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6672 = 5'h4 == rob_head ? T_26182_4_is_load : _GEN_6594; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6688 = 5'h4 == rob_head ? T_26182_4_debug_wdata : _GEN_6610; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6748 = 5'h5 == rob_head ? T_26182_5_is_store : _GEN_6670; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6750 = 5'h5 == rob_head ? T_26182_5_is_load : _GEN_6672; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6766 = 5'h5 == rob_head ? T_26182_5_debug_wdata : _GEN_6688; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6826 = 5'h6 == rob_head ? T_26182_6_is_store : _GEN_6748; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6828 = 5'h6 == rob_head ? T_26182_6_is_load : _GEN_6750; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6844 = 5'h6 == rob_head ? T_26182_6_debug_wdata : _GEN_6766; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6904 = 5'h7 == rob_head ? T_26182_7_is_store : _GEN_6826; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6906 = 5'h7 == rob_head ? T_26182_7_is_load : _GEN_6828; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_6922 = 5'h7 == rob_head ? T_26182_7_debug_wdata : _GEN_6844; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6982 = 5'h8 == rob_head ? T_26182_8_is_store : _GEN_6904; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_6984 = 5'h8 == rob_head ? T_26182_8_is_load : _GEN_6906; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7000 = 5'h8 == rob_head ? T_26182_8_debug_wdata : _GEN_6922; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7060 = 5'h9 == rob_head ? T_26182_9_is_store : _GEN_6982; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7062 = 5'h9 == rob_head ? T_26182_9_is_load : _GEN_6984; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7078 = 5'h9 == rob_head ? T_26182_9_debug_wdata : _GEN_7000; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7138 = 5'ha == rob_head ? T_26182_10_is_store : _GEN_7060; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7140 = 5'ha == rob_head ? T_26182_10_is_load : _GEN_7062; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7156 = 5'ha == rob_head ? T_26182_10_debug_wdata : _GEN_7078; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7216 = 5'hb == rob_head ? T_26182_11_is_store : _GEN_7138; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7218 = 5'hb == rob_head ? T_26182_11_is_load : _GEN_7140; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7234 = 5'hb == rob_head ? T_26182_11_debug_wdata : _GEN_7156; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7294 = 5'hc == rob_head ? T_26182_12_is_store : _GEN_7216; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7296 = 5'hc == rob_head ? T_26182_12_is_load : _GEN_7218; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7312 = 5'hc == rob_head ? T_26182_12_debug_wdata : _GEN_7234; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7372 = 5'hd == rob_head ? T_26182_13_is_store : _GEN_7294; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7374 = 5'hd == rob_head ? T_26182_13_is_load : _GEN_7296; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7390 = 5'hd == rob_head ? T_26182_13_debug_wdata : _GEN_7312; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7450 = 5'he == rob_head ? T_26182_14_is_store : _GEN_7372; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7452 = 5'he == rob_head ? T_26182_14_is_load : _GEN_7374; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7468 = 5'he == rob_head ? T_26182_14_debug_wdata : _GEN_7390; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7528 = 5'hf == rob_head ? T_26182_15_is_store : _GEN_7450; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7530 = 5'hf == rob_head ? T_26182_15_is_load : _GEN_7452; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7546 = 5'hf == rob_head ? T_26182_15_debug_wdata : _GEN_7468; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7606 = 5'h10 == rob_head ? T_26182_16_is_store : _GEN_7528; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7608 = 5'h10 == rob_head ? T_26182_16_is_load : _GEN_7530; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7624 = 5'h10 == rob_head ? T_26182_16_debug_wdata : _GEN_7546; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7684 = 5'h11 == rob_head ? T_26182_17_is_store : _GEN_7606; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7686 = 5'h11 == rob_head ? T_26182_17_is_load : _GEN_7608; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7702 = 5'h11 == rob_head ? T_26182_17_debug_wdata : _GEN_7624; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7762 = 5'h12 == rob_head ? T_26182_18_is_store : _GEN_7684; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7764 = 5'h12 == rob_head ? T_26182_18_is_load : _GEN_7686; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7780 = 5'h12 == rob_head ? T_26182_18_debug_wdata : _GEN_7702; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7840 = 5'h13 == rob_head ? T_26182_19_is_store : _GEN_7762; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7842 = 5'h13 == rob_head ? T_26182_19_is_load : _GEN_7764; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7858 = 5'h13 == rob_head ? T_26182_19_debug_wdata : _GEN_7780; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7918 = 5'h14 == rob_head ? T_26182_20_is_store : _GEN_7840; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7920 = 5'h14 == rob_head ? T_26182_20_is_load : _GEN_7842; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_7936 = 5'h14 == rob_head ? T_26182_20_debug_wdata : _GEN_7858; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7996 = 5'h15 == rob_head ? T_26182_21_is_store : _GEN_7918; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_7998 = 5'h15 == rob_head ? T_26182_21_is_load : _GEN_7920; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_8014 = 5'h15 == rob_head ? T_26182_21_debug_wdata : _GEN_7936; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_8074 = 5'h16 == rob_head ? T_26182_22_is_store : _GEN_7996; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_8076 = 5'h16 == rob_head ? T_26182_22_is_load : _GEN_7998; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_8092 = 5'h16 == rob_head ? T_26182_22_debug_wdata : _GEN_8014; // @[rob.scala 507:28 rob.scala 507:28]
  wire  rob_head_is_store_0 = 5'h17 == rob_head ? T_26182_23_is_store : _GEN_8074; // @[rob.scala 507:28 rob.scala 507:28]
  wire  rob_head_is_load_0 = 5'h17 == rob_head ? T_26182_23_is_load : _GEN_8076; // @[rob.scala 507:28 rob.scala 507:28]
  wire [31:0] _GEN_8196 = 5'h0 == rob_head ? 32'h4033 : _GEN_6181; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8197 = 5'h1 == rob_head ? 32'h4033 : _GEN_6184; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8198 = 5'h2 == rob_head ? 32'h4033 : _GEN_6187; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8199 = 5'h3 == rob_head ? 32'h4033 : _GEN_6190; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8200 = 5'h4 == rob_head ? 32'h4033 : _GEN_6193; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8201 = 5'h5 == rob_head ? 32'h4033 : _GEN_6196; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8202 = 5'h6 == rob_head ? 32'h4033 : _GEN_6199; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8203 = 5'h7 == rob_head ? 32'h4033 : _GEN_6202; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8204 = 5'h8 == rob_head ? 32'h4033 : _GEN_6205; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8205 = 5'h9 == rob_head ? 32'h4033 : _GEN_6208; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8206 = 5'ha == rob_head ? 32'h4033 : _GEN_6211; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8207 = 5'hb == rob_head ? 32'h4033 : _GEN_6214; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8208 = 5'hc == rob_head ? 32'h4033 : _GEN_6217; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8209 = 5'hd == rob_head ? 32'h4033 : _GEN_6220; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8210 = 5'he == rob_head ? 32'h4033 : _GEN_6223; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8211 = 5'hf == rob_head ? 32'h4033 : _GEN_6226; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8212 = 5'h10 == rob_head ? 32'h4033 : _GEN_6229; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8213 = 5'h11 == rob_head ? 32'h4033 : _GEN_6232; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8214 = 5'h12 == rob_head ? 32'h4033 : _GEN_6235; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8215 = 5'h13 == rob_head ? 32'h4033 : _GEN_6238; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8216 = 5'h14 == rob_head ? 32'h4033 : _GEN_6241; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8217 = 5'h15 == rob_head ? 32'h4033 : _GEN_6244; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8218 = 5'h16 == rob_head ? 32'h4033 : _GEN_6247; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8219 = 5'h17 == rob_head ? 32'h4033 : _GEN_6250; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_8220 = T_47546 ? _GEN_8196 : _GEN_6181; // @[rob.scala 514:7]
  wire [31:0] _GEN_8221 = T_47546 ? _GEN_8197 : _GEN_6184; // @[rob.scala 514:7]
  wire [31:0] _GEN_8222 = T_47546 ? _GEN_8198 : _GEN_6187; // @[rob.scala 514:7]
  wire [31:0] _GEN_8223 = T_47546 ? _GEN_8199 : _GEN_6190; // @[rob.scala 514:7]
  wire [31:0] _GEN_8224 = T_47546 ? _GEN_8200 : _GEN_6193; // @[rob.scala 514:7]
  wire [31:0] _GEN_8225 = T_47546 ? _GEN_8201 : _GEN_6196; // @[rob.scala 514:7]
  wire [31:0] _GEN_8226 = T_47546 ? _GEN_8202 : _GEN_6199; // @[rob.scala 514:7]
  wire [31:0] _GEN_8227 = T_47546 ? _GEN_8203 : _GEN_6202; // @[rob.scala 514:7]
  wire [31:0] _GEN_8228 = T_47546 ? _GEN_8204 : _GEN_6205; // @[rob.scala 514:7]
  wire [31:0] _GEN_8229 = T_47546 ? _GEN_8205 : _GEN_6208; // @[rob.scala 514:7]
  wire [31:0] _GEN_8230 = T_47546 ? _GEN_8206 : _GEN_6211; // @[rob.scala 514:7]
  wire [31:0] _GEN_8231 = T_47546 ? _GEN_8207 : _GEN_6214; // @[rob.scala 514:7]
  wire [31:0] _GEN_8232 = T_47546 ? _GEN_8208 : _GEN_6217; // @[rob.scala 514:7]
  wire [31:0] _GEN_8233 = T_47546 ? _GEN_8209 : _GEN_6220; // @[rob.scala 514:7]
  wire [31:0] _GEN_8234 = T_47546 ? _GEN_8210 : _GEN_6223; // @[rob.scala 514:7]
  wire [31:0] _GEN_8235 = T_47546 ? _GEN_8211 : _GEN_6226; // @[rob.scala 514:7]
  wire [31:0] _GEN_8236 = T_47546 ? _GEN_8212 : _GEN_6229; // @[rob.scala 514:7]
  wire [31:0] _GEN_8237 = T_47546 ? _GEN_8213 : _GEN_6232; // @[rob.scala 514:7]
  wire [31:0] _GEN_8238 = T_47546 ? _GEN_8214 : _GEN_6235; // @[rob.scala 514:7]
  wire [31:0] _GEN_8239 = T_47546 ? _GEN_8215 : _GEN_6238; // @[rob.scala 514:7]
  wire [31:0] _GEN_8240 = T_47546 ? _GEN_8216 : _GEN_6241; // @[rob.scala 514:7]
  wire [31:0] _GEN_8241 = T_47546 ? _GEN_8217 : _GEN_6244; // @[rob.scala 514:7]
  wire [31:0] _GEN_8242 = T_47546 ? _GEN_8218 : _GEN_6247; // @[rob.scala 514:7]
  wire [31:0] _GEN_8243 = T_47546 ? _GEN_8219 : _GEN_6250; // @[rob.scala 514:7]
  wire  T_32081 = ~T_47546; // @[rob.scala 514:7]
  wire  T_32082 = T_32081 & T_29097; // @[rob.scala 518:7]
  wire  T_32171 = io_debug_wb_valids_0 & T_28592; // @[rob.scala 529:38]
  wire [63:0] _GEN_8292 = 6'h0 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3806; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8293 = 6'h1 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3807; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8294 = 6'h2 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3808; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8295 = 6'h3 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3809; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8296 = 6'h4 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3810; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8297 = 6'h5 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3811; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8298 = 6'h6 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3812; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8299 = 6'h7 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3813; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8300 = 6'h8 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3814; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8301 = 6'h9 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3815; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8302 = 6'ha == T_28589 ? io_debug_wb_wdata_0 : _GEN_3816; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8303 = 6'hb == T_28589 ? io_debug_wb_wdata_0 : _GEN_3817; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8304 = 6'hc == T_28589 ? io_debug_wb_wdata_0 : _GEN_3818; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8305 = 6'hd == T_28589 ? io_debug_wb_wdata_0 : _GEN_3819; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8306 = 6'he == T_28589 ? io_debug_wb_wdata_0 : _GEN_3820; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8307 = 6'hf == T_28589 ? io_debug_wb_wdata_0 : _GEN_3821; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8308 = 6'h10 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3822; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8309 = 6'h11 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3823; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8310 = 6'h12 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3824; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8311 = 6'h13 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3825; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8312 = 6'h14 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3826; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8313 = 6'h15 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3827; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8314 = 6'h16 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3828; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8315 = 6'h17 == T_28589 ? io_debug_wb_wdata_0 : _GEN_3829; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_8316 = T_32171 ? _GEN_8292 : _GEN_3806; // @[rob.scala 530:10]
  wire [63:0] _GEN_8317 = T_32171 ? _GEN_8293 : _GEN_3807; // @[rob.scala 530:10]
  wire [63:0] _GEN_8318 = T_32171 ? _GEN_8294 : _GEN_3808; // @[rob.scala 530:10]
  wire [63:0] _GEN_8319 = T_32171 ? _GEN_8295 : _GEN_3809; // @[rob.scala 530:10]
  wire [63:0] _GEN_8320 = T_32171 ? _GEN_8296 : _GEN_3810; // @[rob.scala 530:10]
  wire [63:0] _GEN_8321 = T_32171 ? _GEN_8297 : _GEN_3811; // @[rob.scala 530:10]
  wire [63:0] _GEN_8322 = T_32171 ? _GEN_8298 : _GEN_3812; // @[rob.scala 530:10]
  wire [63:0] _GEN_8323 = T_32171 ? _GEN_8299 : _GEN_3813; // @[rob.scala 530:10]
  wire [63:0] _GEN_8324 = T_32171 ? _GEN_8300 : _GEN_3814; // @[rob.scala 530:10]
  wire [63:0] _GEN_8325 = T_32171 ? _GEN_8301 : _GEN_3815; // @[rob.scala 530:10]
  wire [63:0] _GEN_8326 = T_32171 ? _GEN_8302 : _GEN_3816; // @[rob.scala 530:10]
  wire [63:0] _GEN_8327 = T_32171 ? _GEN_8303 : _GEN_3817; // @[rob.scala 530:10]
  wire [63:0] _GEN_8328 = T_32171 ? _GEN_8304 : _GEN_3818; // @[rob.scala 530:10]
  wire [63:0] _GEN_8329 = T_32171 ? _GEN_8305 : _GEN_3819; // @[rob.scala 530:10]
  wire [63:0] _GEN_8330 = T_32171 ? _GEN_8306 : _GEN_3820; // @[rob.scala 530:10]
  wire [63:0] _GEN_8331 = T_32171 ? _GEN_8307 : _GEN_3821; // @[rob.scala 530:10]
  wire [63:0] _GEN_8332 = T_32171 ? _GEN_8308 : _GEN_3822; // @[rob.scala 530:10]
  wire [63:0] _GEN_8333 = T_32171 ? _GEN_8309 : _GEN_3823; // @[rob.scala 530:10]
  wire [63:0] _GEN_8334 = T_32171 ? _GEN_8310 : _GEN_3824; // @[rob.scala 530:10]
  wire [63:0] _GEN_8335 = T_32171 ? _GEN_8311 : _GEN_3825; // @[rob.scala 530:10]
  wire [63:0] _GEN_8336 = T_32171 ? _GEN_8312 : _GEN_3826; // @[rob.scala 530:10]
  wire [63:0] _GEN_8337 = T_32171 ? _GEN_8313 : _GEN_3827; // @[rob.scala 530:10]
  wire [63:0] _GEN_8338 = T_32171 ? _GEN_8314 : _GEN_3828; // @[rob.scala 530:10]
  wire [63:0] _GEN_8339 = T_32171 ? _GEN_8315 : _GEN_3829; // @[rob.scala 530:10]
  wire  _GEN_8341 = 6'h1 == T_28589 ? T_23706_1 : T_23706_0; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8342 = 6'h2 == T_28589 ? T_23706_2 : _GEN_8341; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8343 = 6'h3 == T_28589 ? T_23706_3 : _GEN_8342; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8344 = 6'h4 == T_28589 ? T_23706_4 : _GEN_8343; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8345 = 6'h5 == T_28589 ? T_23706_5 : _GEN_8344; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8346 = 6'h6 == T_28589 ? T_23706_6 : _GEN_8345; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8347 = 6'h7 == T_28589 ? T_23706_7 : _GEN_8346; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8348 = 6'h8 == T_28589 ? T_23706_8 : _GEN_8347; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8349 = 6'h9 == T_28589 ? T_23706_9 : _GEN_8348; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8350 = 6'ha == T_28589 ? T_23706_10 : _GEN_8349; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8351 = 6'hb == T_28589 ? T_23706_11 : _GEN_8350; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8352 = 6'hc == T_28589 ? T_23706_12 : _GEN_8351; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8353 = 6'hd == T_28589 ? T_23706_13 : _GEN_8352; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8354 = 6'he == T_28589 ? T_23706_14 : _GEN_8353; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8355 = 6'hf == T_28589 ? T_23706_15 : _GEN_8354; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8356 = 6'h10 == T_28589 ? T_23706_16 : _GEN_8355; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8357 = 6'h11 == T_28589 ? T_23706_17 : _GEN_8356; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8358 = 6'h12 == T_28589 ? T_23706_18 : _GEN_8357; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8359 = 6'h13 == T_28589 ? T_23706_19 : _GEN_8358; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8360 = 6'h14 == T_28589 ? T_23706_20 : _GEN_8359; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8361 = 6'h15 == T_28589 ? T_23706_21 : _GEN_8360; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8362 = 6'h16 == T_28589 ? T_23706_22 : _GEN_8361; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_8363 = 6'h17 == T_28589 ? T_23706_23 : _GEN_8362; // @[rob.scala 536:22 rob.scala 536:22]
  wire  T_32353 = ~_GEN_8363; // @[rob.scala 536:22]
  wire  T_32354 = T_28593 & T_32353; // @[rob.scala 535:75]
  wire  T_32356 = ~T_32354; // @[rob.scala 535:18]
  wire  T_32357 = T_32356 | reset; // @[rob.scala 535:17]
  wire  T_32359 = ~T_32357; // @[rob.scala 535:17]
  wire [6:0] _GEN_8485 = 6'h1 == T_28589 ? T_26182_1_pdst : T_26182_0_pdst; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8509 = 6'h1 == T_28589 ? T_26182_1_ldst_val : T_26182_0_ldst_val; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_8563 = 6'h2 == T_28589 ? T_26182_2_pdst : _GEN_8485; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8587 = 6'h2 == T_28589 ? T_26182_2_ldst_val : _GEN_8509; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_8641 = 6'h3 == T_28589 ? T_26182_3_pdst : _GEN_8563; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8665 = 6'h3 == T_28589 ? T_26182_3_ldst_val : _GEN_8587; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_8719 = 6'h4 == T_28589 ? T_26182_4_pdst : _GEN_8641; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8743 = 6'h4 == T_28589 ? T_26182_4_ldst_val : _GEN_8665; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_8797 = 6'h5 == T_28589 ? T_26182_5_pdst : _GEN_8719; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8821 = 6'h5 == T_28589 ? T_26182_5_ldst_val : _GEN_8743; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_8875 = 6'h6 == T_28589 ? T_26182_6_pdst : _GEN_8797; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8899 = 6'h6 == T_28589 ? T_26182_6_ldst_val : _GEN_8821; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_8953 = 6'h7 == T_28589 ? T_26182_7_pdst : _GEN_8875; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_8977 = 6'h7 == T_28589 ? T_26182_7_ldst_val : _GEN_8899; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9031 = 6'h8 == T_28589 ? T_26182_8_pdst : _GEN_8953; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9055 = 6'h8 == T_28589 ? T_26182_8_ldst_val : _GEN_8977; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9109 = 6'h9 == T_28589 ? T_26182_9_pdst : _GEN_9031; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9133 = 6'h9 == T_28589 ? T_26182_9_ldst_val : _GEN_9055; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9187 = 6'ha == T_28589 ? T_26182_10_pdst : _GEN_9109; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9211 = 6'ha == T_28589 ? T_26182_10_ldst_val : _GEN_9133; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9265 = 6'hb == T_28589 ? T_26182_11_pdst : _GEN_9187; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9289 = 6'hb == T_28589 ? T_26182_11_ldst_val : _GEN_9211; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9343 = 6'hc == T_28589 ? T_26182_12_pdst : _GEN_9265; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9367 = 6'hc == T_28589 ? T_26182_12_ldst_val : _GEN_9289; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9421 = 6'hd == T_28589 ? T_26182_13_pdst : _GEN_9343; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9445 = 6'hd == T_28589 ? T_26182_13_ldst_val : _GEN_9367; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9499 = 6'he == T_28589 ? T_26182_14_pdst : _GEN_9421; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9523 = 6'he == T_28589 ? T_26182_14_ldst_val : _GEN_9445; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9577 = 6'hf == T_28589 ? T_26182_15_pdst : _GEN_9499; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9601 = 6'hf == T_28589 ? T_26182_15_ldst_val : _GEN_9523; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9655 = 6'h10 == T_28589 ? T_26182_16_pdst : _GEN_9577; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9679 = 6'h10 == T_28589 ? T_26182_16_ldst_val : _GEN_9601; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9733 = 6'h11 == T_28589 ? T_26182_17_pdst : _GEN_9655; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9757 = 6'h11 == T_28589 ? T_26182_17_ldst_val : _GEN_9679; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9811 = 6'h12 == T_28589 ? T_26182_18_pdst : _GEN_9733; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9835 = 6'h12 == T_28589 ? T_26182_18_ldst_val : _GEN_9757; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9889 = 6'h13 == T_28589 ? T_26182_19_pdst : _GEN_9811; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9913 = 6'h13 == T_28589 ? T_26182_19_ldst_val : _GEN_9835; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_9967 = 6'h14 == T_28589 ? T_26182_20_pdst : _GEN_9889; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_9991 = 6'h14 == T_28589 ? T_26182_20_ldst_val : _GEN_9913; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10045 = 6'h15 == T_28589 ? T_26182_21_pdst : _GEN_9967; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10069 = 6'h15 == T_28589 ? T_26182_21_ldst_val : _GEN_9991; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10123 = 6'h16 == T_28589 ? T_26182_22_pdst : _GEN_10045; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10147 = 6'h16 == T_28589 ? T_26182_22_ldst_val : _GEN_10069; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10201 = 6'h17 == T_28589 ? T_26182_23_pdst : _GEN_10123; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10225 = 6'h17 == T_28589 ? T_26182_23_ldst_val : _GEN_10147; // @[rob.scala 538:75 rob.scala 538:75]
  wire  T_32364 = T_28593 & _GEN_10225; // @[rob.scala 538:75]
  wire  T_32365 = _GEN_10201 != io_wb_resps_0_bits_uop_pdst; // @[rob.scala 539:54]
  wire  T_32366 = T_32364 & T_32365; // @[rob.scala 539:37]
  wire  T_32368 = ~T_32366; // @[rob.scala 538:18]
  wire  T_32369 = T_32368 | reset; // @[rob.scala 538:17]
  wire  T_32371 = ~T_32369; // @[rob.scala 538:17]
  wire  T_32375 = io_debug_wb_valids_1 & T_28600; // @[rob.scala 529:38]
  wire [63:0] _GEN_10236 = 6'h0 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8316; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10237 = 6'h1 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8317; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10238 = 6'h2 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8318; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10239 = 6'h3 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8319; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10240 = 6'h4 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8320; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10241 = 6'h5 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8321; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10242 = 6'h6 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8322; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10243 = 6'h7 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8323; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10244 = 6'h8 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8324; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10245 = 6'h9 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8325; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10246 = 6'ha == T_28597 ? io_debug_wb_wdata_1 : _GEN_8326; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10247 = 6'hb == T_28597 ? io_debug_wb_wdata_1 : _GEN_8327; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10248 = 6'hc == T_28597 ? io_debug_wb_wdata_1 : _GEN_8328; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10249 = 6'hd == T_28597 ? io_debug_wb_wdata_1 : _GEN_8329; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10250 = 6'he == T_28597 ? io_debug_wb_wdata_1 : _GEN_8330; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10251 = 6'hf == T_28597 ? io_debug_wb_wdata_1 : _GEN_8331; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10252 = 6'h10 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8332; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10253 = 6'h11 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8333; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10254 = 6'h12 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8334; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10255 = 6'h13 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8335; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10256 = 6'h14 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8336; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10257 = 6'h15 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8337; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10258 = 6'h16 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8338; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10259 = 6'h17 == T_28597 ? io_debug_wb_wdata_1 : _GEN_8339; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_10260 = T_32375 ? _GEN_10236 : _GEN_8316; // @[rob.scala 530:10]
  wire [63:0] _GEN_10261 = T_32375 ? _GEN_10237 : _GEN_8317; // @[rob.scala 530:10]
  wire [63:0] _GEN_10262 = T_32375 ? _GEN_10238 : _GEN_8318; // @[rob.scala 530:10]
  wire [63:0] _GEN_10263 = T_32375 ? _GEN_10239 : _GEN_8319; // @[rob.scala 530:10]
  wire [63:0] _GEN_10264 = T_32375 ? _GEN_10240 : _GEN_8320; // @[rob.scala 530:10]
  wire [63:0] _GEN_10265 = T_32375 ? _GEN_10241 : _GEN_8321; // @[rob.scala 530:10]
  wire [63:0] _GEN_10266 = T_32375 ? _GEN_10242 : _GEN_8322; // @[rob.scala 530:10]
  wire [63:0] _GEN_10267 = T_32375 ? _GEN_10243 : _GEN_8323; // @[rob.scala 530:10]
  wire [63:0] _GEN_10268 = T_32375 ? _GEN_10244 : _GEN_8324; // @[rob.scala 530:10]
  wire [63:0] _GEN_10269 = T_32375 ? _GEN_10245 : _GEN_8325; // @[rob.scala 530:10]
  wire [63:0] _GEN_10270 = T_32375 ? _GEN_10246 : _GEN_8326; // @[rob.scala 530:10]
  wire [63:0] _GEN_10271 = T_32375 ? _GEN_10247 : _GEN_8327; // @[rob.scala 530:10]
  wire [63:0] _GEN_10272 = T_32375 ? _GEN_10248 : _GEN_8328; // @[rob.scala 530:10]
  wire [63:0] _GEN_10273 = T_32375 ? _GEN_10249 : _GEN_8329; // @[rob.scala 530:10]
  wire [63:0] _GEN_10274 = T_32375 ? _GEN_10250 : _GEN_8330; // @[rob.scala 530:10]
  wire [63:0] _GEN_10275 = T_32375 ? _GEN_10251 : _GEN_8331; // @[rob.scala 530:10]
  wire [63:0] _GEN_10276 = T_32375 ? _GEN_10252 : _GEN_8332; // @[rob.scala 530:10]
  wire [63:0] _GEN_10277 = T_32375 ? _GEN_10253 : _GEN_8333; // @[rob.scala 530:10]
  wire [63:0] _GEN_10278 = T_32375 ? _GEN_10254 : _GEN_8334; // @[rob.scala 530:10]
  wire [63:0] _GEN_10279 = T_32375 ? _GEN_10255 : _GEN_8335; // @[rob.scala 530:10]
  wire [63:0] _GEN_10280 = T_32375 ? _GEN_10256 : _GEN_8336; // @[rob.scala 530:10]
  wire [63:0] _GEN_10281 = T_32375 ? _GEN_10257 : _GEN_8337; // @[rob.scala 530:10]
  wire [63:0] _GEN_10282 = T_32375 ? _GEN_10258 : _GEN_8338; // @[rob.scala 530:10]
  wire [63:0] _GEN_10283 = T_32375 ? _GEN_10259 : _GEN_8339; // @[rob.scala 530:10]
  wire  _GEN_10285 = 6'h1 == T_28597 ? T_23706_1 : T_23706_0; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10286 = 6'h2 == T_28597 ? T_23706_2 : _GEN_10285; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10287 = 6'h3 == T_28597 ? T_23706_3 : _GEN_10286; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10288 = 6'h4 == T_28597 ? T_23706_4 : _GEN_10287; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10289 = 6'h5 == T_28597 ? T_23706_5 : _GEN_10288; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10290 = 6'h6 == T_28597 ? T_23706_6 : _GEN_10289; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10291 = 6'h7 == T_28597 ? T_23706_7 : _GEN_10290; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10292 = 6'h8 == T_28597 ? T_23706_8 : _GEN_10291; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10293 = 6'h9 == T_28597 ? T_23706_9 : _GEN_10292; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10294 = 6'ha == T_28597 ? T_23706_10 : _GEN_10293; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10295 = 6'hb == T_28597 ? T_23706_11 : _GEN_10294; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10296 = 6'hc == T_28597 ? T_23706_12 : _GEN_10295; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10297 = 6'hd == T_28597 ? T_23706_13 : _GEN_10296; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10298 = 6'he == T_28597 ? T_23706_14 : _GEN_10297; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10299 = 6'hf == T_28597 ? T_23706_15 : _GEN_10298; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10300 = 6'h10 == T_28597 ? T_23706_16 : _GEN_10299; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10301 = 6'h11 == T_28597 ? T_23706_17 : _GEN_10300; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10302 = 6'h12 == T_28597 ? T_23706_18 : _GEN_10301; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10303 = 6'h13 == T_28597 ? T_23706_19 : _GEN_10302; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10304 = 6'h14 == T_28597 ? T_23706_20 : _GEN_10303; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10305 = 6'h15 == T_28597 ? T_23706_21 : _GEN_10304; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10306 = 6'h16 == T_28597 ? T_23706_22 : _GEN_10305; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_10307 = 6'h17 == T_28597 ? T_23706_23 : _GEN_10306; // @[rob.scala 536:22 rob.scala 536:22]
  wire  T_32557 = ~_GEN_10307; // @[rob.scala 536:22]
  wire  T_32558 = T_28601 & T_32557; // @[rob.scala 535:75]
  wire  T_32560 = ~T_32558; // @[rob.scala 535:18]
  wire  T_32561 = T_32560 | reset; // @[rob.scala 535:17]
  wire  T_32563 = ~T_32561; // @[rob.scala 535:17]
  wire [6:0] _GEN_10429 = 6'h1 == T_28597 ? T_26182_1_pdst : T_26182_0_pdst; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10453 = 6'h1 == T_28597 ? T_26182_1_ldst_val : T_26182_0_ldst_val; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10507 = 6'h2 == T_28597 ? T_26182_2_pdst : _GEN_10429; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10531 = 6'h2 == T_28597 ? T_26182_2_ldst_val : _GEN_10453; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10585 = 6'h3 == T_28597 ? T_26182_3_pdst : _GEN_10507; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10609 = 6'h3 == T_28597 ? T_26182_3_ldst_val : _GEN_10531; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10663 = 6'h4 == T_28597 ? T_26182_4_pdst : _GEN_10585; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10687 = 6'h4 == T_28597 ? T_26182_4_ldst_val : _GEN_10609; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10741 = 6'h5 == T_28597 ? T_26182_5_pdst : _GEN_10663; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10765 = 6'h5 == T_28597 ? T_26182_5_ldst_val : _GEN_10687; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10819 = 6'h6 == T_28597 ? T_26182_6_pdst : _GEN_10741; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10843 = 6'h6 == T_28597 ? T_26182_6_ldst_val : _GEN_10765; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10897 = 6'h7 == T_28597 ? T_26182_7_pdst : _GEN_10819; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10921 = 6'h7 == T_28597 ? T_26182_7_ldst_val : _GEN_10843; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_10975 = 6'h8 == T_28597 ? T_26182_8_pdst : _GEN_10897; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_10999 = 6'h8 == T_28597 ? T_26182_8_ldst_val : _GEN_10921; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11053 = 6'h9 == T_28597 ? T_26182_9_pdst : _GEN_10975; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11077 = 6'h9 == T_28597 ? T_26182_9_ldst_val : _GEN_10999; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11131 = 6'ha == T_28597 ? T_26182_10_pdst : _GEN_11053; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11155 = 6'ha == T_28597 ? T_26182_10_ldst_val : _GEN_11077; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11209 = 6'hb == T_28597 ? T_26182_11_pdst : _GEN_11131; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11233 = 6'hb == T_28597 ? T_26182_11_ldst_val : _GEN_11155; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11287 = 6'hc == T_28597 ? T_26182_12_pdst : _GEN_11209; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11311 = 6'hc == T_28597 ? T_26182_12_ldst_val : _GEN_11233; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11365 = 6'hd == T_28597 ? T_26182_13_pdst : _GEN_11287; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11389 = 6'hd == T_28597 ? T_26182_13_ldst_val : _GEN_11311; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11443 = 6'he == T_28597 ? T_26182_14_pdst : _GEN_11365; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11467 = 6'he == T_28597 ? T_26182_14_ldst_val : _GEN_11389; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11521 = 6'hf == T_28597 ? T_26182_15_pdst : _GEN_11443; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11545 = 6'hf == T_28597 ? T_26182_15_ldst_val : _GEN_11467; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11599 = 6'h10 == T_28597 ? T_26182_16_pdst : _GEN_11521; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11623 = 6'h10 == T_28597 ? T_26182_16_ldst_val : _GEN_11545; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11677 = 6'h11 == T_28597 ? T_26182_17_pdst : _GEN_11599; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11701 = 6'h11 == T_28597 ? T_26182_17_ldst_val : _GEN_11623; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11755 = 6'h12 == T_28597 ? T_26182_18_pdst : _GEN_11677; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11779 = 6'h12 == T_28597 ? T_26182_18_ldst_val : _GEN_11701; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11833 = 6'h13 == T_28597 ? T_26182_19_pdst : _GEN_11755; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11857 = 6'h13 == T_28597 ? T_26182_19_ldst_val : _GEN_11779; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11911 = 6'h14 == T_28597 ? T_26182_20_pdst : _GEN_11833; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_11935 = 6'h14 == T_28597 ? T_26182_20_ldst_val : _GEN_11857; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_11989 = 6'h15 == T_28597 ? T_26182_21_pdst : _GEN_11911; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12013 = 6'h15 == T_28597 ? T_26182_21_ldst_val : _GEN_11935; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12067 = 6'h16 == T_28597 ? T_26182_22_pdst : _GEN_11989; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12091 = 6'h16 == T_28597 ? T_26182_22_ldst_val : _GEN_12013; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12145 = 6'h17 == T_28597 ? T_26182_23_pdst : _GEN_12067; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12169 = 6'h17 == T_28597 ? T_26182_23_ldst_val : _GEN_12091; // @[rob.scala 538:75 rob.scala 538:75]
  wire  T_32568 = T_28601 & _GEN_12169; // @[rob.scala 538:75]
  wire  T_32569 = _GEN_12145 != io_wb_resps_1_bits_uop_pdst; // @[rob.scala 539:54]
  wire  T_32570 = T_32568 & T_32569; // @[rob.scala 539:37]
  wire  T_32572 = ~T_32570; // @[rob.scala 538:18]
  wire  T_32573 = T_32572 | reset; // @[rob.scala 538:17]
  wire  T_32575 = ~T_32573; // @[rob.scala 538:17]
  wire  T_32579 = io_debug_wb_valids_2 & T_28608; // @[rob.scala 529:38]
  wire  _GEN_12229 = 6'h1 == T_28605 ? T_23706_1 : T_23706_0; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12230 = 6'h2 == T_28605 ? T_23706_2 : _GEN_12229; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12231 = 6'h3 == T_28605 ? T_23706_3 : _GEN_12230; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12232 = 6'h4 == T_28605 ? T_23706_4 : _GEN_12231; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12233 = 6'h5 == T_28605 ? T_23706_5 : _GEN_12232; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12234 = 6'h6 == T_28605 ? T_23706_6 : _GEN_12233; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12235 = 6'h7 == T_28605 ? T_23706_7 : _GEN_12234; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12236 = 6'h8 == T_28605 ? T_23706_8 : _GEN_12235; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12237 = 6'h9 == T_28605 ? T_23706_9 : _GEN_12236; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12238 = 6'ha == T_28605 ? T_23706_10 : _GEN_12237; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12239 = 6'hb == T_28605 ? T_23706_11 : _GEN_12238; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12240 = 6'hc == T_28605 ? T_23706_12 : _GEN_12239; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12241 = 6'hd == T_28605 ? T_23706_13 : _GEN_12240; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12242 = 6'he == T_28605 ? T_23706_14 : _GEN_12241; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12243 = 6'hf == T_28605 ? T_23706_15 : _GEN_12242; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12244 = 6'h10 == T_28605 ? T_23706_16 : _GEN_12243; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12245 = 6'h11 == T_28605 ? T_23706_17 : _GEN_12244; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12246 = 6'h12 == T_28605 ? T_23706_18 : _GEN_12245; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12247 = 6'h13 == T_28605 ? T_23706_19 : _GEN_12246; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12248 = 6'h14 == T_28605 ? T_23706_20 : _GEN_12247; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12249 = 6'h15 == T_28605 ? T_23706_21 : _GEN_12248; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12250 = 6'h16 == T_28605 ? T_23706_22 : _GEN_12249; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_12251 = 6'h17 == T_28605 ? T_23706_23 : _GEN_12250; // @[rob.scala 536:22 rob.scala 536:22]
  wire  T_32761 = ~_GEN_12251; // @[rob.scala 536:22]
  wire  T_32762 = T_28609 & T_32761; // @[rob.scala 535:75]
  wire  T_32764 = ~T_32762; // @[rob.scala 535:18]
  wire  T_32765 = T_32764 | reset; // @[rob.scala 535:17]
  wire  T_32767 = ~T_32765; // @[rob.scala 535:17]
  wire [6:0] _GEN_12373 = 6'h1 == T_28605 ? T_26182_1_pdst : T_26182_0_pdst; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12397 = 6'h1 == T_28605 ? T_26182_1_ldst_val : T_26182_0_ldst_val; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12451 = 6'h2 == T_28605 ? T_26182_2_pdst : _GEN_12373; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12475 = 6'h2 == T_28605 ? T_26182_2_ldst_val : _GEN_12397; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12529 = 6'h3 == T_28605 ? T_26182_3_pdst : _GEN_12451; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12553 = 6'h3 == T_28605 ? T_26182_3_ldst_val : _GEN_12475; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12607 = 6'h4 == T_28605 ? T_26182_4_pdst : _GEN_12529; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12631 = 6'h4 == T_28605 ? T_26182_4_ldst_val : _GEN_12553; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12685 = 6'h5 == T_28605 ? T_26182_5_pdst : _GEN_12607; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12709 = 6'h5 == T_28605 ? T_26182_5_ldst_val : _GEN_12631; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12763 = 6'h6 == T_28605 ? T_26182_6_pdst : _GEN_12685; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12787 = 6'h6 == T_28605 ? T_26182_6_ldst_val : _GEN_12709; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12841 = 6'h7 == T_28605 ? T_26182_7_pdst : _GEN_12763; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12865 = 6'h7 == T_28605 ? T_26182_7_ldst_val : _GEN_12787; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12919 = 6'h8 == T_28605 ? T_26182_8_pdst : _GEN_12841; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_12943 = 6'h8 == T_28605 ? T_26182_8_ldst_val : _GEN_12865; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_12997 = 6'h9 == T_28605 ? T_26182_9_pdst : _GEN_12919; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13021 = 6'h9 == T_28605 ? T_26182_9_ldst_val : _GEN_12943; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13075 = 6'ha == T_28605 ? T_26182_10_pdst : _GEN_12997; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13099 = 6'ha == T_28605 ? T_26182_10_ldst_val : _GEN_13021; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13153 = 6'hb == T_28605 ? T_26182_11_pdst : _GEN_13075; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13177 = 6'hb == T_28605 ? T_26182_11_ldst_val : _GEN_13099; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13231 = 6'hc == T_28605 ? T_26182_12_pdst : _GEN_13153; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13255 = 6'hc == T_28605 ? T_26182_12_ldst_val : _GEN_13177; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13309 = 6'hd == T_28605 ? T_26182_13_pdst : _GEN_13231; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13333 = 6'hd == T_28605 ? T_26182_13_ldst_val : _GEN_13255; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13387 = 6'he == T_28605 ? T_26182_14_pdst : _GEN_13309; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13411 = 6'he == T_28605 ? T_26182_14_ldst_val : _GEN_13333; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13465 = 6'hf == T_28605 ? T_26182_15_pdst : _GEN_13387; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13489 = 6'hf == T_28605 ? T_26182_15_ldst_val : _GEN_13411; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13543 = 6'h10 == T_28605 ? T_26182_16_pdst : _GEN_13465; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13567 = 6'h10 == T_28605 ? T_26182_16_ldst_val : _GEN_13489; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13621 = 6'h11 == T_28605 ? T_26182_17_pdst : _GEN_13543; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13645 = 6'h11 == T_28605 ? T_26182_17_ldst_val : _GEN_13567; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13699 = 6'h12 == T_28605 ? T_26182_18_pdst : _GEN_13621; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13723 = 6'h12 == T_28605 ? T_26182_18_ldst_val : _GEN_13645; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13777 = 6'h13 == T_28605 ? T_26182_19_pdst : _GEN_13699; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13801 = 6'h13 == T_28605 ? T_26182_19_ldst_val : _GEN_13723; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13855 = 6'h14 == T_28605 ? T_26182_20_pdst : _GEN_13777; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13879 = 6'h14 == T_28605 ? T_26182_20_ldst_val : _GEN_13801; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_13933 = 6'h15 == T_28605 ? T_26182_21_pdst : _GEN_13855; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_13957 = 6'h15 == T_28605 ? T_26182_21_ldst_val : _GEN_13879; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_14011 = 6'h16 == T_28605 ? T_26182_22_pdst : _GEN_13933; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_14035 = 6'h16 == T_28605 ? T_26182_22_ldst_val : _GEN_13957; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_14089 = 6'h17 == T_28605 ? T_26182_23_pdst : _GEN_14011; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_14113 = 6'h17 == T_28605 ? T_26182_23_ldst_val : _GEN_14035; // @[rob.scala 538:75 rob.scala 538:75]
  wire  T_32772 = T_28609 & _GEN_14113; // @[rob.scala 538:75]
  wire  T_32773 = _GEN_14089 != io_wb_resps_2_bits_uop_pdst; // @[rob.scala 539:54]
  wire  T_32774 = T_32772 & T_32773; // @[rob.scala 539:37]
  wire  T_32776 = ~T_32774; // @[rob.scala 538:18]
  wire  T_32777 = T_32776 | reset; // @[rob.scala 538:17]
  wire  T_32779 = ~T_32777; // @[rob.scala 538:17]
  wire [39:0] T_32960 = {T_23555_T_32958_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_32955 = {{24'd0}, T_32960}; // @[rob.scala 899:26]
  wire [39:0] T_32967 = T_32955[39:0]; // @[rob.scala 906:20]
  wire  T_32968 = T_32967[39]; // @[util.scala 114:43]
  wire [23:0] T_32972 = T_32968 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_32973 = {T_32972,T_32967}; // @[Cat.scala 20:58]
  wire [64:0] T_32975 = {{1'd0}, T_32973}; // @[rob.scala 554:94]
  wire [63:0] T_32976 = T_32975[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33080 = {T_23558_T_33078_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_33069 = {{24'd0}, T_33080}; // @[rob.scala 899:26]
  wire [39:0] T_33081 = T_33069[39:0]; // @[rob.scala 906:20]
  wire  T_33082 = T_33081[39]; // @[util.scala 114:43]
  wire [23:0] T_33086 = T_33082 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33087 = {T_33086,T_33081}; // @[Cat.scala 20:58]
  wire [64:0] T_33089 = {{1'd0}, T_33087}; // @[rob.scala 554:94]
  wire [63:0] T_33090 = T_33089[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33188 = {T_23555_T_33186_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_33183 = {{24'd0}, T_33188}; // @[rob.scala 899:26]
  wire [39:0] T_33195 = T_33183[39:0]; // @[rob.scala 906:20]
  wire  T_33196 = T_33195[39]; // @[util.scala 114:43]
  wire [23:0] T_33200 = T_33196 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33201 = {T_33200,T_33195}; // @[Cat.scala 20:58]
  wire [64:0] T_33203 = {{1'd0}, T_33201}; // @[rob.scala 554:94]
  wire [63:0] T_33204 = T_33203[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33308 = {T_23558_T_33306_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_33297 = {{24'd0}, T_33308}; // @[rob.scala 899:26]
  wire [39:0] T_33309 = T_33297[39:0]; // @[rob.scala 906:20]
  wire  T_33310 = T_33309[39]; // @[util.scala 114:43]
  wire [23:0] T_33314 = T_33310 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33315 = {T_33314,T_33309}; // @[Cat.scala 20:58]
  wire [64:0] T_33317 = {{1'd0}, T_33315}; // @[rob.scala 554:94]
  wire [63:0] T_33318 = T_33317[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33416 = {T_23555_T_33414_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_33411 = {{24'd0}, T_33416}; // @[rob.scala 899:26]
  wire [39:0] T_33423 = T_33411[39:0]; // @[rob.scala 906:20]
  wire  T_33424 = T_33423[39]; // @[util.scala 114:43]
  wire [23:0] T_33428 = T_33424 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33429 = {T_33428,T_33423}; // @[Cat.scala 20:58]
  wire [64:0] T_33431 = {{1'd0}, T_33429}; // @[rob.scala 554:94]
  wire [63:0] T_33432 = T_33431[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33536 = {T_23558_T_33534_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_33525 = {{24'd0}, T_33536}; // @[rob.scala 899:26]
  wire [39:0] T_33537 = T_33525[39:0]; // @[rob.scala 906:20]
  wire  T_33538 = T_33537[39]; // @[util.scala 114:43]
  wire [23:0] T_33542 = T_33538 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33543 = {T_33542,T_33537}; // @[Cat.scala 20:58]
  wire [64:0] T_33545 = {{1'd0}, T_33543}; // @[rob.scala 554:94]
  wire [63:0] T_33546 = T_33545[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33644 = {T_23555_T_33642_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_33639 = {{24'd0}, T_33644}; // @[rob.scala 899:26]
  wire [39:0] T_33651 = T_33639[39:0]; // @[rob.scala 906:20]
  wire  T_33652 = T_33651[39]; // @[util.scala 114:43]
  wire [23:0] T_33656 = T_33652 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33657 = {T_33656,T_33651}; // @[Cat.scala 20:58]
  wire [64:0] T_33659 = {{1'd0}, T_33657}; // @[rob.scala 554:94]
  wire [63:0] T_33660 = T_33659[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33764 = {T_23558_T_33762_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_33753 = {{24'd0}, T_33764}; // @[rob.scala 899:26]
  wire [39:0] T_33765 = T_33753[39:0]; // @[rob.scala 906:20]
  wire  T_33766 = T_33765[39]; // @[util.scala 114:43]
  wire [23:0] T_33770 = T_33766 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33771 = {T_33770,T_33765}; // @[Cat.scala 20:58]
  wire [64:0] T_33773 = {{1'd0}, T_33771}; // @[rob.scala 554:94]
  wire [63:0] T_33774 = T_33773[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33872 = {T_23555_T_33870_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_33867 = {{24'd0}, T_33872}; // @[rob.scala 899:26]
  wire [39:0] T_33879 = T_33867[39:0]; // @[rob.scala 906:20]
  wire  T_33880 = T_33879[39]; // @[util.scala 114:43]
  wire [23:0] T_33884 = T_33880 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33885 = {T_33884,T_33879}; // @[Cat.scala 20:58]
  wire [64:0] T_33887 = {{1'd0}, T_33885}; // @[rob.scala 554:94]
  wire [63:0] T_33888 = T_33887[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_33992 = {T_23558_T_33990_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_33981 = {{24'd0}, T_33992}; // @[rob.scala 899:26]
  wire [39:0] T_33993 = T_33981[39:0]; // @[rob.scala 906:20]
  wire  T_33994 = T_33993[39]; // @[util.scala 114:43]
  wire [23:0] T_33998 = T_33994 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_33999 = {T_33998,T_33993}; // @[Cat.scala 20:58]
  wire [64:0] T_34001 = {{1'd0}, T_33999}; // @[rob.scala 554:94]
  wire [63:0] T_34002 = T_34001[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34100 = {T_23555_T_34098_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_34095 = {{24'd0}, T_34100}; // @[rob.scala 899:26]
  wire [39:0] T_34107 = T_34095[39:0]; // @[rob.scala 906:20]
  wire  T_34108 = T_34107[39]; // @[util.scala 114:43]
  wire [23:0] T_34112 = T_34108 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34113 = {T_34112,T_34107}; // @[Cat.scala 20:58]
  wire [64:0] T_34115 = {{1'd0}, T_34113}; // @[rob.scala 554:94]
  wire [63:0] T_34116 = T_34115[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34220 = {T_23558_T_34218_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_34209 = {{24'd0}, T_34220}; // @[rob.scala 899:26]
  wire [39:0] T_34221 = T_34209[39:0]; // @[rob.scala 906:20]
  wire  T_34222 = T_34221[39]; // @[util.scala 114:43]
  wire [23:0] T_34226 = T_34222 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34227 = {T_34226,T_34221}; // @[Cat.scala 20:58]
  wire [64:0] T_34229 = {{1'd0}, T_34227}; // @[rob.scala 554:94]
  wire [63:0] T_34230 = T_34229[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34328 = {T_23555_T_34326_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_34323 = {{24'd0}, T_34328}; // @[rob.scala 899:26]
  wire [39:0] T_34335 = T_34323[39:0]; // @[rob.scala 906:20]
  wire  T_34336 = T_34335[39]; // @[util.scala 114:43]
  wire [23:0] T_34340 = T_34336 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34341 = {T_34340,T_34335}; // @[Cat.scala 20:58]
  wire [64:0] T_34343 = {{1'd0}, T_34341}; // @[rob.scala 554:94]
  wire [63:0] T_34344 = T_34343[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34448 = {T_23558_T_34446_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_34437 = {{24'd0}, T_34448}; // @[rob.scala 899:26]
  wire [39:0] T_34449 = T_34437[39:0]; // @[rob.scala 906:20]
  wire  T_34450 = T_34449[39]; // @[util.scala 114:43]
  wire [23:0] T_34454 = T_34450 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34455 = {T_34454,T_34449}; // @[Cat.scala 20:58]
  wire [64:0] T_34457 = {{1'd0}, T_34455}; // @[rob.scala 554:94]
  wire [63:0] T_34458 = T_34457[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34556 = {T_23555_T_34554_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_34551 = {{24'd0}, T_34556}; // @[rob.scala 899:26]
  wire [39:0] T_34563 = T_34551[39:0]; // @[rob.scala 906:20]
  wire  T_34564 = T_34563[39]; // @[util.scala 114:43]
  wire [23:0] T_34568 = T_34564 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34569 = {T_34568,T_34563}; // @[Cat.scala 20:58]
  wire [64:0] T_34571 = {{1'd0}, T_34569}; // @[rob.scala 554:94]
  wire [63:0] T_34572 = T_34571[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34676 = {T_23558_T_34674_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_34665 = {{24'd0}, T_34676}; // @[rob.scala 899:26]
  wire [39:0] T_34677 = T_34665[39:0]; // @[rob.scala 906:20]
  wire  T_34678 = T_34677[39]; // @[util.scala 114:43]
  wire [23:0] T_34682 = T_34678 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34683 = {T_34682,T_34677}; // @[Cat.scala 20:58]
  wire [64:0] T_34685 = {{1'd0}, T_34683}; // @[rob.scala 554:94]
  wire [63:0] T_34686 = T_34685[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34784 = {T_23555_T_34782_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_34779 = {{24'd0}, T_34784}; // @[rob.scala 899:26]
  wire [39:0] T_34791 = T_34779[39:0]; // @[rob.scala 906:20]
  wire  T_34792 = T_34791[39]; // @[util.scala 114:43]
  wire [23:0] T_34796 = T_34792 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34797 = {T_34796,T_34791}; // @[Cat.scala 20:58]
  wire [64:0] T_34799 = {{1'd0}, T_34797}; // @[rob.scala 554:94]
  wire [63:0] T_34800 = T_34799[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_34904 = {T_23558_T_34902_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_34893 = {{24'd0}, T_34904}; // @[rob.scala 899:26]
  wire [39:0] T_34905 = T_34893[39:0]; // @[rob.scala 906:20]
  wire  T_34906 = T_34905[39]; // @[util.scala 114:43]
  wire [23:0] T_34910 = T_34906 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_34911 = {T_34910,T_34905}; // @[Cat.scala 20:58]
  wire [64:0] T_34913 = {{1'd0}, T_34911}; // @[rob.scala 554:94]
  wire [63:0] T_34914 = T_34913[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_35012 = {T_23555_T_35010_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_35007 = {{24'd0}, T_35012}; // @[rob.scala 899:26]
  wire [39:0] T_35019 = T_35007[39:0]; // @[rob.scala 906:20]
  wire  T_35020 = T_35019[39]; // @[util.scala 114:43]
  wire [23:0] T_35024 = T_35020 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_35025 = {T_35024,T_35019}; // @[Cat.scala 20:58]
  wire [64:0] T_35027 = {{1'd0}, T_35025}; // @[rob.scala 554:94]
  wire [63:0] T_35028 = T_35027[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_35132 = {T_23558_T_35130_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_35121 = {{24'd0}, T_35132}; // @[rob.scala 899:26]
  wire [39:0] T_35133 = T_35121[39:0]; // @[rob.scala 906:20]
  wire  T_35134 = T_35133[39]; // @[util.scala 114:43]
  wire [23:0] T_35138 = T_35134 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_35139 = {T_35138,T_35133}; // @[Cat.scala 20:58]
  wire [64:0] T_35141 = {{1'd0}, T_35139}; // @[rob.scala 554:94]
  wire [63:0] T_35142 = T_35141[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_35240 = {T_23555_T_35238_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_35235 = {{24'd0}, T_35240}; // @[rob.scala 899:26]
  wire [39:0] T_35247 = T_35235[39:0]; // @[rob.scala 906:20]
  wire  T_35248 = T_35247[39]; // @[util.scala 114:43]
  wire [23:0] T_35252 = T_35248 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_35253 = {T_35252,T_35247}; // @[Cat.scala 20:58]
  wire [64:0] T_35255 = {{1'd0}, T_35253}; // @[rob.scala 554:94]
  wire [63:0] T_35256 = T_35255[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_35360 = {T_23558_T_35358_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_35349 = {{24'd0}, T_35360}; // @[rob.scala 899:26]
  wire [39:0] T_35361 = T_35349[39:0]; // @[rob.scala 906:20]
  wire  T_35362 = T_35361[39]; // @[util.scala 114:43]
  wire [23:0] T_35366 = T_35362 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_35367 = {T_35366,T_35361}; // @[Cat.scala 20:58]
  wire [64:0] T_35369 = {{1'd0}, T_35367}; // @[rob.scala 554:94]
  wire [63:0] T_35370 = T_35369[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_35468 = {T_23555_T_35466_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_35463 = {{24'd0}, T_35468}; // @[rob.scala 899:26]
  wire [39:0] T_35475 = T_35463[39:0]; // @[rob.scala 906:20]
  wire  T_35476 = T_35475[39]; // @[util.scala 114:43]
  wire [23:0] T_35480 = T_35476 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_35481 = {T_35480,T_35475}; // @[Cat.scala 20:58]
  wire [64:0] T_35483 = {{1'd0}, T_35481}; // @[rob.scala 554:94]
  wire [63:0] T_35484 = T_35483[63:0]; // @[rob.scala 554:94]
  wire [39:0] T_35588 = {T_23558_T_35586_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_35577 = {{24'd0}, T_35588}; // @[rob.scala 899:26]
  wire [39:0] T_35589 = T_35577[39:0]; // @[rob.scala 906:20]
  wire  T_35590 = T_35589[39]; // @[util.scala 114:43]
  wire [23:0] T_35594 = T_35590 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_35595 = {T_35594,T_35589}; // @[Cat.scala 20:58]
  wire [64:0] T_35597 = {{1'd0}, T_35595}; // @[rob.scala 554:94]
  wire [63:0] T_35598 = T_35597[63:0]; // @[rob.scala 554:94]
  reg  T_38110_0_valid;
  reg [1:0] T_38110_0_iw_state;
  reg [8:0] T_38110_0_uopc;
  reg [31:0] T_38110_0_inst;
  reg [39:0] T_38110_0_pc;
  reg [7:0] T_38110_0_fu_code;
  reg [3:0] T_38110_0_ctrl_br_type;
  reg [1:0] T_38110_0_ctrl_op1_sel;
  reg [2:0] T_38110_0_ctrl_op2_sel;
  reg [2:0] T_38110_0_ctrl_imm_sel;
  reg [3:0] T_38110_0_ctrl_op_fcn;
  reg  T_38110_0_ctrl_fcn_dw;
  reg  T_38110_0_ctrl_rf_wen;
  reg [2:0] T_38110_0_ctrl_csr_cmd;
  reg  T_38110_0_ctrl_is_load;
  reg  T_38110_0_ctrl_is_sta;
  reg  T_38110_0_ctrl_is_std;
  reg [1:0] T_38110_0_wakeup_delay;
  reg  T_38110_0_allocate_brtag;
  reg  T_38110_0_is_br_or_jmp;
  reg  T_38110_0_is_jump;
  reg  T_38110_0_is_jal;
  reg  T_38110_0_is_ret;
  reg  T_38110_0_is_call;
  reg [7:0] T_38110_0_br_mask;
  reg [2:0] T_38110_0_br_tag;
  reg  T_38110_0_br_prediction_bpd_predict_val;
  reg  T_38110_0_br_prediction_bpd_predict_taken;
  reg  T_38110_0_br_prediction_btb_hit;
  reg  T_38110_0_br_prediction_btb_predicted;
  reg  T_38110_0_br_prediction_is_br_or_jalr;
  reg  T_38110_0_stat_brjmp_mispredicted;
  reg  T_38110_0_stat_btb_made_pred;
  reg  T_38110_0_stat_btb_mispredicted;
  reg  T_38110_0_stat_bpd_made_pred;
  reg  T_38110_0_stat_bpd_mispredicted;
  reg [2:0] T_38110_0_fetch_pc_lob;
  reg [19:0] T_38110_0_imm_packed;
  reg [11:0] T_38110_0_csr_addr;
  reg [5:0] T_38110_0_rob_idx;
  reg [3:0] T_38110_0_ldq_idx;
  reg [3:0] T_38110_0_stq_idx;
  reg [4:0] T_38110_0_brob_idx;
  reg [6:0] T_38110_0_pdst;
  reg [6:0] T_38110_0_pop1;
  reg [6:0] T_38110_0_pop2;
  reg [6:0] T_38110_0_pop3;
  reg  T_38110_0_prs1_busy;
  reg  T_38110_0_prs2_busy;
  reg  T_38110_0_prs3_busy;
  reg [6:0] T_38110_0_stale_pdst;
  reg  T_38110_0_exception;
  reg [63:0] T_38110_0_exc_cause;
  reg  T_38110_0_bypassable;
  reg [3:0] T_38110_0_mem_cmd;
  reg [2:0] T_38110_0_mem_typ;
  reg  T_38110_0_is_fence;
  reg  T_38110_0_is_fencei;
  reg  T_38110_0_is_store;
  reg  T_38110_0_is_amo;
  reg  T_38110_0_is_load;
  reg  T_38110_0_is_unique;
  reg  T_38110_0_flush_on_commit;
  reg [5:0] T_38110_0_ldst;
  reg [5:0] T_38110_0_lrs1;
  reg [5:0] T_38110_0_lrs2;
  reg [5:0] T_38110_0_lrs3;
  reg  T_38110_0_ldst_val;
  reg [1:0] T_38110_0_dst_rtype;
  reg [1:0] T_38110_0_lrs1_rtype;
  reg [1:0] T_38110_0_lrs2_rtype;
  reg  T_38110_0_frs3_en;
  reg  T_38110_0_fp_val;
  reg  T_38110_0_fp_single;
  reg  T_38110_0_xcpt_if;
  reg  T_38110_0_replay_if;
  reg [63:0] T_38110_0_debug_wdata;
  reg [31:0] T_38110_0_debug_events_fetch_seq;
  reg  T_38110_1_valid;
  reg [1:0] T_38110_1_iw_state;
  reg [8:0] T_38110_1_uopc;
  reg [31:0] T_38110_1_inst;
  reg [39:0] T_38110_1_pc;
  reg [7:0] T_38110_1_fu_code;
  reg [3:0] T_38110_1_ctrl_br_type;
  reg [1:0] T_38110_1_ctrl_op1_sel;
  reg [2:0] T_38110_1_ctrl_op2_sel;
  reg [2:0] T_38110_1_ctrl_imm_sel;
  reg [3:0] T_38110_1_ctrl_op_fcn;
  reg  T_38110_1_ctrl_fcn_dw;
  reg  T_38110_1_ctrl_rf_wen;
  reg [2:0] T_38110_1_ctrl_csr_cmd;
  reg  T_38110_1_ctrl_is_load;
  reg  T_38110_1_ctrl_is_sta;
  reg  T_38110_1_ctrl_is_std;
  reg [1:0] T_38110_1_wakeup_delay;
  reg  T_38110_1_allocate_brtag;
  reg  T_38110_1_is_br_or_jmp;
  reg  T_38110_1_is_jump;
  reg  T_38110_1_is_jal;
  reg  T_38110_1_is_ret;
  reg  T_38110_1_is_call;
  reg [7:0] T_38110_1_br_mask;
  reg [2:0] T_38110_1_br_tag;
  reg  T_38110_1_br_prediction_bpd_predict_val;
  reg  T_38110_1_br_prediction_bpd_predict_taken;
  reg  T_38110_1_br_prediction_btb_hit;
  reg  T_38110_1_br_prediction_btb_predicted;
  reg  T_38110_1_br_prediction_is_br_or_jalr;
  reg  T_38110_1_stat_brjmp_mispredicted;
  reg  T_38110_1_stat_btb_made_pred;
  reg  T_38110_1_stat_btb_mispredicted;
  reg  T_38110_1_stat_bpd_made_pred;
  reg  T_38110_1_stat_bpd_mispredicted;
  reg [2:0] T_38110_1_fetch_pc_lob;
  reg [19:0] T_38110_1_imm_packed;
  reg [11:0] T_38110_1_csr_addr;
  reg [5:0] T_38110_1_rob_idx;
  reg [3:0] T_38110_1_ldq_idx;
  reg [3:0] T_38110_1_stq_idx;
  reg [4:0] T_38110_1_brob_idx;
  reg [6:0] T_38110_1_pdst;
  reg [6:0] T_38110_1_pop1;
  reg [6:0] T_38110_1_pop2;
  reg [6:0] T_38110_1_pop3;
  reg  T_38110_1_prs1_busy;
  reg  T_38110_1_prs2_busy;
  reg  T_38110_1_prs3_busy;
  reg [6:0] T_38110_1_stale_pdst;
  reg  T_38110_1_exception;
  reg [63:0] T_38110_1_exc_cause;
  reg  T_38110_1_bypassable;
  reg [3:0] T_38110_1_mem_cmd;
  reg [2:0] T_38110_1_mem_typ;
  reg  T_38110_1_is_fence;
  reg  T_38110_1_is_fencei;
  reg  T_38110_1_is_store;
  reg  T_38110_1_is_amo;
  reg  T_38110_1_is_load;
  reg  T_38110_1_is_unique;
  reg  T_38110_1_flush_on_commit;
  reg [5:0] T_38110_1_ldst;
  reg [5:0] T_38110_1_lrs1;
  reg [5:0] T_38110_1_lrs2;
  reg [5:0] T_38110_1_lrs3;
  reg  T_38110_1_ldst_val;
  reg [1:0] T_38110_1_dst_rtype;
  reg [1:0] T_38110_1_lrs1_rtype;
  reg [1:0] T_38110_1_lrs2_rtype;
  reg  T_38110_1_frs3_en;
  reg  T_38110_1_fp_val;
  reg  T_38110_1_fp_single;
  reg  T_38110_1_xcpt_if;
  reg  T_38110_1_replay_if;
  reg [63:0] T_38110_1_debug_wdata;
  reg [31:0] T_38110_1_debug_events_fetch_seq;
  reg  T_38110_2_valid;
  reg [1:0] T_38110_2_iw_state;
  reg [8:0] T_38110_2_uopc;
  reg [31:0] T_38110_2_inst;
  reg [39:0] T_38110_2_pc;
  reg [7:0] T_38110_2_fu_code;
  reg [3:0] T_38110_2_ctrl_br_type;
  reg [1:0] T_38110_2_ctrl_op1_sel;
  reg [2:0] T_38110_2_ctrl_op2_sel;
  reg [2:0] T_38110_2_ctrl_imm_sel;
  reg [3:0] T_38110_2_ctrl_op_fcn;
  reg  T_38110_2_ctrl_fcn_dw;
  reg  T_38110_2_ctrl_rf_wen;
  reg [2:0] T_38110_2_ctrl_csr_cmd;
  reg  T_38110_2_ctrl_is_load;
  reg  T_38110_2_ctrl_is_sta;
  reg  T_38110_2_ctrl_is_std;
  reg [1:0] T_38110_2_wakeup_delay;
  reg  T_38110_2_allocate_brtag;
  reg  T_38110_2_is_br_or_jmp;
  reg  T_38110_2_is_jump;
  reg  T_38110_2_is_jal;
  reg  T_38110_2_is_ret;
  reg  T_38110_2_is_call;
  reg [7:0] T_38110_2_br_mask;
  reg [2:0] T_38110_2_br_tag;
  reg  T_38110_2_br_prediction_bpd_predict_val;
  reg  T_38110_2_br_prediction_bpd_predict_taken;
  reg  T_38110_2_br_prediction_btb_hit;
  reg  T_38110_2_br_prediction_btb_predicted;
  reg  T_38110_2_br_prediction_is_br_or_jalr;
  reg  T_38110_2_stat_brjmp_mispredicted;
  reg  T_38110_2_stat_btb_made_pred;
  reg  T_38110_2_stat_btb_mispredicted;
  reg  T_38110_2_stat_bpd_made_pred;
  reg  T_38110_2_stat_bpd_mispredicted;
  reg [2:0] T_38110_2_fetch_pc_lob;
  reg [19:0] T_38110_2_imm_packed;
  reg [11:0] T_38110_2_csr_addr;
  reg [5:0] T_38110_2_rob_idx;
  reg [3:0] T_38110_2_ldq_idx;
  reg [3:0] T_38110_2_stq_idx;
  reg [4:0] T_38110_2_brob_idx;
  reg [6:0] T_38110_2_pdst;
  reg [6:0] T_38110_2_pop1;
  reg [6:0] T_38110_2_pop2;
  reg [6:0] T_38110_2_pop3;
  reg  T_38110_2_prs1_busy;
  reg  T_38110_2_prs2_busy;
  reg  T_38110_2_prs3_busy;
  reg [6:0] T_38110_2_stale_pdst;
  reg  T_38110_2_exception;
  reg [63:0] T_38110_2_exc_cause;
  reg  T_38110_2_bypassable;
  reg [3:0] T_38110_2_mem_cmd;
  reg [2:0] T_38110_2_mem_typ;
  reg  T_38110_2_is_fence;
  reg  T_38110_2_is_fencei;
  reg  T_38110_2_is_store;
  reg  T_38110_2_is_amo;
  reg  T_38110_2_is_load;
  reg  T_38110_2_is_unique;
  reg  T_38110_2_flush_on_commit;
  reg [5:0] T_38110_2_ldst;
  reg [5:0] T_38110_2_lrs1;
  reg [5:0] T_38110_2_lrs2;
  reg [5:0] T_38110_2_lrs3;
  reg  T_38110_2_ldst_val;
  reg [1:0] T_38110_2_dst_rtype;
  reg [1:0] T_38110_2_lrs1_rtype;
  reg [1:0] T_38110_2_lrs2_rtype;
  reg  T_38110_2_frs3_en;
  reg  T_38110_2_fp_val;
  reg  T_38110_2_fp_single;
  reg  T_38110_2_xcpt_if;
  reg  T_38110_2_replay_if;
  reg [63:0] T_38110_2_debug_wdata;
  reg [31:0] T_38110_2_debug_events_fetch_seq;
  reg  T_38110_3_valid;
  reg [1:0] T_38110_3_iw_state;
  reg [8:0] T_38110_3_uopc;
  reg [31:0] T_38110_3_inst;
  reg [39:0] T_38110_3_pc;
  reg [7:0] T_38110_3_fu_code;
  reg [3:0] T_38110_3_ctrl_br_type;
  reg [1:0] T_38110_3_ctrl_op1_sel;
  reg [2:0] T_38110_3_ctrl_op2_sel;
  reg [2:0] T_38110_3_ctrl_imm_sel;
  reg [3:0] T_38110_3_ctrl_op_fcn;
  reg  T_38110_3_ctrl_fcn_dw;
  reg  T_38110_3_ctrl_rf_wen;
  reg [2:0] T_38110_3_ctrl_csr_cmd;
  reg  T_38110_3_ctrl_is_load;
  reg  T_38110_3_ctrl_is_sta;
  reg  T_38110_3_ctrl_is_std;
  reg [1:0] T_38110_3_wakeup_delay;
  reg  T_38110_3_allocate_brtag;
  reg  T_38110_3_is_br_or_jmp;
  reg  T_38110_3_is_jump;
  reg  T_38110_3_is_jal;
  reg  T_38110_3_is_ret;
  reg  T_38110_3_is_call;
  reg [7:0] T_38110_3_br_mask;
  reg [2:0] T_38110_3_br_tag;
  reg  T_38110_3_br_prediction_bpd_predict_val;
  reg  T_38110_3_br_prediction_bpd_predict_taken;
  reg  T_38110_3_br_prediction_btb_hit;
  reg  T_38110_3_br_prediction_btb_predicted;
  reg  T_38110_3_br_prediction_is_br_or_jalr;
  reg  T_38110_3_stat_brjmp_mispredicted;
  reg  T_38110_3_stat_btb_made_pred;
  reg  T_38110_3_stat_btb_mispredicted;
  reg  T_38110_3_stat_bpd_made_pred;
  reg  T_38110_3_stat_bpd_mispredicted;
  reg [2:0] T_38110_3_fetch_pc_lob;
  reg [19:0] T_38110_3_imm_packed;
  reg [11:0] T_38110_3_csr_addr;
  reg [5:0] T_38110_3_rob_idx;
  reg [3:0] T_38110_3_ldq_idx;
  reg [3:0] T_38110_3_stq_idx;
  reg [4:0] T_38110_3_brob_idx;
  reg [6:0] T_38110_3_pdst;
  reg [6:0] T_38110_3_pop1;
  reg [6:0] T_38110_3_pop2;
  reg [6:0] T_38110_3_pop3;
  reg  T_38110_3_prs1_busy;
  reg  T_38110_3_prs2_busy;
  reg  T_38110_3_prs3_busy;
  reg [6:0] T_38110_3_stale_pdst;
  reg  T_38110_3_exception;
  reg [63:0] T_38110_3_exc_cause;
  reg  T_38110_3_bypassable;
  reg [3:0] T_38110_3_mem_cmd;
  reg [2:0] T_38110_3_mem_typ;
  reg  T_38110_3_is_fence;
  reg  T_38110_3_is_fencei;
  reg  T_38110_3_is_store;
  reg  T_38110_3_is_amo;
  reg  T_38110_3_is_load;
  reg  T_38110_3_is_unique;
  reg  T_38110_3_flush_on_commit;
  reg [5:0] T_38110_3_ldst;
  reg [5:0] T_38110_3_lrs1;
  reg [5:0] T_38110_3_lrs2;
  reg [5:0] T_38110_3_lrs3;
  reg  T_38110_3_ldst_val;
  reg [1:0] T_38110_3_dst_rtype;
  reg [1:0] T_38110_3_lrs1_rtype;
  reg [1:0] T_38110_3_lrs2_rtype;
  reg  T_38110_3_frs3_en;
  reg  T_38110_3_fp_val;
  reg  T_38110_3_fp_single;
  reg  T_38110_3_xcpt_if;
  reg  T_38110_3_replay_if;
  reg [63:0] T_38110_3_debug_wdata;
  reg [31:0] T_38110_3_debug_events_fetch_seq;
  reg  T_38110_4_valid;
  reg [1:0] T_38110_4_iw_state;
  reg [8:0] T_38110_4_uopc;
  reg [31:0] T_38110_4_inst;
  reg [39:0] T_38110_4_pc;
  reg [7:0] T_38110_4_fu_code;
  reg [3:0] T_38110_4_ctrl_br_type;
  reg [1:0] T_38110_4_ctrl_op1_sel;
  reg [2:0] T_38110_4_ctrl_op2_sel;
  reg [2:0] T_38110_4_ctrl_imm_sel;
  reg [3:0] T_38110_4_ctrl_op_fcn;
  reg  T_38110_4_ctrl_fcn_dw;
  reg  T_38110_4_ctrl_rf_wen;
  reg [2:0] T_38110_4_ctrl_csr_cmd;
  reg  T_38110_4_ctrl_is_load;
  reg  T_38110_4_ctrl_is_sta;
  reg  T_38110_4_ctrl_is_std;
  reg [1:0] T_38110_4_wakeup_delay;
  reg  T_38110_4_allocate_brtag;
  reg  T_38110_4_is_br_or_jmp;
  reg  T_38110_4_is_jump;
  reg  T_38110_4_is_jal;
  reg  T_38110_4_is_ret;
  reg  T_38110_4_is_call;
  reg [7:0] T_38110_4_br_mask;
  reg [2:0] T_38110_4_br_tag;
  reg  T_38110_4_br_prediction_bpd_predict_val;
  reg  T_38110_4_br_prediction_bpd_predict_taken;
  reg  T_38110_4_br_prediction_btb_hit;
  reg  T_38110_4_br_prediction_btb_predicted;
  reg  T_38110_4_br_prediction_is_br_or_jalr;
  reg  T_38110_4_stat_brjmp_mispredicted;
  reg  T_38110_4_stat_btb_made_pred;
  reg  T_38110_4_stat_btb_mispredicted;
  reg  T_38110_4_stat_bpd_made_pred;
  reg  T_38110_4_stat_bpd_mispredicted;
  reg [2:0] T_38110_4_fetch_pc_lob;
  reg [19:0] T_38110_4_imm_packed;
  reg [11:0] T_38110_4_csr_addr;
  reg [5:0] T_38110_4_rob_idx;
  reg [3:0] T_38110_4_ldq_idx;
  reg [3:0] T_38110_4_stq_idx;
  reg [4:0] T_38110_4_brob_idx;
  reg [6:0] T_38110_4_pdst;
  reg [6:0] T_38110_4_pop1;
  reg [6:0] T_38110_4_pop2;
  reg [6:0] T_38110_4_pop3;
  reg  T_38110_4_prs1_busy;
  reg  T_38110_4_prs2_busy;
  reg  T_38110_4_prs3_busy;
  reg [6:0] T_38110_4_stale_pdst;
  reg  T_38110_4_exception;
  reg [63:0] T_38110_4_exc_cause;
  reg  T_38110_4_bypassable;
  reg [3:0] T_38110_4_mem_cmd;
  reg [2:0] T_38110_4_mem_typ;
  reg  T_38110_4_is_fence;
  reg  T_38110_4_is_fencei;
  reg  T_38110_4_is_store;
  reg  T_38110_4_is_amo;
  reg  T_38110_4_is_load;
  reg  T_38110_4_is_unique;
  reg  T_38110_4_flush_on_commit;
  reg [5:0] T_38110_4_ldst;
  reg [5:0] T_38110_4_lrs1;
  reg [5:0] T_38110_4_lrs2;
  reg [5:0] T_38110_4_lrs3;
  reg  T_38110_4_ldst_val;
  reg [1:0] T_38110_4_dst_rtype;
  reg [1:0] T_38110_4_lrs1_rtype;
  reg [1:0] T_38110_4_lrs2_rtype;
  reg  T_38110_4_frs3_en;
  reg  T_38110_4_fp_val;
  reg  T_38110_4_fp_single;
  reg  T_38110_4_xcpt_if;
  reg  T_38110_4_replay_if;
  reg [63:0] T_38110_4_debug_wdata;
  reg [31:0] T_38110_4_debug_events_fetch_seq;
  reg  T_38110_5_valid;
  reg [1:0] T_38110_5_iw_state;
  reg [8:0] T_38110_5_uopc;
  reg [31:0] T_38110_5_inst;
  reg [39:0] T_38110_5_pc;
  reg [7:0] T_38110_5_fu_code;
  reg [3:0] T_38110_5_ctrl_br_type;
  reg [1:0] T_38110_5_ctrl_op1_sel;
  reg [2:0] T_38110_5_ctrl_op2_sel;
  reg [2:0] T_38110_5_ctrl_imm_sel;
  reg [3:0] T_38110_5_ctrl_op_fcn;
  reg  T_38110_5_ctrl_fcn_dw;
  reg  T_38110_5_ctrl_rf_wen;
  reg [2:0] T_38110_5_ctrl_csr_cmd;
  reg  T_38110_5_ctrl_is_load;
  reg  T_38110_5_ctrl_is_sta;
  reg  T_38110_5_ctrl_is_std;
  reg [1:0] T_38110_5_wakeup_delay;
  reg  T_38110_5_allocate_brtag;
  reg  T_38110_5_is_br_or_jmp;
  reg  T_38110_5_is_jump;
  reg  T_38110_5_is_jal;
  reg  T_38110_5_is_ret;
  reg  T_38110_5_is_call;
  reg [7:0] T_38110_5_br_mask;
  reg [2:0] T_38110_5_br_tag;
  reg  T_38110_5_br_prediction_bpd_predict_val;
  reg  T_38110_5_br_prediction_bpd_predict_taken;
  reg  T_38110_5_br_prediction_btb_hit;
  reg  T_38110_5_br_prediction_btb_predicted;
  reg  T_38110_5_br_prediction_is_br_or_jalr;
  reg  T_38110_5_stat_brjmp_mispredicted;
  reg  T_38110_5_stat_btb_made_pred;
  reg  T_38110_5_stat_btb_mispredicted;
  reg  T_38110_5_stat_bpd_made_pred;
  reg  T_38110_5_stat_bpd_mispredicted;
  reg [2:0] T_38110_5_fetch_pc_lob;
  reg [19:0] T_38110_5_imm_packed;
  reg [11:0] T_38110_5_csr_addr;
  reg [5:0] T_38110_5_rob_idx;
  reg [3:0] T_38110_5_ldq_idx;
  reg [3:0] T_38110_5_stq_idx;
  reg [4:0] T_38110_5_brob_idx;
  reg [6:0] T_38110_5_pdst;
  reg [6:0] T_38110_5_pop1;
  reg [6:0] T_38110_5_pop2;
  reg [6:0] T_38110_5_pop3;
  reg  T_38110_5_prs1_busy;
  reg  T_38110_5_prs2_busy;
  reg  T_38110_5_prs3_busy;
  reg [6:0] T_38110_5_stale_pdst;
  reg  T_38110_5_exception;
  reg [63:0] T_38110_5_exc_cause;
  reg  T_38110_5_bypassable;
  reg [3:0] T_38110_5_mem_cmd;
  reg [2:0] T_38110_5_mem_typ;
  reg  T_38110_5_is_fence;
  reg  T_38110_5_is_fencei;
  reg  T_38110_5_is_store;
  reg  T_38110_5_is_amo;
  reg  T_38110_5_is_load;
  reg  T_38110_5_is_unique;
  reg  T_38110_5_flush_on_commit;
  reg [5:0] T_38110_5_ldst;
  reg [5:0] T_38110_5_lrs1;
  reg [5:0] T_38110_5_lrs2;
  reg [5:0] T_38110_5_lrs3;
  reg  T_38110_5_ldst_val;
  reg [1:0] T_38110_5_dst_rtype;
  reg [1:0] T_38110_5_lrs1_rtype;
  reg [1:0] T_38110_5_lrs2_rtype;
  reg  T_38110_5_frs3_en;
  reg  T_38110_5_fp_val;
  reg  T_38110_5_fp_single;
  reg  T_38110_5_xcpt_if;
  reg  T_38110_5_replay_if;
  reg [63:0] T_38110_5_debug_wdata;
  reg [31:0] T_38110_5_debug_events_fetch_seq;
  reg  T_38110_6_valid;
  reg [1:0] T_38110_6_iw_state;
  reg [8:0] T_38110_6_uopc;
  reg [31:0] T_38110_6_inst;
  reg [39:0] T_38110_6_pc;
  reg [7:0] T_38110_6_fu_code;
  reg [3:0] T_38110_6_ctrl_br_type;
  reg [1:0] T_38110_6_ctrl_op1_sel;
  reg [2:0] T_38110_6_ctrl_op2_sel;
  reg [2:0] T_38110_6_ctrl_imm_sel;
  reg [3:0] T_38110_6_ctrl_op_fcn;
  reg  T_38110_6_ctrl_fcn_dw;
  reg  T_38110_6_ctrl_rf_wen;
  reg [2:0] T_38110_6_ctrl_csr_cmd;
  reg  T_38110_6_ctrl_is_load;
  reg  T_38110_6_ctrl_is_sta;
  reg  T_38110_6_ctrl_is_std;
  reg [1:0] T_38110_6_wakeup_delay;
  reg  T_38110_6_allocate_brtag;
  reg  T_38110_6_is_br_or_jmp;
  reg  T_38110_6_is_jump;
  reg  T_38110_6_is_jal;
  reg  T_38110_6_is_ret;
  reg  T_38110_6_is_call;
  reg [7:0] T_38110_6_br_mask;
  reg [2:0] T_38110_6_br_tag;
  reg  T_38110_6_br_prediction_bpd_predict_val;
  reg  T_38110_6_br_prediction_bpd_predict_taken;
  reg  T_38110_6_br_prediction_btb_hit;
  reg  T_38110_6_br_prediction_btb_predicted;
  reg  T_38110_6_br_prediction_is_br_or_jalr;
  reg  T_38110_6_stat_brjmp_mispredicted;
  reg  T_38110_6_stat_btb_made_pred;
  reg  T_38110_6_stat_btb_mispredicted;
  reg  T_38110_6_stat_bpd_made_pred;
  reg  T_38110_6_stat_bpd_mispredicted;
  reg [2:0] T_38110_6_fetch_pc_lob;
  reg [19:0] T_38110_6_imm_packed;
  reg [11:0] T_38110_6_csr_addr;
  reg [5:0] T_38110_6_rob_idx;
  reg [3:0] T_38110_6_ldq_idx;
  reg [3:0] T_38110_6_stq_idx;
  reg [4:0] T_38110_6_brob_idx;
  reg [6:0] T_38110_6_pdst;
  reg [6:0] T_38110_6_pop1;
  reg [6:0] T_38110_6_pop2;
  reg [6:0] T_38110_6_pop3;
  reg  T_38110_6_prs1_busy;
  reg  T_38110_6_prs2_busy;
  reg  T_38110_6_prs3_busy;
  reg [6:0] T_38110_6_stale_pdst;
  reg  T_38110_6_exception;
  reg [63:0] T_38110_6_exc_cause;
  reg  T_38110_6_bypassable;
  reg [3:0] T_38110_6_mem_cmd;
  reg [2:0] T_38110_6_mem_typ;
  reg  T_38110_6_is_fence;
  reg  T_38110_6_is_fencei;
  reg  T_38110_6_is_store;
  reg  T_38110_6_is_amo;
  reg  T_38110_6_is_load;
  reg  T_38110_6_is_unique;
  reg  T_38110_6_flush_on_commit;
  reg [5:0] T_38110_6_ldst;
  reg [5:0] T_38110_6_lrs1;
  reg [5:0] T_38110_6_lrs2;
  reg [5:0] T_38110_6_lrs3;
  reg  T_38110_6_ldst_val;
  reg [1:0] T_38110_6_dst_rtype;
  reg [1:0] T_38110_6_lrs1_rtype;
  reg [1:0] T_38110_6_lrs2_rtype;
  reg  T_38110_6_frs3_en;
  reg  T_38110_6_fp_val;
  reg  T_38110_6_fp_single;
  reg  T_38110_6_xcpt_if;
  reg  T_38110_6_replay_if;
  reg [63:0] T_38110_6_debug_wdata;
  reg [31:0] T_38110_6_debug_events_fetch_seq;
  reg  T_38110_7_valid;
  reg [1:0] T_38110_7_iw_state;
  reg [8:0] T_38110_7_uopc;
  reg [31:0] T_38110_7_inst;
  reg [39:0] T_38110_7_pc;
  reg [7:0] T_38110_7_fu_code;
  reg [3:0] T_38110_7_ctrl_br_type;
  reg [1:0] T_38110_7_ctrl_op1_sel;
  reg [2:0] T_38110_7_ctrl_op2_sel;
  reg [2:0] T_38110_7_ctrl_imm_sel;
  reg [3:0] T_38110_7_ctrl_op_fcn;
  reg  T_38110_7_ctrl_fcn_dw;
  reg  T_38110_7_ctrl_rf_wen;
  reg [2:0] T_38110_7_ctrl_csr_cmd;
  reg  T_38110_7_ctrl_is_load;
  reg  T_38110_7_ctrl_is_sta;
  reg  T_38110_7_ctrl_is_std;
  reg [1:0] T_38110_7_wakeup_delay;
  reg  T_38110_7_allocate_brtag;
  reg  T_38110_7_is_br_or_jmp;
  reg  T_38110_7_is_jump;
  reg  T_38110_7_is_jal;
  reg  T_38110_7_is_ret;
  reg  T_38110_7_is_call;
  reg [7:0] T_38110_7_br_mask;
  reg [2:0] T_38110_7_br_tag;
  reg  T_38110_7_br_prediction_bpd_predict_val;
  reg  T_38110_7_br_prediction_bpd_predict_taken;
  reg  T_38110_7_br_prediction_btb_hit;
  reg  T_38110_7_br_prediction_btb_predicted;
  reg  T_38110_7_br_prediction_is_br_or_jalr;
  reg  T_38110_7_stat_brjmp_mispredicted;
  reg  T_38110_7_stat_btb_made_pred;
  reg  T_38110_7_stat_btb_mispredicted;
  reg  T_38110_7_stat_bpd_made_pred;
  reg  T_38110_7_stat_bpd_mispredicted;
  reg [2:0] T_38110_7_fetch_pc_lob;
  reg [19:0] T_38110_7_imm_packed;
  reg [11:0] T_38110_7_csr_addr;
  reg [5:0] T_38110_7_rob_idx;
  reg [3:0] T_38110_7_ldq_idx;
  reg [3:0] T_38110_7_stq_idx;
  reg [4:0] T_38110_7_brob_idx;
  reg [6:0] T_38110_7_pdst;
  reg [6:0] T_38110_7_pop1;
  reg [6:0] T_38110_7_pop2;
  reg [6:0] T_38110_7_pop3;
  reg  T_38110_7_prs1_busy;
  reg  T_38110_7_prs2_busy;
  reg  T_38110_7_prs3_busy;
  reg [6:0] T_38110_7_stale_pdst;
  reg  T_38110_7_exception;
  reg [63:0] T_38110_7_exc_cause;
  reg  T_38110_7_bypassable;
  reg [3:0] T_38110_7_mem_cmd;
  reg [2:0] T_38110_7_mem_typ;
  reg  T_38110_7_is_fence;
  reg  T_38110_7_is_fencei;
  reg  T_38110_7_is_store;
  reg  T_38110_7_is_amo;
  reg  T_38110_7_is_load;
  reg  T_38110_7_is_unique;
  reg  T_38110_7_flush_on_commit;
  reg [5:0] T_38110_7_ldst;
  reg [5:0] T_38110_7_lrs1;
  reg [5:0] T_38110_7_lrs2;
  reg [5:0] T_38110_7_lrs3;
  reg  T_38110_7_ldst_val;
  reg [1:0] T_38110_7_dst_rtype;
  reg [1:0] T_38110_7_lrs1_rtype;
  reg [1:0] T_38110_7_lrs2_rtype;
  reg  T_38110_7_frs3_en;
  reg  T_38110_7_fp_val;
  reg  T_38110_7_fp_single;
  reg  T_38110_7_xcpt_if;
  reg  T_38110_7_replay_if;
  reg [63:0] T_38110_7_debug_wdata;
  reg [31:0] T_38110_7_debug_events_fetch_seq;
  reg  T_38110_8_valid;
  reg [1:0] T_38110_8_iw_state;
  reg [8:0] T_38110_8_uopc;
  reg [31:0] T_38110_8_inst;
  reg [39:0] T_38110_8_pc;
  reg [7:0] T_38110_8_fu_code;
  reg [3:0] T_38110_8_ctrl_br_type;
  reg [1:0] T_38110_8_ctrl_op1_sel;
  reg [2:0] T_38110_8_ctrl_op2_sel;
  reg [2:0] T_38110_8_ctrl_imm_sel;
  reg [3:0] T_38110_8_ctrl_op_fcn;
  reg  T_38110_8_ctrl_fcn_dw;
  reg  T_38110_8_ctrl_rf_wen;
  reg [2:0] T_38110_8_ctrl_csr_cmd;
  reg  T_38110_8_ctrl_is_load;
  reg  T_38110_8_ctrl_is_sta;
  reg  T_38110_8_ctrl_is_std;
  reg [1:0] T_38110_8_wakeup_delay;
  reg  T_38110_8_allocate_brtag;
  reg  T_38110_8_is_br_or_jmp;
  reg  T_38110_8_is_jump;
  reg  T_38110_8_is_jal;
  reg  T_38110_8_is_ret;
  reg  T_38110_8_is_call;
  reg [7:0] T_38110_8_br_mask;
  reg [2:0] T_38110_8_br_tag;
  reg  T_38110_8_br_prediction_bpd_predict_val;
  reg  T_38110_8_br_prediction_bpd_predict_taken;
  reg  T_38110_8_br_prediction_btb_hit;
  reg  T_38110_8_br_prediction_btb_predicted;
  reg  T_38110_8_br_prediction_is_br_or_jalr;
  reg  T_38110_8_stat_brjmp_mispredicted;
  reg  T_38110_8_stat_btb_made_pred;
  reg  T_38110_8_stat_btb_mispredicted;
  reg  T_38110_8_stat_bpd_made_pred;
  reg  T_38110_8_stat_bpd_mispredicted;
  reg [2:0] T_38110_8_fetch_pc_lob;
  reg [19:0] T_38110_8_imm_packed;
  reg [11:0] T_38110_8_csr_addr;
  reg [5:0] T_38110_8_rob_idx;
  reg [3:0] T_38110_8_ldq_idx;
  reg [3:0] T_38110_8_stq_idx;
  reg [4:0] T_38110_8_brob_idx;
  reg [6:0] T_38110_8_pdst;
  reg [6:0] T_38110_8_pop1;
  reg [6:0] T_38110_8_pop2;
  reg [6:0] T_38110_8_pop3;
  reg  T_38110_8_prs1_busy;
  reg  T_38110_8_prs2_busy;
  reg  T_38110_8_prs3_busy;
  reg [6:0] T_38110_8_stale_pdst;
  reg  T_38110_8_exception;
  reg [63:0] T_38110_8_exc_cause;
  reg  T_38110_8_bypassable;
  reg [3:0] T_38110_8_mem_cmd;
  reg [2:0] T_38110_8_mem_typ;
  reg  T_38110_8_is_fence;
  reg  T_38110_8_is_fencei;
  reg  T_38110_8_is_store;
  reg  T_38110_8_is_amo;
  reg  T_38110_8_is_load;
  reg  T_38110_8_is_unique;
  reg  T_38110_8_flush_on_commit;
  reg [5:0] T_38110_8_ldst;
  reg [5:0] T_38110_8_lrs1;
  reg [5:0] T_38110_8_lrs2;
  reg [5:0] T_38110_8_lrs3;
  reg  T_38110_8_ldst_val;
  reg [1:0] T_38110_8_dst_rtype;
  reg [1:0] T_38110_8_lrs1_rtype;
  reg [1:0] T_38110_8_lrs2_rtype;
  reg  T_38110_8_frs3_en;
  reg  T_38110_8_fp_val;
  reg  T_38110_8_fp_single;
  reg  T_38110_8_xcpt_if;
  reg  T_38110_8_replay_if;
  reg [63:0] T_38110_8_debug_wdata;
  reg [31:0] T_38110_8_debug_events_fetch_seq;
  reg  T_38110_9_valid;
  reg [1:0] T_38110_9_iw_state;
  reg [8:0] T_38110_9_uopc;
  reg [31:0] T_38110_9_inst;
  reg [39:0] T_38110_9_pc;
  reg [7:0] T_38110_9_fu_code;
  reg [3:0] T_38110_9_ctrl_br_type;
  reg [1:0] T_38110_9_ctrl_op1_sel;
  reg [2:0] T_38110_9_ctrl_op2_sel;
  reg [2:0] T_38110_9_ctrl_imm_sel;
  reg [3:0] T_38110_9_ctrl_op_fcn;
  reg  T_38110_9_ctrl_fcn_dw;
  reg  T_38110_9_ctrl_rf_wen;
  reg [2:0] T_38110_9_ctrl_csr_cmd;
  reg  T_38110_9_ctrl_is_load;
  reg  T_38110_9_ctrl_is_sta;
  reg  T_38110_9_ctrl_is_std;
  reg [1:0] T_38110_9_wakeup_delay;
  reg  T_38110_9_allocate_brtag;
  reg  T_38110_9_is_br_or_jmp;
  reg  T_38110_9_is_jump;
  reg  T_38110_9_is_jal;
  reg  T_38110_9_is_ret;
  reg  T_38110_9_is_call;
  reg [7:0] T_38110_9_br_mask;
  reg [2:0] T_38110_9_br_tag;
  reg  T_38110_9_br_prediction_bpd_predict_val;
  reg  T_38110_9_br_prediction_bpd_predict_taken;
  reg  T_38110_9_br_prediction_btb_hit;
  reg  T_38110_9_br_prediction_btb_predicted;
  reg  T_38110_9_br_prediction_is_br_or_jalr;
  reg  T_38110_9_stat_brjmp_mispredicted;
  reg  T_38110_9_stat_btb_made_pred;
  reg  T_38110_9_stat_btb_mispredicted;
  reg  T_38110_9_stat_bpd_made_pred;
  reg  T_38110_9_stat_bpd_mispredicted;
  reg [2:0] T_38110_9_fetch_pc_lob;
  reg [19:0] T_38110_9_imm_packed;
  reg [11:0] T_38110_9_csr_addr;
  reg [5:0] T_38110_9_rob_idx;
  reg [3:0] T_38110_9_ldq_idx;
  reg [3:0] T_38110_9_stq_idx;
  reg [4:0] T_38110_9_brob_idx;
  reg [6:0] T_38110_9_pdst;
  reg [6:0] T_38110_9_pop1;
  reg [6:0] T_38110_9_pop2;
  reg [6:0] T_38110_9_pop3;
  reg  T_38110_9_prs1_busy;
  reg  T_38110_9_prs2_busy;
  reg  T_38110_9_prs3_busy;
  reg [6:0] T_38110_9_stale_pdst;
  reg  T_38110_9_exception;
  reg [63:0] T_38110_9_exc_cause;
  reg  T_38110_9_bypassable;
  reg [3:0] T_38110_9_mem_cmd;
  reg [2:0] T_38110_9_mem_typ;
  reg  T_38110_9_is_fence;
  reg  T_38110_9_is_fencei;
  reg  T_38110_9_is_store;
  reg  T_38110_9_is_amo;
  reg  T_38110_9_is_load;
  reg  T_38110_9_is_unique;
  reg  T_38110_9_flush_on_commit;
  reg [5:0] T_38110_9_ldst;
  reg [5:0] T_38110_9_lrs1;
  reg [5:0] T_38110_9_lrs2;
  reg [5:0] T_38110_9_lrs3;
  reg  T_38110_9_ldst_val;
  reg [1:0] T_38110_9_dst_rtype;
  reg [1:0] T_38110_9_lrs1_rtype;
  reg [1:0] T_38110_9_lrs2_rtype;
  reg  T_38110_9_frs3_en;
  reg  T_38110_9_fp_val;
  reg  T_38110_9_fp_single;
  reg  T_38110_9_xcpt_if;
  reg  T_38110_9_replay_if;
  reg [63:0] T_38110_9_debug_wdata;
  reg [31:0] T_38110_9_debug_events_fetch_seq;
  reg  T_38110_10_valid;
  reg [1:0] T_38110_10_iw_state;
  reg [8:0] T_38110_10_uopc;
  reg [31:0] T_38110_10_inst;
  reg [39:0] T_38110_10_pc;
  reg [7:0] T_38110_10_fu_code;
  reg [3:0] T_38110_10_ctrl_br_type;
  reg [1:0] T_38110_10_ctrl_op1_sel;
  reg [2:0] T_38110_10_ctrl_op2_sel;
  reg [2:0] T_38110_10_ctrl_imm_sel;
  reg [3:0] T_38110_10_ctrl_op_fcn;
  reg  T_38110_10_ctrl_fcn_dw;
  reg  T_38110_10_ctrl_rf_wen;
  reg [2:0] T_38110_10_ctrl_csr_cmd;
  reg  T_38110_10_ctrl_is_load;
  reg  T_38110_10_ctrl_is_sta;
  reg  T_38110_10_ctrl_is_std;
  reg [1:0] T_38110_10_wakeup_delay;
  reg  T_38110_10_allocate_brtag;
  reg  T_38110_10_is_br_or_jmp;
  reg  T_38110_10_is_jump;
  reg  T_38110_10_is_jal;
  reg  T_38110_10_is_ret;
  reg  T_38110_10_is_call;
  reg [7:0] T_38110_10_br_mask;
  reg [2:0] T_38110_10_br_tag;
  reg  T_38110_10_br_prediction_bpd_predict_val;
  reg  T_38110_10_br_prediction_bpd_predict_taken;
  reg  T_38110_10_br_prediction_btb_hit;
  reg  T_38110_10_br_prediction_btb_predicted;
  reg  T_38110_10_br_prediction_is_br_or_jalr;
  reg  T_38110_10_stat_brjmp_mispredicted;
  reg  T_38110_10_stat_btb_made_pred;
  reg  T_38110_10_stat_btb_mispredicted;
  reg  T_38110_10_stat_bpd_made_pred;
  reg  T_38110_10_stat_bpd_mispredicted;
  reg [2:0] T_38110_10_fetch_pc_lob;
  reg [19:0] T_38110_10_imm_packed;
  reg [11:0] T_38110_10_csr_addr;
  reg [5:0] T_38110_10_rob_idx;
  reg [3:0] T_38110_10_ldq_idx;
  reg [3:0] T_38110_10_stq_idx;
  reg [4:0] T_38110_10_brob_idx;
  reg [6:0] T_38110_10_pdst;
  reg [6:0] T_38110_10_pop1;
  reg [6:0] T_38110_10_pop2;
  reg [6:0] T_38110_10_pop3;
  reg  T_38110_10_prs1_busy;
  reg  T_38110_10_prs2_busy;
  reg  T_38110_10_prs3_busy;
  reg [6:0] T_38110_10_stale_pdst;
  reg  T_38110_10_exception;
  reg [63:0] T_38110_10_exc_cause;
  reg  T_38110_10_bypassable;
  reg [3:0] T_38110_10_mem_cmd;
  reg [2:0] T_38110_10_mem_typ;
  reg  T_38110_10_is_fence;
  reg  T_38110_10_is_fencei;
  reg  T_38110_10_is_store;
  reg  T_38110_10_is_amo;
  reg  T_38110_10_is_load;
  reg  T_38110_10_is_unique;
  reg  T_38110_10_flush_on_commit;
  reg [5:0] T_38110_10_ldst;
  reg [5:0] T_38110_10_lrs1;
  reg [5:0] T_38110_10_lrs2;
  reg [5:0] T_38110_10_lrs3;
  reg  T_38110_10_ldst_val;
  reg [1:0] T_38110_10_dst_rtype;
  reg [1:0] T_38110_10_lrs1_rtype;
  reg [1:0] T_38110_10_lrs2_rtype;
  reg  T_38110_10_frs3_en;
  reg  T_38110_10_fp_val;
  reg  T_38110_10_fp_single;
  reg  T_38110_10_xcpt_if;
  reg  T_38110_10_replay_if;
  reg [63:0] T_38110_10_debug_wdata;
  reg [31:0] T_38110_10_debug_events_fetch_seq;
  reg  T_38110_11_valid;
  reg [1:0] T_38110_11_iw_state;
  reg [8:0] T_38110_11_uopc;
  reg [31:0] T_38110_11_inst;
  reg [39:0] T_38110_11_pc;
  reg [7:0] T_38110_11_fu_code;
  reg [3:0] T_38110_11_ctrl_br_type;
  reg [1:0] T_38110_11_ctrl_op1_sel;
  reg [2:0] T_38110_11_ctrl_op2_sel;
  reg [2:0] T_38110_11_ctrl_imm_sel;
  reg [3:0] T_38110_11_ctrl_op_fcn;
  reg  T_38110_11_ctrl_fcn_dw;
  reg  T_38110_11_ctrl_rf_wen;
  reg [2:0] T_38110_11_ctrl_csr_cmd;
  reg  T_38110_11_ctrl_is_load;
  reg  T_38110_11_ctrl_is_sta;
  reg  T_38110_11_ctrl_is_std;
  reg [1:0] T_38110_11_wakeup_delay;
  reg  T_38110_11_allocate_brtag;
  reg  T_38110_11_is_br_or_jmp;
  reg  T_38110_11_is_jump;
  reg  T_38110_11_is_jal;
  reg  T_38110_11_is_ret;
  reg  T_38110_11_is_call;
  reg [7:0] T_38110_11_br_mask;
  reg [2:0] T_38110_11_br_tag;
  reg  T_38110_11_br_prediction_bpd_predict_val;
  reg  T_38110_11_br_prediction_bpd_predict_taken;
  reg  T_38110_11_br_prediction_btb_hit;
  reg  T_38110_11_br_prediction_btb_predicted;
  reg  T_38110_11_br_prediction_is_br_or_jalr;
  reg  T_38110_11_stat_brjmp_mispredicted;
  reg  T_38110_11_stat_btb_made_pred;
  reg  T_38110_11_stat_btb_mispredicted;
  reg  T_38110_11_stat_bpd_made_pred;
  reg  T_38110_11_stat_bpd_mispredicted;
  reg [2:0] T_38110_11_fetch_pc_lob;
  reg [19:0] T_38110_11_imm_packed;
  reg [11:0] T_38110_11_csr_addr;
  reg [5:0] T_38110_11_rob_idx;
  reg [3:0] T_38110_11_ldq_idx;
  reg [3:0] T_38110_11_stq_idx;
  reg [4:0] T_38110_11_brob_idx;
  reg [6:0] T_38110_11_pdst;
  reg [6:0] T_38110_11_pop1;
  reg [6:0] T_38110_11_pop2;
  reg [6:0] T_38110_11_pop3;
  reg  T_38110_11_prs1_busy;
  reg  T_38110_11_prs2_busy;
  reg  T_38110_11_prs3_busy;
  reg [6:0] T_38110_11_stale_pdst;
  reg  T_38110_11_exception;
  reg [63:0] T_38110_11_exc_cause;
  reg  T_38110_11_bypassable;
  reg [3:0] T_38110_11_mem_cmd;
  reg [2:0] T_38110_11_mem_typ;
  reg  T_38110_11_is_fence;
  reg  T_38110_11_is_fencei;
  reg  T_38110_11_is_store;
  reg  T_38110_11_is_amo;
  reg  T_38110_11_is_load;
  reg  T_38110_11_is_unique;
  reg  T_38110_11_flush_on_commit;
  reg [5:0] T_38110_11_ldst;
  reg [5:0] T_38110_11_lrs1;
  reg [5:0] T_38110_11_lrs2;
  reg [5:0] T_38110_11_lrs3;
  reg  T_38110_11_ldst_val;
  reg [1:0] T_38110_11_dst_rtype;
  reg [1:0] T_38110_11_lrs1_rtype;
  reg [1:0] T_38110_11_lrs2_rtype;
  reg  T_38110_11_frs3_en;
  reg  T_38110_11_fp_val;
  reg  T_38110_11_fp_single;
  reg  T_38110_11_xcpt_if;
  reg  T_38110_11_replay_if;
  reg [63:0] T_38110_11_debug_wdata;
  reg [31:0] T_38110_11_debug_events_fetch_seq;
  reg  T_38110_12_valid;
  reg [1:0] T_38110_12_iw_state;
  reg [8:0] T_38110_12_uopc;
  reg [31:0] T_38110_12_inst;
  reg [39:0] T_38110_12_pc;
  reg [7:0] T_38110_12_fu_code;
  reg [3:0] T_38110_12_ctrl_br_type;
  reg [1:0] T_38110_12_ctrl_op1_sel;
  reg [2:0] T_38110_12_ctrl_op2_sel;
  reg [2:0] T_38110_12_ctrl_imm_sel;
  reg [3:0] T_38110_12_ctrl_op_fcn;
  reg  T_38110_12_ctrl_fcn_dw;
  reg  T_38110_12_ctrl_rf_wen;
  reg [2:0] T_38110_12_ctrl_csr_cmd;
  reg  T_38110_12_ctrl_is_load;
  reg  T_38110_12_ctrl_is_sta;
  reg  T_38110_12_ctrl_is_std;
  reg [1:0] T_38110_12_wakeup_delay;
  reg  T_38110_12_allocate_brtag;
  reg  T_38110_12_is_br_or_jmp;
  reg  T_38110_12_is_jump;
  reg  T_38110_12_is_jal;
  reg  T_38110_12_is_ret;
  reg  T_38110_12_is_call;
  reg [7:0] T_38110_12_br_mask;
  reg [2:0] T_38110_12_br_tag;
  reg  T_38110_12_br_prediction_bpd_predict_val;
  reg  T_38110_12_br_prediction_bpd_predict_taken;
  reg  T_38110_12_br_prediction_btb_hit;
  reg  T_38110_12_br_prediction_btb_predicted;
  reg  T_38110_12_br_prediction_is_br_or_jalr;
  reg  T_38110_12_stat_brjmp_mispredicted;
  reg  T_38110_12_stat_btb_made_pred;
  reg  T_38110_12_stat_btb_mispredicted;
  reg  T_38110_12_stat_bpd_made_pred;
  reg  T_38110_12_stat_bpd_mispredicted;
  reg [2:0] T_38110_12_fetch_pc_lob;
  reg [19:0] T_38110_12_imm_packed;
  reg [11:0] T_38110_12_csr_addr;
  reg [5:0] T_38110_12_rob_idx;
  reg [3:0] T_38110_12_ldq_idx;
  reg [3:0] T_38110_12_stq_idx;
  reg [4:0] T_38110_12_brob_idx;
  reg [6:0] T_38110_12_pdst;
  reg [6:0] T_38110_12_pop1;
  reg [6:0] T_38110_12_pop2;
  reg [6:0] T_38110_12_pop3;
  reg  T_38110_12_prs1_busy;
  reg  T_38110_12_prs2_busy;
  reg  T_38110_12_prs3_busy;
  reg [6:0] T_38110_12_stale_pdst;
  reg  T_38110_12_exception;
  reg [63:0] T_38110_12_exc_cause;
  reg  T_38110_12_bypassable;
  reg [3:0] T_38110_12_mem_cmd;
  reg [2:0] T_38110_12_mem_typ;
  reg  T_38110_12_is_fence;
  reg  T_38110_12_is_fencei;
  reg  T_38110_12_is_store;
  reg  T_38110_12_is_amo;
  reg  T_38110_12_is_load;
  reg  T_38110_12_is_unique;
  reg  T_38110_12_flush_on_commit;
  reg [5:0] T_38110_12_ldst;
  reg [5:0] T_38110_12_lrs1;
  reg [5:0] T_38110_12_lrs2;
  reg [5:0] T_38110_12_lrs3;
  reg  T_38110_12_ldst_val;
  reg [1:0] T_38110_12_dst_rtype;
  reg [1:0] T_38110_12_lrs1_rtype;
  reg [1:0] T_38110_12_lrs2_rtype;
  reg  T_38110_12_frs3_en;
  reg  T_38110_12_fp_val;
  reg  T_38110_12_fp_single;
  reg  T_38110_12_xcpt_if;
  reg  T_38110_12_replay_if;
  reg [63:0] T_38110_12_debug_wdata;
  reg [31:0] T_38110_12_debug_events_fetch_seq;
  reg  T_38110_13_valid;
  reg [1:0] T_38110_13_iw_state;
  reg [8:0] T_38110_13_uopc;
  reg [31:0] T_38110_13_inst;
  reg [39:0] T_38110_13_pc;
  reg [7:0] T_38110_13_fu_code;
  reg [3:0] T_38110_13_ctrl_br_type;
  reg [1:0] T_38110_13_ctrl_op1_sel;
  reg [2:0] T_38110_13_ctrl_op2_sel;
  reg [2:0] T_38110_13_ctrl_imm_sel;
  reg [3:0] T_38110_13_ctrl_op_fcn;
  reg  T_38110_13_ctrl_fcn_dw;
  reg  T_38110_13_ctrl_rf_wen;
  reg [2:0] T_38110_13_ctrl_csr_cmd;
  reg  T_38110_13_ctrl_is_load;
  reg  T_38110_13_ctrl_is_sta;
  reg  T_38110_13_ctrl_is_std;
  reg [1:0] T_38110_13_wakeup_delay;
  reg  T_38110_13_allocate_brtag;
  reg  T_38110_13_is_br_or_jmp;
  reg  T_38110_13_is_jump;
  reg  T_38110_13_is_jal;
  reg  T_38110_13_is_ret;
  reg  T_38110_13_is_call;
  reg [7:0] T_38110_13_br_mask;
  reg [2:0] T_38110_13_br_tag;
  reg  T_38110_13_br_prediction_bpd_predict_val;
  reg  T_38110_13_br_prediction_bpd_predict_taken;
  reg  T_38110_13_br_prediction_btb_hit;
  reg  T_38110_13_br_prediction_btb_predicted;
  reg  T_38110_13_br_prediction_is_br_or_jalr;
  reg  T_38110_13_stat_brjmp_mispredicted;
  reg  T_38110_13_stat_btb_made_pred;
  reg  T_38110_13_stat_btb_mispredicted;
  reg  T_38110_13_stat_bpd_made_pred;
  reg  T_38110_13_stat_bpd_mispredicted;
  reg [2:0] T_38110_13_fetch_pc_lob;
  reg [19:0] T_38110_13_imm_packed;
  reg [11:0] T_38110_13_csr_addr;
  reg [5:0] T_38110_13_rob_idx;
  reg [3:0] T_38110_13_ldq_idx;
  reg [3:0] T_38110_13_stq_idx;
  reg [4:0] T_38110_13_brob_idx;
  reg [6:0] T_38110_13_pdst;
  reg [6:0] T_38110_13_pop1;
  reg [6:0] T_38110_13_pop2;
  reg [6:0] T_38110_13_pop3;
  reg  T_38110_13_prs1_busy;
  reg  T_38110_13_prs2_busy;
  reg  T_38110_13_prs3_busy;
  reg [6:0] T_38110_13_stale_pdst;
  reg  T_38110_13_exception;
  reg [63:0] T_38110_13_exc_cause;
  reg  T_38110_13_bypassable;
  reg [3:0] T_38110_13_mem_cmd;
  reg [2:0] T_38110_13_mem_typ;
  reg  T_38110_13_is_fence;
  reg  T_38110_13_is_fencei;
  reg  T_38110_13_is_store;
  reg  T_38110_13_is_amo;
  reg  T_38110_13_is_load;
  reg  T_38110_13_is_unique;
  reg  T_38110_13_flush_on_commit;
  reg [5:0] T_38110_13_ldst;
  reg [5:0] T_38110_13_lrs1;
  reg [5:0] T_38110_13_lrs2;
  reg [5:0] T_38110_13_lrs3;
  reg  T_38110_13_ldst_val;
  reg [1:0] T_38110_13_dst_rtype;
  reg [1:0] T_38110_13_lrs1_rtype;
  reg [1:0] T_38110_13_lrs2_rtype;
  reg  T_38110_13_frs3_en;
  reg  T_38110_13_fp_val;
  reg  T_38110_13_fp_single;
  reg  T_38110_13_xcpt_if;
  reg  T_38110_13_replay_if;
  reg [63:0] T_38110_13_debug_wdata;
  reg [31:0] T_38110_13_debug_events_fetch_seq;
  reg  T_38110_14_valid;
  reg [1:0] T_38110_14_iw_state;
  reg [8:0] T_38110_14_uopc;
  reg [31:0] T_38110_14_inst;
  reg [39:0] T_38110_14_pc;
  reg [7:0] T_38110_14_fu_code;
  reg [3:0] T_38110_14_ctrl_br_type;
  reg [1:0] T_38110_14_ctrl_op1_sel;
  reg [2:0] T_38110_14_ctrl_op2_sel;
  reg [2:0] T_38110_14_ctrl_imm_sel;
  reg [3:0] T_38110_14_ctrl_op_fcn;
  reg  T_38110_14_ctrl_fcn_dw;
  reg  T_38110_14_ctrl_rf_wen;
  reg [2:0] T_38110_14_ctrl_csr_cmd;
  reg  T_38110_14_ctrl_is_load;
  reg  T_38110_14_ctrl_is_sta;
  reg  T_38110_14_ctrl_is_std;
  reg [1:0] T_38110_14_wakeup_delay;
  reg  T_38110_14_allocate_brtag;
  reg  T_38110_14_is_br_or_jmp;
  reg  T_38110_14_is_jump;
  reg  T_38110_14_is_jal;
  reg  T_38110_14_is_ret;
  reg  T_38110_14_is_call;
  reg [7:0] T_38110_14_br_mask;
  reg [2:0] T_38110_14_br_tag;
  reg  T_38110_14_br_prediction_bpd_predict_val;
  reg  T_38110_14_br_prediction_bpd_predict_taken;
  reg  T_38110_14_br_prediction_btb_hit;
  reg  T_38110_14_br_prediction_btb_predicted;
  reg  T_38110_14_br_prediction_is_br_or_jalr;
  reg  T_38110_14_stat_brjmp_mispredicted;
  reg  T_38110_14_stat_btb_made_pred;
  reg  T_38110_14_stat_btb_mispredicted;
  reg  T_38110_14_stat_bpd_made_pred;
  reg  T_38110_14_stat_bpd_mispredicted;
  reg [2:0] T_38110_14_fetch_pc_lob;
  reg [19:0] T_38110_14_imm_packed;
  reg [11:0] T_38110_14_csr_addr;
  reg [5:0] T_38110_14_rob_idx;
  reg [3:0] T_38110_14_ldq_idx;
  reg [3:0] T_38110_14_stq_idx;
  reg [4:0] T_38110_14_brob_idx;
  reg [6:0] T_38110_14_pdst;
  reg [6:0] T_38110_14_pop1;
  reg [6:0] T_38110_14_pop2;
  reg [6:0] T_38110_14_pop3;
  reg  T_38110_14_prs1_busy;
  reg  T_38110_14_prs2_busy;
  reg  T_38110_14_prs3_busy;
  reg [6:0] T_38110_14_stale_pdst;
  reg  T_38110_14_exception;
  reg [63:0] T_38110_14_exc_cause;
  reg  T_38110_14_bypassable;
  reg [3:0] T_38110_14_mem_cmd;
  reg [2:0] T_38110_14_mem_typ;
  reg  T_38110_14_is_fence;
  reg  T_38110_14_is_fencei;
  reg  T_38110_14_is_store;
  reg  T_38110_14_is_amo;
  reg  T_38110_14_is_load;
  reg  T_38110_14_is_unique;
  reg  T_38110_14_flush_on_commit;
  reg [5:0] T_38110_14_ldst;
  reg [5:0] T_38110_14_lrs1;
  reg [5:0] T_38110_14_lrs2;
  reg [5:0] T_38110_14_lrs3;
  reg  T_38110_14_ldst_val;
  reg [1:0] T_38110_14_dst_rtype;
  reg [1:0] T_38110_14_lrs1_rtype;
  reg [1:0] T_38110_14_lrs2_rtype;
  reg  T_38110_14_frs3_en;
  reg  T_38110_14_fp_val;
  reg  T_38110_14_fp_single;
  reg  T_38110_14_xcpt_if;
  reg  T_38110_14_replay_if;
  reg [63:0] T_38110_14_debug_wdata;
  reg [31:0] T_38110_14_debug_events_fetch_seq;
  reg  T_38110_15_valid;
  reg [1:0] T_38110_15_iw_state;
  reg [8:0] T_38110_15_uopc;
  reg [31:0] T_38110_15_inst;
  reg [39:0] T_38110_15_pc;
  reg [7:0] T_38110_15_fu_code;
  reg [3:0] T_38110_15_ctrl_br_type;
  reg [1:0] T_38110_15_ctrl_op1_sel;
  reg [2:0] T_38110_15_ctrl_op2_sel;
  reg [2:0] T_38110_15_ctrl_imm_sel;
  reg [3:0] T_38110_15_ctrl_op_fcn;
  reg  T_38110_15_ctrl_fcn_dw;
  reg  T_38110_15_ctrl_rf_wen;
  reg [2:0] T_38110_15_ctrl_csr_cmd;
  reg  T_38110_15_ctrl_is_load;
  reg  T_38110_15_ctrl_is_sta;
  reg  T_38110_15_ctrl_is_std;
  reg [1:0] T_38110_15_wakeup_delay;
  reg  T_38110_15_allocate_brtag;
  reg  T_38110_15_is_br_or_jmp;
  reg  T_38110_15_is_jump;
  reg  T_38110_15_is_jal;
  reg  T_38110_15_is_ret;
  reg  T_38110_15_is_call;
  reg [7:0] T_38110_15_br_mask;
  reg [2:0] T_38110_15_br_tag;
  reg  T_38110_15_br_prediction_bpd_predict_val;
  reg  T_38110_15_br_prediction_bpd_predict_taken;
  reg  T_38110_15_br_prediction_btb_hit;
  reg  T_38110_15_br_prediction_btb_predicted;
  reg  T_38110_15_br_prediction_is_br_or_jalr;
  reg  T_38110_15_stat_brjmp_mispredicted;
  reg  T_38110_15_stat_btb_made_pred;
  reg  T_38110_15_stat_btb_mispredicted;
  reg  T_38110_15_stat_bpd_made_pred;
  reg  T_38110_15_stat_bpd_mispredicted;
  reg [2:0] T_38110_15_fetch_pc_lob;
  reg [19:0] T_38110_15_imm_packed;
  reg [11:0] T_38110_15_csr_addr;
  reg [5:0] T_38110_15_rob_idx;
  reg [3:0] T_38110_15_ldq_idx;
  reg [3:0] T_38110_15_stq_idx;
  reg [4:0] T_38110_15_brob_idx;
  reg [6:0] T_38110_15_pdst;
  reg [6:0] T_38110_15_pop1;
  reg [6:0] T_38110_15_pop2;
  reg [6:0] T_38110_15_pop3;
  reg  T_38110_15_prs1_busy;
  reg  T_38110_15_prs2_busy;
  reg  T_38110_15_prs3_busy;
  reg [6:0] T_38110_15_stale_pdst;
  reg  T_38110_15_exception;
  reg [63:0] T_38110_15_exc_cause;
  reg  T_38110_15_bypassable;
  reg [3:0] T_38110_15_mem_cmd;
  reg [2:0] T_38110_15_mem_typ;
  reg  T_38110_15_is_fence;
  reg  T_38110_15_is_fencei;
  reg  T_38110_15_is_store;
  reg  T_38110_15_is_amo;
  reg  T_38110_15_is_load;
  reg  T_38110_15_is_unique;
  reg  T_38110_15_flush_on_commit;
  reg [5:0] T_38110_15_ldst;
  reg [5:0] T_38110_15_lrs1;
  reg [5:0] T_38110_15_lrs2;
  reg [5:0] T_38110_15_lrs3;
  reg  T_38110_15_ldst_val;
  reg [1:0] T_38110_15_dst_rtype;
  reg [1:0] T_38110_15_lrs1_rtype;
  reg [1:0] T_38110_15_lrs2_rtype;
  reg  T_38110_15_frs3_en;
  reg  T_38110_15_fp_val;
  reg  T_38110_15_fp_single;
  reg  T_38110_15_xcpt_if;
  reg  T_38110_15_replay_if;
  reg [63:0] T_38110_15_debug_wdata;
  reg [31:0] T_38110_15_debug_events_fetch_seq;
  reg  T_38110_16_valid;
  reg [1:0] T_38110_16_iw_state;
  reg [8:0] T_38110_16_uopc;
  reg [31:0] T_38110_16_inst;
  reg [39:0] T_38110_16_pc;
  reg [7:0] T_38110_16_fu_code;
  reg [3:0] T_38110_16_ctrl_br_type;
  reg [1:0] T_38110_16_ctrl_op1_sel;
  reg [2:0] T_38110_16_ctrl_op2_sel;
  reg [2:0] T_38110_16_ctrl_imm_sel;
  reg [3:0] T_38110_16_ctrl_op_fcn;
  reg  T_38110_16_ctrl_fcn_dw;
  reg  T_38110_16_ctrl_rf_wen;
  reg [2:0] T_38110_16_ctrl_csr_cmd;
  reg  T_38110_16_ctrl_is_load;
  reg  T_38110_16_ctrl_is_sta;
  reg  T_38110_16_ctrl_is_std;
  reg [1:0] T_38110_16_wakeup_delay;
  reg  T_38110_16_allocate_brtag;
  reg  T_38110_16_is_br_or_jmp;
  reg  T_38110_16_is_jump;
  reg  T_38110_16_is_jal;
  reg  T_38110_16_is_ret;
  reg  T_38110_16_is_call;
  reg [7:0] T_38110_16_br_mask;
  reg [2:0] T_38110_16_br_tag;
  reg  T_38110_16_br_prediction_bpd_predict_val;
  reg  T_38110_16_br_prediction_bpd_predict_taken;
  reg  T_38110_16_br_prediction_btb_hit;
  reg  T_38110_16_br_prediction_btb_predicted;
  reg  T_38110_16_br_prediction_is_br_or_jalr;
  reg  T_38110_16_stat_brjmp_mispredicted;
  reg  T_38110_16_stat_btb_made_pred;
  reg  T_38110_16_stat_btb_mispredicted;
  reg  T_38110_16_stat_bpd_made_pred;
  reg  T_38110_16_stat_bpd_mispredicted;
  reg [2:0] T_38110_16_fetch_pc_lob;
  reg [19:0] T_38110_16_imm_packed;
  reg [11:0] T_38110_16_csr_addr;
  reg [5:0] T_38110_16_rob_idx;
  reg [3:0] T_38110_16_ldq_idx;
  reg [3:0] T_38110_16_stq_idx;
  reg [4:0] T_38110_16_brob_idx;
  reg [6:0] T_38110_16_pdst;
  reg [6:0] T_38110_16_pop1;
  reg [6:0] T_38110_16_pop2;
  reg [6:0] T_38110_16_pop3;
  reg  T_38110_16_prs1_busy;
  reg  T_38110_16_prs2_busy;
  reg  T_38110_16_prs3_busy;
  reg [6:0] T_38110_16_stale_pdst;
  reg  T_38110_16_exception;
  reg [63:0] T_38110_16_exc_cause;
  reg  T_38110_16_bypassable;
  reg [3:0] T_38110_16_mem_cmd;
  reg [2:0] T_38110_16_mem_typ;
  reg  T_38110_16_is_fence;
  reg  T_38110_16_is_fencei;
  reg  T_38110_16_is_store;
  reg  T_38110_16_is_amo;
  reg  T_38110_16_is_load;
  reg  T_38110_16_is_unique;
  reg  T_38110_16_flush_on_commit;
  reg [5:0] T_38110_16_ldst;
  reg [5:0] T_38110_16_lrs1;
  reg [5:0] T_38110_16_lrs2;
  reg [5:0] T_38110_16_lrs3;
  reg  T_38110_16_ldst_val;
  reg [1:0] T_38110_16_dst_rtype;
  reg [1:0] T_38110_16_lrs1_rtype;
  reg [1:0] T_38110_16_lrs2_rtype;
  reg  T_38110_16_frs3_en;
  reg  T_38110_16_fp_val;
  reg  T_38110_16_fp_single;
  reg  T_38110_16_xcpt_if;
  reg  T_38110_16_replay_if;
  reg [63:0] T_38110_16_debug_wdata;
  reg [31:0] T_38110_16_debug_events_fetch_seq;
  reg  T_38110_17_valid;
  reg [1:0] T_38110_17_iw_state;
  reg [8:0] T_38110_17_uopc;
  reg [31:0] T_38110_17_inst;
  reg [39:0] T_38110_17_pc;
  reg [7:0] T_38110_17_fu_code;
  reg [3:0] T_38110_17_ctrl_br_type;
  reg [1:0] T_38110_17_ctrl_op1_sel;
  reg [2:0] T_38110_17_ctrl_op2_sel;
  reg [2:0] T_38110_17_ctrl_imm_sel;
  reg [3:0] T_38110_17_ctrl_op_fcn;
  reg  T_38110_17_ctrl_fcn_dw;
  reg  T_38110_17_ctrl_rf_wen;
  reg [2:0] T_38110_17_ctrl_csr_cmd;
  reg  T_38110_17_ctrl_is_load;
  reg  T_38110_17_ctrl_is_sta;
  reg  T_38110_17_ctrl_is_std;
  reg [1:0] T_38110_17_wakeup_delay;
  reg  T_38110_17_allocate_brtag;
  reg  T_38110_17_is_br_or_jmp;
  reg  T_38110_17_is_jump;
  reg  T_38110_17_is_jal;
  reg  T_38110_17_is_ret;
  reg  T_38110_17_is_call;
  reg [7:0] T_38110_17_br_mask;
  reg [2:0] T_38110_17_br_tag;
  reg  T_38110_17_br_prediction_bpd_predict_val;
  reg  T_38110_17_br_prediction_bpd_predict_taken;
  reg  T_38110_17_br_prediction_btb_hit;
  reg  T_38110_17_br_prediction_btb_predicted;
  reg  T_38110_17_br_prediction_is_br_or_jalr;
  reg  T_38110_17_stat_brjmp_mispredicted;
  reg  T_38110_17_stat_btb_made_pred;
  reg  T_38110_17_stat_btb_mispredicted;
  reg  T_38110_17_stat_bpd_made_pred;
  reg  T_38110_17_stat_bpd_mispredicted;
  reg [2:0] T_38110_17_fetch_pc_lob;
  reg [19:0] T_38110_17_imm_packed;
  reg [11:0] T_38110_17_csr_addr;
  reg [5:0] T_38110_17_rob_idx;
  reg [3:0] T_38110_17_ldq_idx;
  reg [3:0] T_38110_17_stq_idx;
  reg [4:0] T_38110_17_brob_idx;
  reg [6:0] T_38110_17_pdst;
  reg [6:0] T_38110_17_pop1;
  reg [6:0] T_38110_17_pop2;
  reg [6:0] T_38110_17_pop3;
  reg  T_38110_17_prs1_busy;
  reg  T_38110_17_prs2_busy;
  reg  T_38110_17_prs3_busy;
  reg [6:0] T_38110_17_stale_pdst;
  reg  T_38110_17_exception;
  reg [63:0] T_38110_17_exc_cause;
  reg  T_38110_17_bypassable;
  reg [3:0] T_38110_17_mem_cmd;
  reg [2:0] T_38110_17_mem_typ;
  reg  T_38110_17_is_fence;
  reg  T_38110_17_is_fencei;
  reg  T_38110_17_is_store;
  reg  T_38110_17_is_amo;
  reg  T_38110_17_is_load;
  reg  T_38110_17_is_unique;
  reg  T_38110_17_flush_on_commit;
  reg [5:0] T_38110_17_ldst;
  reg [5:0] T_38110_17_lrs1;
  reg [5:0] T_38110_17_lrs2;
  reg [5:0] T_38110_17_lrs3;
  reg  T_38110_17_ldst_val;
  reg [1:0] T_38110_17_dst_rtype;
  reg [1:0] T_38110_17_lrs1_rtype;
  reg [1:0] T_38110_17_lrs2_rtype;
  reg  T_38110_17_frs3_en;
  reg  T_38110_17_fp_val;
  reg  T_38110_17_fp_single;
  reg  T_38110_17_xcpt_if;
  reg  T_38110_17_replay_if;
  reg [63:0] T_38110_17_debug_wdata;
  reg [31:0] T_38110_17_debug_events_fetch_seq;
  reg  T_38110_18_valid;
  reg [1:0] T_38110_18_iw_state;
  reg [8:0] T_38110_18_uopc;
  reg [31:0] T_38110_18_inst;
  reg [39:0] T_38110_18_pc;
  reg [7:0] T_38110_18_fu_code;
  reg [3:0] T_38110_18_ctrl_br_type;
  reg [1:0] T_38110_18_ctrl_op1_sel;
  reg [2:0] T_38110_18_ctrl_op2_sel;
  reg [2:0] T_38110_18_ctrl_imm_sel;
  reg [3:0] T_38110_18_ctrl_op_fcn;
  reg  T_38110_18_ctrl_fcn_dw;
  reg  T_38110_18_ctrl_rf_wen;
  reg [2:0] T_38110_18_ctrl_csr_cmd;
  reg  T_38110_18_ctrl_is_load;
  reg  T_38110_18_ctrl_is_sta;
  reg  T_38110_18_ctrl_is_std;
  reg [1:0] T_38110_18_wakeup_delay;
  reg  T_38110_18_allocate_brtag;
  reg  T_38110_18_is_br_or_jmp;
  reg  T_38110_18_is_jump;
  reg  T_38110_18_is_jal;
  reg  T_38110_18_is_ret;
  reg  T_38110_18_is_call;
  reg [7:0] T_38110_18_br_mask;
  reg [2:0] T_38110_18_br_tag;
  reg  T_38110_18_br_prediction_bpd_predict_val;
  reg  T_38110_18_br_prediction_bpd_predict_taken;
  reg  T_38110_18_br_prediction_btb_hit;
  reg  T_38110_18_br_prediction_btb_predicted;
  reg  T_38110_18_br_prediction_is_br_or_jalr;
  reg  T_38110_18_stat_brjmp_mispredicted;
  reg  T_38110_18_stat_btb_made_pred;
  reg  T_38110_18_stat_btb_mispredicted;
  reg  T_38110_18_stat_bpd_made_pred;
  reg  T_38110_18_stat_bpd_mispredicted;
  reg [2:0] T_38110_18_fetch_pc_lob;
  reg [19:0] T_38110_18_imm_packed;
  reg [11:0] T_38110_18_csr_addr;
  reg [5:0] T_38110_18_rob_idx;
  reg [3:0] T_38110_18_ldq_idx;
  reg [3:0] T_38110_18_stq_idx;
  reg [4:0] T_38110_18_brob_idx;
  reg [6:0] T_38110_18_pdst;
  reg [6:0] T_38110_18_pop1;
  reg [6:0] T_38110_18_pop2;
  reg [6:0] T_38110_18_pop3;
  reg  T_38110_18_prs1_busy;
  reg  T_38110_18_prs2_busy;
  reg  T_38110_18_prs3_busy;
  reg [6:0] T_38110_18_stale_pdst;
  reg  T_38110_18_exception;
  reg [63:0] T_38110_18_exc_cause;
  reg  T_38110_18_bypassable;
  reg [3:0] T_38110_18_mem_cmd;
  reg [2:0] T_38110_18_mem_typ;
  reg  T_38110_18_is_fence;
  reg  T_38110_18_is_fencei;
  reg  T_38110_18_is_store;
  reg  T_38110_18_is_amo;
  reg  T_38110_18_is_load;
  reg  T_38110_18_is_unique;
  reg  T_38110_18_flush_on_commit;
  reg [5:0] T_38110_18_ldst;
  reg [5:0] T_38110_18_lrs1;
  reg [5:0] T_38110_18_lrs2;
  reg [5:0] T_38110_18_lrs3;
  reg  T_38110_18_ldst_val;
  reg [1:0] T_38110_18_dst_rtype;
  reg [1:0] T_38110_18_lrs1_rtype;
  reg [1:0] T_38110_18_lrs2_rtype;
  reg  T_38110_18_frs3_en;
  reg  T_38110_18_fp_val;
  reg  T_38110_18_fp_single;
  reg  T_38110_18_xcpt_if;
  reg  T_38110_18_replay_if;
  reg [63:0] T_38110_18_debug_wdata;
  reg [31:0] T_38110_18_debug_events_fetch_seq;
  reg  T_38110_19_valid;
  reg [1:0] T_38110_19_iw_state;
  reg [8:0] T_38110_19_uopc;
  reg [31:0] T_38110_19_inst;
  reg [39:0] T_38110_19_pc;
  reg [7:0] T_38110_19_fu_code;
  reg [3:0] T_38110_19_ctrl_br_type;
  reg [1:0] T_38110_19_ctrl_op1_sel;
  reg [2:0] T_38110_19_ctrl_op2_sel;
  reg [2:0] T_38110_19_ctrl_imm_sel;
  reg [3:0] T_38110_19_ctrl_op_fcn;
  reg  T_38110_19_ctrl_fcn_dw;
  reg  T_38110_19_ctrl_rf_wen;
  reg [2:0] T_38110_19_ctrl_csr_cmd;
  reg  T_38110_19_ctrl_is_load;
  reg  T_38110_19_ctrl_is_sta;
  reg  T_38110_19_ctrl_is_std;
  reg [1:0] T_38110_19_wakeup_delay;
  reg  T_38110_19_allocate_brtag;
  reg  T_38110_19_is_br_or_jmp;
  reg  T_38110_19_is_jump;
  reg  T_38110_19_is_jal;
  reg  T_38110_19_is_ret;
  reg  T_38110_19_is_call;
  reg [7:0] T_38110_19_br_mask;
  reg [2:0] T_38110_19_br_tag;
  reg  T_38110_19_br_prediction_bpd_predict_val;
  reg  T_38110_19_br_prediction_bpd_predict_taken;
  reg  T_38110_19_br_prediction_btb_hit;
  reg  T_38110_19_br_prediction_btb_predicted;
  reg  T_38110_19_br_prediction_is_br_or_jalr;
  reg  T_38110_19_stat_brjmp_mispredicted;
  reg  T_38110_19_stat_btb_made_pred;
  reg  T_38110_19_stat_btb_mispredicted;
  reg  T_38110_19_stat_bpd_made_pred;
  reg  T_38110_19_stat_bpd_mispredicted;
  reg [2:0] T_38110_19_fetch_pc_lob;
  reg [19:0] T_38110_19_imm_packed;
  reg [11:0] T_38110_19_csr_addr;
  reg [5:0] T_38110_19_rob_idx;
  reg [3:0] T_38110_19_ldq_idx;
  reg [3:0] T_38110_19_stq_idx;
  reg [4:0] T_38110_19_brob_idx;
  reg [6:0] T_38110_19_pdst;
  reg [6:0] T_38110_19_pop1;
  reg [6:0] T_38110_19_pop2;
  reg [6:0] T_38110_19_pop3;
  reg  T_38110_19_prs1_busy;
  reg  T_38110_19_prs2_busy;
  reg  T_38110_19_prs3_busy;
  reg [6:0] T_38110_19_stale_pdst;
  reg  T_38110_19_exception;
  reg [63:0] T_38110_19_exc_cause;
  reg  T_38110_19_bypassable;
  reg [3:0] T_38110_19_mem_cmd;
  reg [2:0] T_38110_19_mem_typ;
  reg  T_38110_19_is_fence;
  reg  T_38110_19_is_fencei;
  reg  T_38110_19_is_store;
  reg  T_38110_19_is_amo;
  reg  T_38110_19_is_load;
  reg  T_38110_19_is_unique;
  reg  T_38110_19_flush_on_commit;
  reg [5:0] T_38110_19_ldst;
  reg [5:0] T_38110_19_lrs1;
  reg [5:0] T_38110_19_lrs2;
  reg [5:0] T_38110_19_lrs3;
  reg  T_38110_19_ldst_val;
  reg [1:0] T_38110_19_dst_rtype;
  reg [1:0] T_38110_19_lrs1_rtype;
  reg [1:0] T_38110_19_lrs2_rtype;
  reg  T_38110_19_frs3_en;
  reg  T_38110_19_fp_val;
  reg  T_38110_19_fp_single;
  reg  T_38110_19_xcpt_if;
  reg  T_38110_19_replay_if;
  reg [63:0] T_38110_19_debug_wdata;
  reg [31:0] T_38110_19_debug_events_fetch_seq;
  reg  T_38110_20_valid;
  reg [1:0] T_38110_20_iw_state;
  reg [8:0] T_38110_20_uopc;
  reg [31:0] T_38110_20_inst;
  reg [39:0] T_38110_20_pc;
  reg [7:0] T_38110_20_fu_code;
  reg [3:0] T_38110_20_ctrl_br_type;
  reg [1:0] T_38110_20_ctrl_op1_sel;
  reg [2:0] T_38110_20_ctrl_op2_sel;
  reg [2:0] T_38110_20_ctrl_imm_sel;
  reg [3:0] T_38110_20_ctrl_op_fcn;
  reg  T_38110_20_ctrl_fcn_dw;
  reg  T_38110_20_ctrl_rf_wen;
  reg [2:0] T_38110_20_ctrl_csr_cmd;
  reg  T_38110_20_ctrl_is_load;
  reg  T_38110_20_ctrl_is_sta;
  reg  T_38110_20_ctrl_is_std;
  reg [1:0] T_38110_20_wakeup_delay;
  reg  T_38110_20_allocate_brtag;
  reg  T_38110_20_is_br_or_jmp;
  reg  T_38110_20_is_jump;
  reg  T_38110_20_is_jal;
  reg  T_38110_20_is_ret;
  reg  T_38110_20_is_call;
  reg [7:0] T_38110_20_br_mask;
  reg [2:0] T_38110_20_br_tag;
  reg  T_38110_20_br_prediction_bpd_predict_val;
  reg  T_38110_20_br_prediction_bpd_predict_taken;
  reg  T_38110_20_br_prediction_btb_hit;
  reg  T_38110_20_br_prediction_btb_predicted;
  reg  T_38110_20_br_prediction_is_br_or_jalr;
  reg  T_38110_20_stat_brjmp_mispredicted;
  reg  T_38110_20_stat_btb_made_pred;
  reg  T_38110_20_stat_btb_mispredicted;
  reg  T_38110_20_stat_bpd_made_pred;
  reg  T_38110_20_stat_bpd_mispredicted;
  reg [2:0] T_38110_20_fetch_pc_lob;
  reg [19:0] T_38110_20_imm_packed;
  reg [11:0] T_38110_20_csr_addr;
  reg [5:0] T_38110_20_rob_idx;
  reg [3:0] T_38110_20_ldq_idx;
  reg [3:0] T_38110_20_stq_idx;
  reg [4:0] T_38110_20_brob_idx;
  reg [6:0] T_38110_20_pdst;
  reg [6:0] T_38110_20_pop1;
  reg [6:0] T_38110_20_pop2;
  reg [6:0] T_38110_20_pop3;
  reg  T_38110_20_prs1_busy;
  reg  T_38110_20_prs2_busy;
  reg  T_38110_20_prs3_busy;
  reg [6:0] T_38110_20_stale_pdst;
  reg  T_38110_20_exception;
  reg [63:0] T_38110_20_exc_cause;
  reg  T_38110_20_bypassable;
  reg [3:0] T_38110_20_mem_cmd;
  reg [2:0] T_38110_20_mem_typ;
  reg  T_38110_20_is_fence;
  reg  T_38110_20_is_fencei;
  reg  T_38110_20_is_store;
  reg  T_38110_20_is_amo;
  reg  T_38110_20_is_load;
  reg  T_38110_20_is_unique;
  reg  T_38110_20_flush_on_commit;
  reg [5:0] T_38110_20_ldst;
  reg [5:0] T_38110_20_lrs1;
  reg [5:0] T_38110_20_lrs2;
  reg [5:0] T_38110_20_lrs3;
  reg  T_38110_20_ldst_val;
  reg [1:0] T_38110_20_dst_rtype;
  reg [1:0] T_38110_20_lrs1_rtype;
  reg [1:0] T_38110_20_lrs2_rtype;
  reg  T_38110_20_frs3_en;
  reg  T_38110_20_fp_val;
  reg  T_38110_20_fp_single;
  reg  T_38110_20_xcpt_if;
  reg  T_38110_20_replay_if;
  reg [63:0] T_38110_20_debug_wdata;
  reg [31:0] T_38110_20_debug_events_fetch_seq;
  reg  T_38110_21_valid;
  reg [1:0] T_38110_21_iw_state;
  reg [8:0] T_38110_21_uopc;
  reg [31:0] T_38110_21_inst;
  reg [39:0] T_38110_21_pc;
  reg [7:0] T_38110_21_fu_code;
  reg [3:0] T_38110_21_ctrl_br_type;
  reg [1:0] T_38110_21_ctrl_op1_sel;
  reg [2:0] T_38110_21_ctrl_op2_sel;
  reg [2:0] T_38110_21_ctrl_imm_sel;
  reg [3:0] T_38110_21_ctrl_op_fcn;
  reg  T_38110_21_ctrl_fcn_dw;
  reg  T_38110_21_ctrl_rf_wen;
  reg [2:0] T_38110_21_ctrl_csr_cmd;
  reg  T_38110_21_ctrl_is_load;
  reg  T_38110_21_ctrl_is_sta;
  reg  T_38110_21_ctrl_is_std;
  reg [1:0] T_38110_21_wakeup_delay;
  reg  T_38110_21_allocate_brtag;
  reg  T_38110_21_is_br_or_jmp;
  reg  T_38110_21_is_jump;
  reg  T_38110_21_is_jal;
  reg  T_38110_21_is_ret;
  reg  T_38110_21_is_call;
  reg [7:0] T_38110_21_br_mask;
  reg [2:0] T_38110_21_br_tag;
  reg  T_38110_21_br_prediction_bpd_predict_val;
  reg  T_38110_21_br_prediction_bpd_predict_taken;
  reg  T_38110_21_br_prediction_btb_hit;
  reg  T_38110_21_br_prediction_btb_predicted;
  reg  T_38110_21_br_prediction_is_br_or_jalr;
  reg  T_38110_21_stat_brjmp_mispredicted;
  reg  T_38110_21_stat_btb_made_pred;
  reg  T_38110_21_stat_btb_mispredicted;
  reg  T_38110_21_stat_bpd_made_pred;
  reg  T_38110_21_stat_bpd_mispredicted;
  reg [2:0] T_38110_21_fetch_pc_lob;
  reg [19:0] T_38110_21_imm_packed;
  reg [11:0] T_38110_21_csr_addr;
  reg [5:0] T_38110_21_rob_idx;
  reg [3:0] T_38110_21_ldq_idx;
  reg [3:0] T_38110_21_stq_idx;
  reg [4:0] T_38110_21_brob_idx;
  reg [6:0] T_38110_21_pdst;
  reg [6:0] T_38110_21_pop1;
  reg [6:0] T_38110_21_pop2;
  reg [6:0] T_38110_21_pop3;
  reg  T_38110_21_prs1_busy;
  reg  T_38110_21_prs2_busy;
  reg  T_38110_21_prs3_busy;
  reg [6:0] T_38110_21_stale_pdst;
  reg  T_38110_21_exception;
  reg [63:0] T_38110_21_exc_cause;
  reg  T_38110_21_bypassable;
  reg [3:0] T_38110_21_mem_cmd;
  reg [2:0] T_38110_21_mem_typ;
  reg  T_38110_21_is_fence;
  reg  T_38110_21_is_fencei;
  reg  T_38110_21_is_store;
  reg  T_38110_21_is_amo;
  reg  T_38110_21_is_load;
  reg  T_38110_21_is_unique;
  reg  T_38110_21_flush_on_commit;
  reg [5:0] T_38110_21_ldst;
  reg [5:0] T_38110_21_lrs1;
  reg [5:0] T_38110_21_lrs2;
  reg [5:0] T_38110_21_lrs3;
  reg  T_38110_21_ldst_val;
  reg [1:0] T_38110_21_dst_rtype;
  reg [1:0] T_38110_21_lrs1_rtype;
  reg [1:0] T_38110_21_lrs2_rtype;
  reg  T_38110_21_frs3_en;
  reg  T_38110_21_fp_val;
  reg  T_38110_21_fp_single;
  reg  T_38110_21_xcpt_if;
  reg  T_38110_21_replay_if;
  reg [63:0] T_38110_21_debug_wdata;
  reg [31:0] T_38110_21_debug_events_fetch_seq;
  reg  T_38110_22_valid;
  reg [1:0] T_38110_22_iw_state;
  reg [8:0] T_38110_22_uopc;
  reg [31:0] T_38110_22_inst;
  reg [39:0] T_38110_22_pc;
  reg [7:0] T_38110_22_fu_code;
  reg [3:0] T_38110_22_ctrl_br_type;
  reg [1:0] T_38110_22_ctrl_op1_sel;
  reg [2:0] T_38110_22_ctrl_op2_sel;
  reg [2:0] T_38110_22_ctrl_imm_sel;
  reg [3:0] T_38110_22_ctrl_op_fcn;
  reg  T_38110_22_ctrl_fcn_dw;
  reg  T_38110_22_ctrl_rf_wen;
  reg [2:0] T_38110_22_ctrl_csr_cmd;
  reg  T_38110_22_ctrl_is_load;
  reg  T_38110_22_ctrl_is_sta;
  reg  T_38110_22_ctrl_is_std;
  reg [1:0] T_38110_22_wakeup_delay;
  reg  T_38110_22_allocate_brtag;
  reg  T_38110_22_is_br_or_jmp;
  reg  T_38110_22_is_jump;
  reg  T_38110_22_is_jal;
  reg  T_38110_22_is_ret;
  reg  T_38110_22_is_call;
  reg [7:0] T_38110_22_br_mask;
  reg [2:0] T_38110_22_br_tag;
  reg  T_38110_22_br_prediction_bpd_predict_val;
  reg  T_38110_22_br_prediction_bpd_predict_taken;
  reg  T_38110_22_br_prediction_btb_hit;
  reg  T_38110_22_br_prediction_btb_predicted;
  reg  T_38110_22_br_prediction_is_br_or_jalr;
  reg  T_38110_22_stat_brjmp_mispredicted;
  reg  T_38110_22_stat_btb_made_pred;
  reg  T_38110_22_stat_btb_mispredicted;
  reg  T_38110_22_stat_bpd_made_pred;
  reg  T_38110_22_stat_bpd_mispredicted;
  reg [2:0] T_38110_22_fetch_pc_lob;
  reg [19:0] T_38110_22_imm_packed;
  reg [11:0] T_38110_22_csr_addr;
  reg [5:0] T_38110_22_rob_idx;
  reg [3:0] T_38110_22_ldq_idx;
  reg [3:0] T_38110_22_stq_idx;
  reg [4:0] T_38110_22_brob_idx;
  reg [6:0] T_38110_22_pdst;
  reg [6:0] T_38110_22_pop1;
  reg [6:0] T_38110_22_pop2;
  reg [6:0] T_38110_22_pop3;
  reg  T_38110_22_prs1_busy;
  reg  T_38110_22_prs2_busy;
  reg  T_38110_22_prs3_busy;
  reg [6:0] T_38110_22_stale_pdst;
  reg  T_38110_22_exception;
  reg [63:0] T_38110_22_exc_cause;
  reg  T_38110_22_bypassable;
  reg [3:0] T_38110_22_mem_cmd;
  reg [2:0] T_38110_22_mem_typ;
  reg  T_38110_22_is_fence;
  reg  T_38110_22_is_fencei;
  reg  T_38110_22_is_store;
  reg  T_38110_22_is_amo;
  reg  T_38110_22_is_load;
  reg  T_38110_22_is_unique;
  reg  T_38110_22_flush_on_commit;
  reg [5:0] T_38110_22_ldst;
  reg [5:0] T_38110_22_lrs1;
  reg [5:0] T_38110_22_lrs2;
  reg [5:0] T_38110_22_lrs3;
  reg  T_38110_22_ldst_val;
  reg [1:0] T_38110_22_dst_rtype;
  reg [1:0] T_38110_22_lrs1_rtype;
  reg [1:0] T_38110_22_lrs2_rtype;
  reg  T_38110_22_frs3_en;
  reg  T_38110_22_fp_val;
  reg  T_38110_22_fp_single;
  reg  T_38110_22_xcpt_if;
  reg  T_38110_22_replay_if;
  reg [63:0] T_38110_22_debug_wdata;
  reg [31:0] T_38110_22_debug_events_fetch_seq;
  reg  T_38110_23_valid;
  reg [1:0] T_38110_23_iw_state;
  reg [8:0] T_38110_23_uopc;
  reg [31:0] T_38110_23_inst;
  reg [39:0] T_38110_23_pc;
  reg [7:0] T_38110_23_fu_code;
  reg [3:0] T_38110_23_ctrl_br_type;
  reg [1:0] T_38110_23_ctrl_op1_sel;
  reg [2:0] T_38110_23_ctrl_op2_sel;
  reg [2:0] T_38110_23_ctrl_imm_sel;
  reg [3:0] T_38110_23_ctrl_op_fcn;
  reg  T_38110_23_ctrl_fcn_dw;
  reg  T_38110_23_ctrl_rf_wen;
  reg [2:0] T_38110_23_ctrl_csr_cmd;
  reg  T_38110_23_ctrl_is_load;
  reg  T_38110_23_ctrl_is_sta;
  reg  T_38110_23_ctrl_is_std;
  reg [1:0] T_38110_23_wakeup_delay;
  reg  T_38110_23_allocate_brtag;
  reg  T_38110_23_is_br_or_jmp;
  reg  T_38110_23_is_jump;
  reg  T_38110_23_is_jal;
  reg  T_38110_23_is_ret;
  reg  T_38110_23_is_call;
  reg [7:0] T_38110_23_br_mask;
  reg [2:0] T_38110_23_br_tag;
  reg  T_38110_23_br_prediction_bpd_predict_val;
  reg  T_38110_23_br_prediction_bpd_predict_taken;
  reg  T_38110_23_br_prediction_btb_hit;
  reg  T_38110_23_br_prediction_btb_predicted;
  reg  T_38110_23_br_prediction_is_br_or_jalr;
  reg  T_38110_23_stat_brjmp_mispredicted;
  reg  T_38110_23_stat_btb_made_pred;
  reg  T_38110_23_stat_btb_mispredicted;
  reg  T_38110_23_stat_bpd_made_pred;
  reg  T_38110_23_stat_bpd_mispredicted;
  reg [2:0] T_38110_23_fetch_pc_lob;
  reg [19:0] T_38110_23_imm_packed;
  reg [11:0] T_38110_23_csr_addr;
  reg [5:0] T_38110_23_rob_idx;
  reg [3:0] T_38110_23_ldq_idx;
  reg [3:0] T_38110_23_stq_idx;
  reg [4:0] T_38110_23_brob_idx;
  reg [6:0] T_38110_23_pdst;
  reg [6:0] T_38110_23_pop1;
  reg [6:0] T_38110_23_pop2;
  reg [6:0] T_38110_23_pop3;
  reg  T_38110_23_prs1_busy;
  reg  T_38110_23_prs2_busy;
  reg  T_38110_23_prs3_busy;
  reg [6:0] T_38110_23_stale_pdst;
  reg  T_38110_23_exception;
  reg [63:0] T_38110_23_exc_cause;
  reg  T_38110_23_bypassable;
  reg [3:0] T_38110_23_mem_cmd;
  reg [2:0] T_38110_23_mem_typ;
  reg  T_38110_23_is_fence;
  reg  T_38110_23_is_fencei;
  reg  T_38110_23_is_store;
  reg  T_38110_23_is_amo;
  reg  T_38110_23_is_load;
  reg  T_38110_23_is_unique;
  reg  T_38110_23_flush_on_commit;
  reg [5:0] T_38110_23_ldst;
  reg [5:0] T_38110_23_lrs1;
  reg [5:0] T_38110_23_lrs2;
  reg [5:0] T_38110_23_lrs3;
  reg  T_38110_23_ldst_val;
  reg [1:0] T_38110_23_dst_rtype;
  reg [1:0] T_38110_23_lrs1_rtype;
  reg [1:0] T_38110_23_lrs2_rtype;
  reg  T_38110_23_frs3_en;
  reg  T_38110_23_fp_val;
  reg  T_38110_23_fp_single;
  reg  T_38110_23_xcpt_if;
  reg  T_38110_23_replay_if;
  reg [63:0] T_38110_23_debug_wdata;
  reg [31:0] T_38110_23_debug_events_fetch_seq;
  wire  _GEN_14176 = 5'h0 == rob_tail | T_35634_0; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14177 = 5'h1 == rob_tail | T_35634_1; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14178 = 5'h2 == rob_tail | T_35634_2; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14179 = 5'h3 == rob_tail | T_35634_3; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14180 = 5'h4 == rob_tail | T_35634_4; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14181 = 5'h5 == rob_tail | T_35634_5; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14182 = 5'h6 == rob_tail | T_35634_6; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14183 = 5'h7 == rob_tail | T_35634_7; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14184 = 5'h8 == rob_tail | T_35634_8; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14185 = 5'h9 == rob_tail | T_35634_9; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14186 = 5'ha == rob_tail | T_35634_10; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14187 = 5'hb == rob_tail | T_35634_11; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14188 = 5'hc == rob_tail | T_35634_12; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14189 = 5'hd == rob_tail | T_35634_13; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14190 = 5'he == rob_tail | T_35634_14; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14191 = 5'hf == rob_tail | T_35634_15; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14192 = 5'h10 == rob_tail | T_35634_16; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14193 = 5'h11 == rob_tail | T_35634_17; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14194 = 5'h12 == rob_tail | T_35634_18; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14195 = 5'h13 == rob_tail | T_35634_19; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14196 = 5'h14 == rob_tail | T_35634_20; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14197 = 5'h15 == rob_tail | T_35634_21; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14198 = 5'h16 == rob_tail | T_35634_22; // @[rob.scala 347:34 rob.scala 347:34]
  wire  _GEN_14199 = 5'h17 == rob_tail | T_35634_23; // @[rob.scala 347:34 rob.scala 347:34]
  wire [31:0] _GEN_14272 = 5'h0 == rob_tail ? io_dis_uops_1_inst : T_38110_0_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14273 = 5'h1 == rob_tail ? io_dis_uops_1_inst : T_38110_1_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14274 = 5'h2 == rob_tail ? io_dis_uops_1_inst : T_38110_2_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14275 = 5'h3 == rob_tail ? io_dis_uops_1_inst : T_38110_3_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14276 = 5'h4 == rob_tail ? io_dis_uops_1_inst : T_38110_4_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14277 = 5'h5 == rob_tail ? io_dis_uops_1_inst : T_38110_5_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14278 = 5'h6 == rob_tail ? io_dis_uops_1_inst : T_38110_6_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14279 = 5'h7 == rob_tail ? io_dis_uops_1_inst : T_38110_7_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14280 = 5'h8 == rob_tail ? io_dis_uops_1_inst : T_38110_8_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14281 = 5'h9 == rob_tail ? io_dis_uops_1_inst : T_38110_9_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14282 = 5'ha == rob_tail ? io_dis_uops_1_inst : T_38110_10_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14283 = 5'hb == rob_tail ? io_dis_uops_1_inst : T_38110_11_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14284 = 5'hc == rob_tail ? io_dis_uops_1_inst : T_38110_12_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14285 = 5'hd == rob_tail ? io_dis_uops_1_inst : T_38110_13_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14286 = 5'he == rob_tail ? io_dis_uops_1_inst : T_38110_14_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14287 = 5'hf == rob_tail ? io_dis_uops_1_inst : T_38110_15_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14288 = 5'h10 == rob_tail ? io_dis_uops_1_inst : T_38110_16_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14289 = 5'h11 == rob_tail ? io_dis_uops_1_inst : T_38110_17_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14290 = 5'h12 == rob_tail ? io_dis_uops_1_inst : T_38110_18_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14291 = 5'h13 == rob_tail ? io_dis_uops_1_inst : T_38110_19_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14292 = 5'h14 == rob_tail ? io_dis_uops_1_inst : T_38110_20_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14293 = 5'h15 == rob_tail ? io_dis_uops_1_inst : T_38110_21_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14294 = 5'h16 == rob_tail ? io_dis_uops_1_inst : T_38110_22_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire [31:0] _GEN_14295 = 5'h17 == rob_tail ? io_dis_uops_1_inst : T_38110_23_inst; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14944 = 5'h0 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_0_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14945 = 5'h1 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_1_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14946 = 5'h2 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_2_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14947 = 5'h3 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_3_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14948 = 5'h4 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_4_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14949 = 5'h5 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_5_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14950 = 5'h6 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_6_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14951 = 5'h7 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_7_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14952 = 5'h8 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_8_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14953 = 5'h9 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_9_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14954 = 5'ha == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_10_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14955 = 5'hb == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_11_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14956 = 5'hc == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_12_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14957 = 5'hd == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_13_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14958 = 5'he == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_14_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14959 = 5'hf == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_15_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14960 = 5'h10 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_16_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14961 = 5'h11 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_17_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14962 = 5'h12 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_18_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14963 = 5'h13 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_19_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14964 = 5'h14 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_20_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14965 = 5'h15 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_21_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14966 = 5'h16 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_22_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14967 = 5'h17 == rob_tail ? io_dis_uops_1_stat_brjmp_mispredicted : T_38110_23_stat_brjmp_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14968 = 5'h0 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_0_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14969 = 5'h1 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_1_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14970 = 5'h2 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_2_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14971 = 5'h3 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_3_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14972 = 5'h4 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_4_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14973 = 5'h5 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_5_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14974 = 5'h6 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_6_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14975 = 5'h7 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_7_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14976 = 5'h8 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_8_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14977 = 5'h9 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_9_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14978 = 5'ha == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_10_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14979 = 5'hb == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_11_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14980 = 5'hc == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_12_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14981 = 5'hd == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_13_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14982 = 5'he == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_14_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14983 = 5'hf == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_15_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14984 = 5'h10 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_16_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14985 = 5'h11 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_17_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14986 = 5'h12 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_18_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14987 = 5'h13 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_19_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14988 = 5'h14 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_20_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14989 = 5'h15 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_21_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14990 = 5'h16 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_22_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14991 = 5'h17 == rob_tail ? io_dis_uops_1_stat_btb_made_pred : T_38110_23_stat_btb_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14992 = 5'h0 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_0_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14993 = 5'h1 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_1_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14994 = 5'h2 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_2_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14995 = 5'h3 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_3_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14996 = 5'h4 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_4_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14997 = 5'h5 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_5_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14998 = 5'h6 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_6_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_14999 = 5'h7 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_7_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15000 = 5'h8 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_8_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15001 = 5'h9 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_9_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15002 = 5'ha == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_10_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15003 = 5'hb == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_11_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15004 = 5'hc == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_12_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15005 = 5'hd == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_13_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15006 = 5'he == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_14_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15007 = 5'hf == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_15_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15008 = 5'h10 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_16_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15009 = 5'h11 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_17_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15010 = 5'h12 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_18_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15011 = 5'h13 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_19_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15012 = 5'h14 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_20_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15013 = 5'h15 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_21_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15014 = 5'h16 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_22_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15015 = 5'h17 == rob_tail ? io_dis_uops_1_stat_btb_mispredicted : T_38110_23_stat_btb_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15016 = 5'h0 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_0_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15017 = 5'h1 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_1_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15018 = 5'h2 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_2_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15019 = 5'h3 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_3_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15020 = 5'h4 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_4_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15021 = 5'h5 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_5_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15022 = 5'h6 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_6_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15023 = 5'h7 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_7_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15024 = 5'h8 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_8_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15025 = 5'h9 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_9_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15026 = 5'ha == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_10_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15027 = 5'hb == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_11_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15028 = 5'hc == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_12_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15029 = 5'hd == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_13_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15030 = 5'he == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_14_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15031 = 5'hf == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_15_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15032 = 5'h10 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_16_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15033 = 5'h11 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_17_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15034 = 5'h12 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_18_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15035 = 5'h13 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_19_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15036 = 5'h14 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_20_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15037 = 5'h15 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_21_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15038 = 5'h16 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_22_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15039 = 5'h17 == rob_tail ? io_dis_uops_1_stat_bpd_made_pred : T_38110_23_stat_bpd_made_pred; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15040 = 5'h0 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_0_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15041 = 5'h1 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_1_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15042 = 5'h2 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_2_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15043 = 5'h3 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_3_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15044 = 5'h4 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_4_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15045 = 5'h5 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_5_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15046 = 5'h6 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_6_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15047 = 5'h7 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_7_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15048 = 5'h8 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_8_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15049 = 5'h9 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_9_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15050 = 5'ha == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_10_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15051 = 5'hb == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_11_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15052 = 5'hc == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_12_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15053 = 5'hd == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_13_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15054 = 5'he == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_14_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15055 = 5'hf == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_15_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15056 = 5'h10 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_16_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15057 = 5'h11 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_17_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15058 = 5'h12 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_18_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15059 = 5'h13 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_19_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15060 = 5'h14 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_20_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15061 = 5'h15 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_21_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15062 = 5'h16 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_22_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_15063 = 5'h17 == rob_tail ? io_dis_uops_1_stat_bpd_mispredicted : T_38110_23_stat_bpd_mispredicted; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16024 = 5'h0 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_0_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16025 = 5'h1 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_1_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16026 = 5'h2 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_2_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16027 = 5'h3 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_3_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16028 = 5'h4 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_4_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16029 = 5'h5 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_5_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16030 = 5'h6 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_6_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16031 = 5'h7 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_7_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16032 = 5'h8 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_8_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16033 = 5'h9 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_9_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16034 = 5'ha == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_10_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16035 = 5'hb == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_11_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16036 = 5'hc == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_12_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16037 = 5'hd == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_13_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16038 = 5'he == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_14_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16039 = 5'hf == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_15_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16040 = 5'h10 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_16_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16041 = 5'h11 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_17_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16042 = 5'h12 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_18_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16043 = 5'h13 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_19_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16044 = 5'h14 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_20_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16045 = 5'h15 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_21_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16046 = 5'h16 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_22_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire [63:0] _GEN_16047 = 5'h17 == rob_tail ? io_dis_uops_1_debug_wdata : T_38110_23_debug_wdata; // @[rob.scala 350:34 rob.scala 350:34]
  wire  _GEN_16072 = 5'h0 == rob_tail ? 1'h0 : _GEN_14944; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16073 = 5'h1 == rob_tail ? 1'h0 : _GEN_14945; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16074 = 5'h2 == rob_tail ? 1'h0 : _GEN_14946; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16075 = 5'h3 == rob_tail ? 1'h0 : _GEN_14947; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16076 = 5'h4 == rob_tail ? 1'h0 : _GEN_14948; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16077 = 5'h5 == rob_tail ? 1'h0 : _GEN_14949; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16078 = 5'h6 == rob_tail ? 1'h0 : _GEN_14950; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16079 = 5'h7 == rob_tail ? 1'h0 : _GEN_14951; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16080 = 5'h8 == rob_tail ? 1'h0 : _GEN_14952; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16081 = 5'h9 == rob_tail ? 1'h0 : _GEN_14953; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16082 = 5'ha == rob_tail ? 1'h0 : _GEN_14954; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16083 = 5'hb == rob_tail ? 1'h0 : _GEN_14955; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16084 = 5'hc == rob_tail ? 1'h0 : _GEN_14956; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16085 = 5'hd == rob_tail ? 1'h0 : _GEN_14957; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16086 = 5'he == rob_tail ? 1'h0 : _GEN_14958; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16087 = 5'hf == rob_tail ? 1'h0 : _GEN_14959; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16088 = 5'h10 == rob_tail ? 1'h0 : _GEN_14960; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16089 = 5'h11 == rob_tail ? 1'h0 : _GEN_14961; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16090 = 5'h12 == rob_tail ? 1'h0 : _GEN_14962; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16091 = 5'h13 == rob_tail ? 1'h0 : _GEN_14963; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16092 = 5'h14 == rob_tail ? 1'h0 : _GEN_14964; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16093 = 5'h15 == rob_tail ? 1'h0 : _GEN_14965; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16094 = 5'h16 == rob_tail ? 1'h0 : _GEN_14966; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16095 = 5'h17 == rob_tail ? 1'h0 : _GEN_14967; // @[rob.scala 353:52 rob.scala 353:52]
  wire  _GEN_16096 = io_dis_valids_1 ? _GEN_14176 : T_35634_0; // @[rob.scala 346:7]
  wire  _GEN_16097 = io_dis_valids_1 ? _GEN_14177 : T_35634_1; // @[rob.scala 346:7]
  wire  _GEN_16098 = io_dis_valids_1 ? _GEN_14178 : T_35634_2; // @[rob.scala 346:7]
  wire  _GEN_16099 = io_dis_valids_1 ? _GEN_14179 : T_35634_3; // @[rob.scala 346:7]
  wire  _GEN_16100 = io_dis_valids_1 ? _GEN_14180 : T_35634_4; // @[rob.scala 346:7]
  wire  _GEN_16101 = io_dis_valids_1 ? _GEN_14181 : T_35634_5; // @[rob.scala 346:7]
  wire  _GEN_16102 = io_dis_valids_1 ? _GEN_14182 : T_35634_6; // @[rob.scala 346:7]
  wire  _GEN_16103 = io_dis_valids_1 ? _GEN_14183 : T_35634_7; // @[rob.scala 346:7]
  wire  _GEN_16104 = io_dis_valids_1 ? _GEN_14184 : T_35634_8; // @[rob.scala 346:7]
  wire  _GEN_16105 = io_dis_valids_1 ? _GEN_14185 : T_35634_9; // @[rob.scala 346:7]
  wire  _GEN_16106 = io_dis_valids_1 ? _GEN_14186 : T_35634_10; // @[rob.scala 346:7]
  wire  _GEN_16107 = io_dis_valids_1 ? _GEN_14187 : T_35634_11; // @[rob.scala 346:7]
  wire  _GEN_16108 = io_dis_valids_1 ? _GEN_14188 : T_35634_12; // @[rob.scala 346:7]
  wire  _GEN_16109 = io_dis_valids_1 ? _GEN_14189 : T_35634_13; // @[rob.scala 346:7]
  wire  _GEN_16110 = io_dis_valids_1 ? _GEN_14190 : T_35634_14; // @[rob.scala 346:7]
  wire  _GEN_16111 = io_dis_valids_1 ? _GEN_14191 : T_35634_15; // @[rob.scala 346:7]
  wire  _GEN_16112 = io_dis_valids_1 ? _GEN_14192 : T_35634_16; // @[rob.scala 346:7]
  wire  _GEN_16113 = io_dis_valids_1 ? _GEN_14193 : T_35634_17; // @[rob.scala 346:7]
  wire  _GEN_16114 = io_dis_valids_1 ? _GEN_14194 : T_35634_18; // @[rob.scala 346:7]
  wire  _GEN_16115 = io_dis_valids_1 ? _GEN_14195 : T_35634_19; // @[rob.scala 346:7]
  wire  _GEN_16116 = io_dis_valids_1 ? _GEN_14196 : T_35634_20; // @[rob.scala 346:7]
  wire  _GEN_16117 = io_dis_valids_1 ? _GEN_14197 : T_35634_21; // @[rob.scala 346:7]
  wire  _GEN_16118 = io_dis_valids_1 ? _GEN_14198 : T_35634_22; // @[rob.scala 346:7]
  wire  _GEN_16119 = io_dis_valids_1 ? _GEN_14199 : T_35634_23; // @[rob.scala 346:7]
  wire [31:0] _GEN_16197 = io_dis_valids_1 ? _GEN_14272 : T_38110_0_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16198 = io_dis_valids_1 ? _GEN_14273 : T_38110_1_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16199 = io_dis_valids_1 ? _GEN_14274 : T_38110_2_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16200 = io_dis_valids_1 ? _GEN_14275 : T_38110_3_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16201 = io_dis_valids_1 ? _GEN_14276 : T_38110_4_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16202 = io_dis_valids_1 ? _GEN_14277 : T_38110_5_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16203 = io_dis_valids_1 ? _GEN_14278 : T_38110_6_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16204 = io_dis_valids_1 ? _GEN_14279 : T_38110_7_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16205 = io_dis_valids_1 ? _GEN_14280 : T_38110_8_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16206 = io_dis_valids_1 ? _GEN_14281 : T_38110_9_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16207 = io_dis_valids_1 ? _GEN_14282 : T_38110_10_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16208 = io_dis_valids_1 ? _GEN_14283 : T_38110_11_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16209 = io_dis_valids_1 ? _GEN_14284 : T_38110_12_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16210 = io_dis_valids_1 ? _GEN_14285 : T_38110_13_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16211 = io_dis_valids_1 ? _GEN_14286 : T_38110_14_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16212 = io_dis_valids_1 ? _GEN_14287 : T_38110_15_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16213 = io_dis_valids_1 ? _GEN_14288 : T_38110_16_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16214 = io_dis_valids_1 ? _GEN_14289 : T_38110_17_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16215 = io_dis_valids_1 ? _GEN_14290 : T_38110_18_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16216 = io_dis_valids_1 ? _GEN_14291 : T_38110_19_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16217 = io_dis_valids_1 ? _GEN_14292 : T_38110_20_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16218 = io_dis_valids_1 ? _GEN_14293 : T_38110_21_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16219 = io_dis_valids_1 ? _GEN_14294 : T_38110_22_inst; // @[rob.scala 346:7]
  wire [31:0] _GEN_16220 = io_dis_valids_1 ? _GEN_14295 : T_38110_23_inst; // @[rob.scala 346:7]
  wire  _GEN_16869 = io_dis_valids_1 ? _GEN_16072 : T_38110_0_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16870 = io_dis_valids_1 ? _GEN_16073 : T_38110_1_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16871 = io_dis_valids_1 ? _GEN_16074 : T_38110_2_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16872 = io_dis_valids_1 ? _GEN_16075 : T_38110_3_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16873 = io_dis_valids_1 ? _GEN_16076 : T_38110_4_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16874 = io_dis_valids_1 ? _GEN_16077 : T_38110_5_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16875 = io_dis_valids_1 ? _GEN_16078 : T_38110_6_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16876 = io_dis_valids_1 ? _GEN_16079 : T_38110_7_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16877 = io_dis_valids_1 ? _GEN_16080 : T_38110_8_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16878 = io_dis_valids_1 ? _GEN_16081 : T_38110_9_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16879 = io_dis_valids_1 ? _GEN_16082 : T_38110_10_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16880 = io_dis_valids_1 ? _GEN_16083 : T_38110_11_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16881 = io_dis_valids_1 ? _GEN_16084 : T_38110_12_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16882 = io_dis_valids_1 ? _GEN_16085 : T_38110_13_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16883 = io_dis_valids_1 ? _GEN_16086 : T_38110_14_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16884 = io_dis_valids_1 ? _GEN_16087 : T_38110_15_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16885 = io_dis_valids_1 ? _GEN_16088 : T_38110_16_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16886 = io_dis_valids_1 ? _GEN_16089 : T_38110_17_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16887 = io_dis_valids_1 ? _GEN_16090 : T_38110_18_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16888 = io_dis_valids_1 ? _GEN_16091 : T_38110_19_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16889 = io_dis_valids_1 ? _GEN_16092 : T_38110_20_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16890 = io_dis_valids_1 ? _GEN_16093 : T_38110_21_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16891 = io_dis_valids_1 ? _GEN_16094 : T_38110_22_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16892 = io_dis_valids_1 ? _GEN_16095 : T_38110_23_stat_brjmp_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16893 = io_dis_valids_1 ? _GEN_14968 : T_38110_0_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16894 = io_dis_valids_1 ? _GEN_14969 : T_38110_1_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16895 = io_dis_valids_1 ? _GEN_14970 : T_38110_2_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16896 = io_dis_valids_1 ? _GEN_14971 : T_38110_3_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16897 = io_dis_valids_1 ? _GEN_14972 : T_38110_4_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16898 = io_dis_valids_1 ? _GEN_14973 : T_38110_5_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16899 = io_dis_valids_1 ? _GEN_14974 : T_38110_6_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16900 = io_dis_valids_1 ? _GEN_14975 : T_38110_7_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16901 = io_dis_valids_1 ? _GEN_14976 : T_38110_8_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16902 = io_dis_valids_1 ? _GEN_14977 : T_38110_9_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16903 = io_dis_valids_1 ? _GEN_14978 : T_38110_10_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16904 = io_dis_valids_1 ? _GEN_14979 : T_38110_11_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16905 = io_dis_valids_1 ? _GEN_14980 : T_38110_12_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16906 = io_dis_valids_1 ? _GEN_14981 : T_38110_13_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16907 = io_dis_valids_1 ? _GEN_14982 : T_38110_14_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16908 = io_dis_valids_1 ? _GEN_14983 : T_38110_15_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16909 = io_dis_valids_1 ? _GEN_14984 : T_38110_16_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16910 = io_dis_valids_1 ? _GEN_14985 : T_38110_17_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16911 = io_dis_valids_1 ? _GEN_14986 : T_38110_18_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16912 = io_dis_valids_1 ? _GEN_14987 : T_38110_19_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16913 = io_dis_valids_1 ? _GEN_14988 : T_38110_20_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16914 = io_dis_valids_1 ? _GEN_14989 : T_38110_21_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16915 = io_dis_valids_1 ? _GEN_14990 : T_38110_22_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16916 = io_dis_valids_1 ? _GEN_14991 : T_38110_23_stat_btb_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16917 = io_dis_valids_1 ? _GEN_14992 : T_38110_0_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16918 = io_dis_valids_1 ? _GEN_14993 : T_38110_1_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16919 = io_dis_valids_1 ? _GEN_14994 : T_38110_2_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16920 = io_dis_valids_1 ? _GEN_14995 : T_38110_3_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16921 = io_dis_valids_1 ? _GEN_14996 : T_38110_4_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16922 = io_dis_valids_1 ? _GEN_14997 : T_38110_5_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16923 = io_dis_valids_1 ? _GEN_14998 : T_38110_6_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16924 = io_dis_valids_1 ? _GEN_14999 : T_38110_7_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16925 = io_dis_valids_1 ? _GEN_15000 : T_38110_8_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16926 = io_dis_valids_1 ? _GEN_15001 : T_38110_9_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16927 = io_dis_valids_1 ? _GEN_15002 : T_38110_10_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16928 = io_dis_valids_1 ? _GEN_15003 : T_38110_11_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16929 = io_dis_valids_1 ? _GEN_15004 : T_38110_12_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16930 = io_dis_valids_1 ? _GEN_15005 : T_38110_13_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16931 = io_dis_valids_1 ? _GEN_15006 : T_38110_14_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16932 = io_dis_valids_1 ? _GEN_15007 : T_38110_15_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16933 = io_dis_valids_1 ? _GEN_15008 : T_38110_16_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16934 = io_dis_valids_1 ? _GEN_15009 : T_38110_17_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16935 = io_dis_valids_1 ? _GEN_15010 : T_38110_18_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16936 = io_dis_valids_1 ? _GEN_15011 : T_38110_19_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16937 = io_dis_valids_1 ? _GEN_15012 : T_38110_20_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16938 = io_dis_valids_1 ? _GEN_15013 : T_38110_21_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16939 = io_dis_valids_1 ? _GEN_15014 : T_38110_22_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16940 = io_dis_valids_1 ? _GEN_15015 : T_38110_23_stat_btb_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16941 = io_dis_valids_1 ? _GEN_15016 : T_38110_0_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16942 = io_dis_valids_1 ? _GEN_15017 : T_38110_1_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16943 = io_dis_valids_1 ? _GEN_15018 : T_38110_2_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16944 = io_dis_valids_1 ? _GEN_15019 : T_38110_3_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16945 = io_dis_valids_1 ? _GEN_15020 : T_38110_4_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16946 = io_dis_valids_1 ? _GEN_15021 : T_38110_5_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16947 = io_dis_valids_1 ? _GEN_15022 : T_38110_6_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16948 = io_dis_valids_1 ? _GEN_15023 : T_38110_7_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16949 = io_dis_valids_1 ? _GEN_15024 : T_38110_8_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16950 = io_dis_valids_1 ? _GEN_15025 : T_38110_9_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16951 = io_dis_valids_1 ? _GEN_15026 : T_38110_10_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16952 = io_dis_valids_1 ? _GEN_15027 : T_38110_11_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16953 = io_dis_valids_1 ? _GEN_15028 : T_38110_12_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16954 = io_dis_valids_1 ? _GEN_15029 : T_38110_13_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16955 = io_dis_valids_1 ? _GEN_15030 : T_38110_14_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16956 = io_dis_valids_1 ? _GEN_15031 : T_38110_15_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16957 = io_dis_valids_1 ? _GEN_15032 : T_38110_16_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16958 = io_dis_valids_1 ? _GEN_15033 : T_38110_17_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16959 = io_dis_valids_1 ? _GEN_15034 : T_38110_18_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16960 = io_dis_valids_1 ? _GEN_15035 : T_38110_19_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16961 = io_dis_valids_1 ? _GEN_15036 : T_38110_20_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16962 = io_dis_valids_1 ? _GEN_15037 : T_38110_21_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16963 = io_dis_valids_1 ? _GEN_15038 : T_38110_22_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16964 = io_dis_valids_1 ? _GEN_15039 : T_38110_23_stat_bpd_made_pred; // @[rob.scala 346:7]
  wire  _GEN_16965 = io_dis_valids_1 ? _GEN_15040 : T_38110_0_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16966 = io_dis_valids_1 ? _GEN_15041 : T_38110_1_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16967 = io_dis_valids_1 ? _GEN_15042 : T_38110_2_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16968 = io_dis_valids_1 ? _GEN_15043 : T_38110_3_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16969 = io_dis_valids_1 ? _GEN_15044 : T_38110_4_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16970 = io_dis_valids_1 ? _GEN_15045 : T_38110_5_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16971 = io_dis_valids_1 ? _GEN_15046 : T_38110_6_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16972 = io_dis_valids_1 ? _GEN_15047 : T_38110_7_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16973 = io_dis_valids_1 ? _GEN_15048 : T_38110_8_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16974 = io_dis_valids_1 ? _GEN_15049 : T_38110_9_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16975 = io_dis_valids_1 ? _GEN_15050 : T_38110_10_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16976 = io_dis_valids_1 ? _GEN_15051 : T_38110_11_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16977 = io_dis_valids_1 ? _GEN_15052 : T_38110_12_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16978 = io_dis_valids_1 ? _GEN_15053 : T_38110_13_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16979 = io_dis_valids_1 ? _GEN_15054 : T_38110_14_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16980 = io_dis_valids_1 ? _GEN_15055 : T_38110_15_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16981 = io_dis_valids_1 ? _GEN_15056 : T_38110_16_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16982 = io_dis_valids_1 ? _GEN_15057 : T_38110_17_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16983 = io_dis_valids_1 ? _GEN_15058 : T_38110_18_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16984 = io_dis_valids_1 ? _GEN_15059 : T_38110_19_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16985 = io_dis_valids_1 ? _GEN_15060 : T_38110_20_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16986 = io_dis_valids_1 ? _GEN_15061 : T_38110_21_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16987 = io_dis_valids_1 ? _GEN_15062 : T_38110_22_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire  _GEN_16988 = io_dis_valids_1 ? _GEN_15063 : T_38110_23_stat_bpd_mispredicted; // @[rob.scala 346:7]
  wire [63:0] _GEN_17949 = io_dis_valids_1 ? _GEN_16024 : T_38110_0_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17950 = io_dis_valids_1 ? _GEN_16025 : T_38110_1_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17951 = io_dis_valids_1 ? _GEN_16026 : T_38110_2_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17952 = io_dis_valids_1 ? _GEN_16027 : T_38110_3_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17953 = io_dis_valids_1 ? _GEN_16028 : T_38110_4_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17954 = io_dis_valids_1 ? _GEN_16029 : T_38110_5_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17955 = io_dis_valids_1 ? _GEN_16030 : T_38110_6_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17956 = io_dis_valids_1 ? _GEN_16031 : T_38110_7_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17957 = io_dis_valids_1 ? _GEN_16032 : T_38110_8_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17958 = io_dis_valids_1 ? _GEN_16033 : T_38110_9_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17959 = io_dis_valids_1 ? _GEN_16034 : T_38110_10_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17960 = io_dis_valids_1 ? _GEN_16035 : T_38110_11_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17961 = io_dis_valids_1 ? _GEN_16036 : T_38110_12_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17962 = io_dis_valids_1 ? _GEN_16037 : T_38110_13_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17963 = io_dis_valids_1 ? _GEN_16038 : T_38110_14_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17964 = io_dis_valids_1 ? _GEN_16039 : T_38110_15_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17965 = io_dis_valids_1 ? _GEN_16040 : T_38110_16_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17966 = io_dis_valids_1 ? _GEN_16041 : T_38110_17_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17967 = io_dis_valids_1 ? _GEN_16042 : T_38110_18_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17968 = io_dis_valids_1 ? _GEN_16043 : T_38110_19_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17969 = io_dis_valids_1 ? _GEN_16044 : T_38110_20_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17970 = io_dis_valids_1 ? _GEN_16045 : T_38110_21_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17971 = io_dis_valids_1 ? _GEN_16046 : T_38110_22_debug_wdata; // @[rob.scala 346:7]
  wire [63:0] _GEN_17972 = io_dis_valids_1 ? _GEN_16047 : T_38110_23_debug_wdata; // @[rob.scala 346:7]
  wire  _GEN_18000 = 5'h1 == rob_tail ? T_35634_1 : T_35634_0; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18001 = 5'h2 == rob_tail ? T_35634_2 : _GEN_18000; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18002 = 5'h3 == rob_tail ? T_35634_3 : _GEN_18001; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18003 = 5'h4 == rob_tail ? T_35634_4 : _GEN_18002; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18004 = 5'h5 == rob_tail ? T_35634_5 : _GEN_18003; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18005 = 5'h6 == rob_tail ? T_35634_6 : _GEN_18004; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18006 = 5'h7 == rob_tail ? T_35634_7 : _GEN_18005; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18007 = 5'h8 == rob_tail ? T_35634_8 : _GEN_18006; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18008 = 5'h9 == rob_tail ? T_35634_9 : _GEN_18007; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18009 = 5'ha == rob_tail ? T_35634_10 : _GEN_18008; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18010 = 5'hb == rob_tail ? T_35634_11 : _GEN_18009; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18011 = 5'hc == rob_tail ? T_35634_12 : _GEN_18010; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18012 = 5'hd == rob_tail ? T_35634_13 : _GEN_18011; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18013 = 5'he == rob_tail ? T_35634_14 : _GEN_18012; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18014 = 5'hf == rob_tail ? T_35634_15 : _GEN_18013; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18015 = 5'h10 == rob_tail ? T_35634_16 : _GEN_18014; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18016 = 5'h11 == rob_tail ? T_35634_17 : _GEN_18015; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18017 = 5'h12 == rob_tail ? T_35634_18 : _GEN_18016; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18018 = 5'h13 == rob_tail ? T_35634_19 : _GEN_18017; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18019 = 5'h14 == rob_tail ? T_35634_20 : _GEN_18018; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18020 = 5'h15 == rob_tail ? T_35634_21 : _GEN_18019; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18021 = 5'h16 == rob_tail ? T_35634_22 : _GEN_18020; // @[rob.scala 355:47 rob.scala 355:47]
  wire  _GEN_18022 = 5'h17 == rob_tail ? T_35634_23 : _GEN_18021; // @[rob.scala 355:47 rob.scala 355:47]
  wire  T_40426 = ~_GEN_18022; // @[rob.scala 355:47]
  wire  T_40427 = T_23559 & T_40426; // @[rob.scala 355:44]
  wire  T_40429 = ~io_dis_valids_1; // @[rob.scala 346:7]
  wire  T_40430 = T_40429 & T_40427; // @[rob.scala 356:7]
  wire [31:0] _GEN_18023 = 5'h0 == rob_tail ? 32'h4033 : _GEN_16197; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18024 = 5'h1 == rob_tail ? 32'h4033 : _GEN_16198; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18025 = 5'h2 == rob_tail ? 32'h4033 : _GEN_16199; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18026 = 5'h3 == rob_tail ? 32'h4033 : _GEN_16200; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18027 = 5'h4 == rob_tail ? 32'h4033 : _GEN_16201; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18028 = 5'h5 == rob_tail ? 32'h4033 : _GEN_16202; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18029 = 5'h6 == rob_tail ? 32'h4033 : _GEN_16203; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18030 = 5'h7 == rob_tail ? 32'h4033 : _GEN_16204; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18031 = 5'h8 == rob_tail ? 32'h4033 : _GEN_16205; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18032 = 5'h9 == rob_tail ? 32'h4033 : _GEN_16206; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18033 = 5'ha == rob_tail ? 32'h4033 : _GEN_16207; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18034 = 5'hb == rob_tail ? 32'h4033 : _GEN_16208; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18035 = 5'hc == rob_tail ? 32'h4033 : _GEN_16209; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18036 = 5'hd == rob_tail ? 32'h4033 : _GEN_16210; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18037 = 5'he == rob_tail ? 32'h4033 : _GEN_16211; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18038 = 5'hf == rob_tail ? 32'h4033 : _GEN_16212; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18039 = 5'h10 == rob_tail ? 32'h4033 : _GEN_16213; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18040 = 5'h11 == rob_tail ? 32'h4033 : _GEN_16214; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18041 = 5'h12 == rob_tail ? 32'h4033 : _GEN_16215; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18042 = 5'h13 == rob_tail ? 32'h4033 : _GEN_16216; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18043 = 5'h14 == rob_tail ? 32'h4033 : _GEN_16217; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18044 = 5'h15 == rob_tail ? 32'h4033 : _GEN_16218; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18045 = 5'h16 == rob_tail ? 32'h4033 : _GEN_16219; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18046 = 5'h17 == rob_tail ? 32'h4033 : _GEN_16220; // @[rob.scala 357:33 rob.scala 357:33]
  wire [31:0] _GEN_18047 = T_40430 ? _GEN_18023 : _GEN_16197; // @[rob.scala 356:7]
  wire [31:0] _GEN_18048 = T_40430 ? _GEN_18024 : _GEN_16198; // @[rob.scala 356:7]
  wire [31:0] _GEN_18049 = T_40430 ? _GEN_18025 : _GEN_16199; // @[rob.scala 356:7]
  wire [31:0] _GEN_18050 = T_40430 ? _GEN_18026 : _GEN_16200; // @[rob.scala 356:7]
  wire [31:0] _GEN_18051 = T_40430 ? _GEN_18027 : _GEN_16201; // @[rob.scala 356:7]
  wire [31:0] _GEN_18052 = T_40430 ? _GEN_18028 : _GEN_16202; // @[rob.scala 356:7]
  wire [31:0] _GEN_18053 = T_40430 ? _GEN_18029 : _GEN_16203; // @[rob.scala 356:7]
  wire [31:0] _GEN_18054 = T_40430 ? _GEN_18030 : _GEN_16204; // @[rob.scala 356:7]
  wire [31:0] _GEN_18055 = T_40430 ? _GEN_18031 : _GEN_16205; // @[rob.scala 356:7]
  wire [31:0] _GEN_18056 = T_40430 ? _GEN_18032 : _GEN_16206; // @[rob.scala 356:7]
  wire [31:0] _GEN_18057 = T_40430 ? _GEN_18033 : _GEN_16207; // @[rob.scala 356:7]
  wire [31:0] _GEN_18058 = T_40430 ? _GEN_18034 : _GEN_16208; // @[rob.scala 356:7]
  wire [31:0] _GEN_18059 = T_40430 ? _GEN_18035 : _GEN_16209; // @[rob.scala 356:7]
  wire [31:0] _GEN_18060 = T_40430 ? _GEN_18036 : _GEN_16210; // @[rob.scala 356:7]
  wire [31:0] _GEN_18061 = T_40430 ? _GEN_18037 : _GEN_16211; // @[rob.scala 356:7]
  wire [31:0] _GEN_18062 = T_40430 ? _GEN_18038 : _GEN_16212; // @[rob.scala 356:7]
  wire [31:0] _GEN_18063 = T_40430 ? _GEN_18039 : _GEN_16213; // @[rob.scala 356:7]
  wire [31:0] _GEN_18064 = T_40430 ? _GEN_18040 : _GEN_16214; // @[rob.scala 356:7]
  wire [31:0] _GEN_18065 = T_40430 ? _GEN_18041 : _GEN_16215; // @[rob.scala 356:7]
  wire [31:0] _GEN_18066 = T_40430 ? _GEN_18042 : _GEN_16216; // @[rob.scala 356:7]
  wire [31:0] _GEN_18067 = T_40430 ? _GEN_18043 : _GEN_16217; // @[rob.scala 356:7]
  wire [31:0] _GEN_18068 = T_40430 ? _GEN_18044 : _GEN_16218; // @[rob.scala 356:7]
  wire [31:0] _GEN_18069 = T_40430 ? _GEN_18045 : _GEN_16219; // @[rob.scala 356:7]
  wire [31:0] _GEN_18070 = T_40430 ? _GEN_18046 : _GEN_16220; // @[rob.scala 356:7]
  wire  T_40521 = io_wb_resps_0_valid & T_28590; // @[rob.scala 368:30]
  wire  T_40529 = io_wb_resps_1_valid & T_28598; // @[rob.scala 368:30]
  wire  T_40537 = io_wb_resps_2_valid & T_28606; // @[rob.scala 368:30]
  wire  T_40551 = io_brinfo_valid & T_28620; // @[rob.scala 400:29]
  wire  _GEN_18375 = 5'h1 == T_29096 ? T_35634_1 : T_35634_0; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18376 = 5'h2 == T_29096 ? T_35634_2 : _GEN_18375; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18377 = 5'h3 == T_29096 ? T_35634_3 : _GEN_18376; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18378 = 5'h4 == T_29096 ? T_35634_4 : _GEN_18377; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18379 = 5'h5 == T_29096 ? T_35634_5 : _GEN_18378; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18380 = 5'h6 == T_29096 ? T_35634_6 : _GEN_18379; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18381 = 5'h7 == T_29096 ? T_35634_7 : _GEN_18380; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18382 = 5'h8 == T_29096 ? T_35634_8 : _GEN_18381; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18383 = 5'h9 == T_29096 ? T_35634_9 : _GEN_18382; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18384 = 5'ha == T_29096 ? T_35634_10 : _GEN_18383; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18385 = 5'hb == T_29096 ? T_35634_11 : _GEN_18384; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18386 = 5'hc == T_29096 ? T_35634_12 : _GEN_18385; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18387 = 5'hd == T_29096 ? T_35634_13 : _GEN_18386; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18388 = 5'he == T_29096 ? T_35634_14 : _GEN_18387; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18389 = 5'hf == T_29096 ? T_35634_15 : _GEN_18388; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18390 = 5'h10 == T_29096 ? T_35634_16 : _GEN_18389; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18391 = 5'h11 == T_29096 ? T_35634_17 : _GEN_18390; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18392 = 5'h12 == T_29096 ? T_35634_18 : _GEN_18391; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18393 = 5'h13 == T_29096 ? T_35634_19 : _GEN_18392; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18394 = 5'h14 == T_29096 ? T_35634_20 : _GEN_18393; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18395 = 5'h15 == T_29096 ? T_35634_21 : _GEN_18394; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18396 = 5'h16 == T_29096 ? T_35634_22 : _GEN_18395; // @[rob.scala 451:58 rob.scala 451:58]
  wire  _GEN_18397 = 5'h17 == T_29096 ? T_35634_23 : _GEN_18396; // @[rob.scala 451:58 rob.scala 451:58]
  wire  T_41027 = T_29097 & _GEN_18397; // @[rob.scala 451:58]
  wire  _GEN_18476 = 5'h1 == T_29096 ? T_38110_1_valid : T_38110_0_valid; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18477 = 5'h1 == T_29096 ? T_38110_1_iw_state : T_38110_0_iw_state; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18478 = 5'h1 == T_29096 ? T_38110_1_uopc : T_38110_0_uopc; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18479 = 5'h1 == T_29096 ? T_38110_1_inst : T_38110_0_inst; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18480 = 5'h1 == T_29096 ? T_38110_1_pc : T_38110_0_pc; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18481 = 5'h1 == T_29096 ? T_38110_1_fu_code : T_38110_0_fu_code; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18482 = 5'h1 == T_29096 ? T_38110_1_ctrl_br_type : T_38110_0_ctrl_br_type; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18483 = 5'h1 == T_29096 ? T_38110_1_ctrl_op1_sel : T_38110_0_ctrl_op1_sel; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18484 = 5'h1 == T_29096 ? T_38110_1_ctrl_op2_sel : T_38110_0_ctrl_op2_sel; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18485 = 5'h1 == T_29096 ? T_38110_1_ctrl_imm_sel : T_38110_0_ctrl_imm_sel; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18486 = 5'h1 == T_29096 ? T_38110_1_ctrl_op_fcn : T_38110_0_ctrl_op_fcn; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18487 = 5'h1 == T_29096 ? T_38110_1_ctrl_fcn_dw : T_38110_0_ctrl_fcn_dw; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18488 = 5'h1 == T_29096 ? T_38110_1_ctrl_rf_wen : T_38110_0_ctrl_rf_wen; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18489 = 5'h1 == T_29096 ? T_38110_1_ctrl_csr_cmd : T_38110_0_ctrl_csr_cmd; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18490 = 5'h1 == T_29096 ? T_38110_1_ctrl_is_load : T_38110_0_ctrl_is_load; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18491 = 5'h1 == T_29096 ? T_38110_1_ctrl_is_sta : T_38110_0_ctrl_is_sta; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18492 = 5'h1 == T_29096 ? T_38110_1_ctrl_is_std : T_38110_0_ctrl_is_std; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18493 = 5'h1 == T_29096 ? T_38110_1_wakeup_delay : T_38110_0_wakeup_delay; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18494 = 5'h1 == T_29096 ? T_38110_1_allocate_brtag : T_38110_0_allocate_brtag; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18495 = 5'h1 == T_29096 ? T_38110_1_is_br_or_jmp : T_38110_0_is_br_or_jmp; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18496 = 5'h1 == T_29096 ? T_38110_1_is_jump : T_38110_0_is_jump; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18497 = 5'h1 == T_29096 ? T_38110_1_is_jal : T_38110_0_is_jal; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18498 = 5'h1 == T_29096 ? T_38110_1_is_ret : T_38110_0_is_ret; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18499 = 5'h1 == T_29096 ? T_38110_1_is_call : T_38110_0_is_call; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18500 = 5'h1 == T_29096 ? T_38110_1_br_mask : T_38110_0_br_mask; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18501 = 5'h1 == T_29096 ? T_38110_1_br_tag : T_38110_0_br_tag; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18502 = 5'h1 == T_29096 ? T_38110_1_br_prediction_bpd_predict_val : T_38110_0_br_prediction_bpd_predict_val
    ; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18503 = 5'h1 == T_29096 ? T_38110_1_br_prediction_bpd_predict_taken :
    T_38110_0_br_prediction_bpd_predict_taken; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18504 = 5'h1 == T_29096 ? T_38110_1_br_prediction_btb_hit : T_38110_0_br_prediction_btb_hit; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18505 = 5'h1 == T_29096 ? T_38110_1_br_prediction_btb_predicted : T_38110_0_br_prediction_btb_predicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18506 = 5'h1 == T_29096 ? T_38110_1_br_prediction_is_br_or_jalr : T_38110_0_br_prediction_is_br_or_jalr; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18507 = 5'h1 == T_29096 ? T_38110_1_stat_brjmp_mispredicted : T_38110_0_stat_brjmp_mispredicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18508 = 5'h1 == T_29096 ? T_38110_1_stat_btb_made_pred : T_38110_0_stat_btb_made_pred; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18509 = 5'h1 == T_29096 ? T_38110_1_stat_btb_mispredicted : T_38110_0_stat_btb_mispredicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18510 = 5'h1 == T_29096 ? T_38110_1_stat_bpd_made_pred : T_38110_0_stat_bpd_made_pred; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18511 = 5'h1 == T_29096 ? T_38110_1_stat_bpd_mispredicted : T_38110_0_stat_bpd_mispredicted; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18512 = 5'h1 == T_29096 ? T_38110_1_fetch_pc_lob : T_38110_0_fetch_pc_lob; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18513 = 5'h1 == T_29096 ? T_38110_1_imm_packed : T_38110_0_imm_packed; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18514 = 5'h1 == T_29096 ? T_38110_1_csr_addr : T_38110_0_csr_addr; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18515 = 5'h1 == T_29096 ? T_38110_1_rob_idx : T_38110_0_rob_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18516 = 5'h1 == T_29096 ? T_38110_1_ldq_idx : T_38110_0_ldq_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18517 = 5'h1 == T_29096 ? T_38110_1_stq_idx : T_38110_0_stq_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18518 = 5'h1 == T_29096 ? T_38110_1_brob_idx : T_38110_0_brob_idx; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18519 = 5'h1 == T_29096 ? T_38110_1_pdst : T_38110_0_pdst; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18520 = 5'h1 == T_29096 ? T_38110_1_pop1 : T_38110_0_pop1; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18521 = 5'h1 == T_29096 ? T_38110_1_pop2 : T_38110_0_pop2; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18522 = 5'h1 == T_29096 ? T_38110_1_pop3 : T_38110_0_pop3; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18523 = 5'h1 == T_29096 ? T_38110_1_prs1_busy : T_38110_0_prs1_busy; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18524 = 5'h1 == T_29096 ? T_38110_1_prs2_busy : T_38110_0_prs2_busy; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18525 = 5'h1 == T_29096 ? T_38110_1_prs3_busy : T_38110_0_prs3_busy; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18526 = 5'h1 == T_29096 ? T_38110_1_stale_pdst : T_38110_0_stale_pdst; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18527 = 5'h1 == T_29096 ? T_38110_1_exception : T_38110_0_exception; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18528 = 5'h1 == T_29096 ? T_38110_1_exc_cause : T_38110_0_exc_cause; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18529 = 5'h1 == T_29096 ? T_38110_1_bypassable : T_38110_0_bypassable; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18530 = 5'h1 == T_29096 ? T_38110_1_mem_cmd : T_38110_0_mem_cmd; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18531 = 5'h1 == T_29096 ? T_38110_1_mem_typ : T_38110_0_mem_typ; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18532 = 5'h1 == T_29096 ? T_38110_1_is_fence : T_38110_0_is_fence; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18533 = 5'h1 == T_29096 ? T_38110_1_is_fencei : T_38110_0_is_fencei; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18534 = 5'h1 == T_29096 ? T_38110_1_is_store : T_38110_0_is_store; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18535 = 5'h1 == T_29096 ? T_38110_1_is_amo : T_38110_0_is_amo; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18536 = 5'h1 == T_29096 ? T_38110_1_is_load : T_38110_0_is_load; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18537 = 5'h1 == T_29096 ? T_38110_1_is_unique : T_38110_0_is_unique; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18538 = 5'h1 == T_29096 ? T_38110_1_flush_on_commit : T_38110_0_flush_on_commit; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18539 = 5'h1 == T_29096 ? T_38110_1_ldst : T_38110_0_ldst; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18540 = 5'h1 == T_29096 ? T_38110_1_lrs1 : T_38110_0_lrs1; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18541 = 5'h1 == T_29096 ? T_38110_1_lrs2 : T_38110_0_lrs2; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18542 = 5'h1 == T_29096 ? T_38110_1_lrs3 : T_38110_0_lrs3; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18543 = 5'h1 == T_29096 ? T_38110_1_ldst_val : T_38110_0_ldst_val; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18544 = 5'h1 == T_29096 ? T_38110_1_dst_rtype : T_38110_0_dst_rtype; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18545 = 5'h1 == T_29096 ? T_38110_1_lrs1_rtype : T_38110_0_lrs1_rtype; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18546 = 5'h1 == T_29096 ? T_38110_1_lrs2_rtype : T_38110_0_lrs2_rtype; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18547 = 5'h1 == T_29096 ? T_38110_1_frs3_en : T_38110_0_frs3_en; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18548 = 5'h1 == T_29096 ? T_38110_1_fp_val : T_38110_0_fp_val; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18549 = 5'h1 == T_29096 ? T_38110_1_fp_single : T_38110_0_fp_single; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18550 = 5'h1 == T_29096 ? T_38110_1_xcpt_if : T_38110_0_xcpt_if; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18551 = 5'h1 == T_29096 ? T_38110_1_replay_if : T_38110_0_replay_if; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18553 = 5'h1 == T_29096 ? T_38110_1_debug_events_fetch_seq : T_38110_0_debug_events_fetch_seq; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18554 = 5'h2 == T_29096 ? T_38110_2_valid : _GEN_18476; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18555 = 5'h2 == T_29096 ? T_38110_2_iw_state : _GEN_18477; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18556 = 5'h2 == T_29096 ? T_38110_2_uopc : _GEN_18478; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18557 = 5'h2 == T_29096 ? T_38110_2_inst : _GEN_18479; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18558 = 5'h2 == T_29096 ? T_38110_2_pc : _GEN_18480; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18559 = 5'h2 == T_29096 ? T_38110_2_fu_code : _GEN_18481; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18560 = 5'h2 == T_29096 ? T_38110_2_ctrl_br_type : _GEN_18482; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18561 = 5'h2 == T_29096 ? T_38110_2_ctrl_op1_sel : _GEN_18483; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18562 = 5'h2 == T_29096 ? T_38110_2_ctrl_op2_sel : _GEN_18484; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18563 = 5'h2 == T_29096 ? T_38110_2_ctrl_imm_sel : _GEN_18485; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18564 = 5'h2 == T_29096 ? T_38110_2_ctrl_op_fcn : _GEN_18486; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18565 = 5'h2 == T_29096 ? T_38110_2_ctrl_fcn_dw : _GEN_18487; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18566 = 5'h2 == T_29096 ? T_38110_2_ctrl_rf_wen : _GEN_18488; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18567 = 5'h2 == T_29096 ? T_38110_2_ctrl_csr_cmd : _GEN_18489; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18568 = 5'h2 == T_29096 ? T_38110_2_ctrl_is_load : _GEN_18490; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18569 = 5'h2 == T_29096 ? T_38110_2_ctrl_is_sta : _GEN_18491; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18570 = 5'h2 == T_29096 ? T_38110_2_ctrl_is_std : _GEN_18492; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18571 = 5'h2 == T_29096 ? T_38110_2_wakeup_delay : _GEN_18493; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18572 = 5'h2 == T_29096 ? T_38110_2_allocate_brtag : _GEN_18494; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18573 = 5'h2 == T_29096 ? T_38110_2_is_br_or_jmp : _GEN_18495; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18574 = 5'h2 == T_29096 ? T_38110_2_is_jump : _GEN_18496; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18575 = 5'h2 == T_29096 ? T_38110_2_is_jal : _GEN_18497; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18576 = 5'h2 == T_29096 ? T_38110_2_is_ret : _GEN_18498; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18577 = 5'h2 == T_29096 ? T_38110_2_is_call : _GEN_18499; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18578 = 5'h2 == T_29096 ? T_38110_2_br_mask : _GEN_18500; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18579 = 5'h2 == T_29096 ? T_38110_2_br_tag : _GEN_18501; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18580 = 5'h2 == T_29096 ? T_38110_2_br_prediction_bpd_predict_val : _GEN_18502; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18581 = 5'h2 == T_29096 ? T_38110_2_br_prediction_bpd_predict_taken : _GEN_18503; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18582 = 5'h2 == T_29096 ? T_38110_2_br_prediction_btb_hit : _GEN_18504; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18583 = 5'h2 == T_29096 ? T_38110_2_br_prediction_btb_predicted : _GEN_18505; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18584 = 5'h2 == T_29096 ? T_38110_2_br_prediction_is_br_or_jalr : _GEN_18506; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18585 = 5'h2 == T_29096 ? T_38110_2_stat_brjmp_mispredicted : _GEN_18507; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18586 = 5'h2 == T_29096 ? T_38110_2_stat_btb_made_pred : _GEN_18508; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18587 = 5'h2 == T_29096 ? T_38110_2_stat_btb_mispredicted : _GEN_18509; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18588 = 5'h2 == T_29096 ? T_38110_2_stat_bpd_made_pred : _GEN_18510; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18589 = 5'h2 == T_29096 ? T_38110_2_stat_bpd_mispredicted : _GEN_18511; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18590 = 5'h2 == T_29096 ? T_38110_2_fetch_pc_lob : _GEN_18512; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18591 = 5'h2 == T_29096 ? T_38110_2_imm_packed : _GEN_18513; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18592 = 5'h2 == T_29096 ? T_38110_2_csr_addr : _GEN_18514; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18593 = 5'h2 == T_29096 ? T_38110_2_rob_idx : _GEN_18515; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18594 = 5'h2 == T_29096 ? T_38110_2_ldq_idx : _GEN_18516; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18595 = 5'h2 == T_29096 ? T_38110_2_stq_idx : _GEN_18517; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18596 = 5'h2 == T_29096 ? T_38110_2_brob_idx : _GEN_18518; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18597 = 5'h2 == T_29096 ? T_38110_2_pdst : _GEN_18519; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18598 = 5'h2 == T_29096 ? T_38110_2_pop1 : _GEN_18520; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18599 = 5'h2 == T_29096 ? T_38110_2_pop2 : _GEN_18521; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18600 = 5'h2 == T_29096 ? T_38110_2_pop3 : _GEN_18522; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18601 = 5'h2 == T_29096 ? T_38110_2_prs1_busy : _GEN_18523; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18602 = 5'h2 == T_29096 ? T_38110_2_prs2_busy : _GEN_18524; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18603 = 5'h2 == T_29096 ? T_38110_2_prs3_busy : _GEN_18525; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18604 = 5'h2 == T_29096 ? T_38110_2_stale_pdst : _GEN_18526; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18605 = 5'h2 == T_29096 ? T_38110_2_exception : _GEN_18527; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18606 = 5'h2 == T_29096 ? T_38110_2_exc_cause : _GEN_18528; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18607 = 5'h2 == T_29096 ? T_38110_2_bypassable : _GEN_18529; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18608 = 5'h2 == T_29096 ? T_38110_2_mem_cmd : _GEN_18530; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18609 = 5'h2 == T_29096 ? T_38110_2_mem_typ : _GEN_18531; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18610 = 5'h2 == T_29096 ? T_38110_2_is_fence : _GEN_18532; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18611 = 5'h2 == T_29096 ? T_38110_2_is_fencei : _GEN_18533; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18612 = 5'h2 == T_29096 ? T_38110_2_is_store : _GEN_18534; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18613 = 5'h2 == T_29096 ? T_38110_2_is_amo : _GEN_18535; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18614 = 5'h2 == T_29096 ? T_38110_2_is_load : _GEN_18536; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18615 = 5'h2 == T_29096 ? T_38110_2_is_unique : _GEN_18537; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18616 = 5'h2 == T_29096 ? T_38110_2_flush_on_commit : _GEN_18538; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18617 = 5'h2 == T_29096 ? T_38110_2_ldst : _GEN_18539; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18618 = 5'h2 == T_29096 ? T_38110_2_lrs1 : _GEN_18540; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18619 = 5'h2 == T_29096 ? T_38110_2_lrs2 : _GEN_18541; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18620 = 5'h2 == T_29096 ? T_38110_2_lrs3 : _GEN_18542; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18621 = 5'h2 == T_29096 ? T_38110_2_ldst_val : _GEN_18543; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18622 = 5'h2 == T_29096 ? T_38110_2_dst_rtype : _GEN_18544; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18623 = 5'h2 == T_29096 ? T_38110_2_lrs1_rtype : _GEN_18545; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18624 = 5'h2 == T_29096 ? T_38110_2_lrs2_rtype : _GEN_18546; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18625 = 5'h2 == T_29096 ? T_38110_2_frs3_en : _GEN_18547; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18626 = 5'h2 == T_29096 ? T_38110_2_fp_val : _GEN_18548; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18627 = 5'h2 == T_29096 ? T_38110_2_fp_single : _GEN_18549; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18628 = 5'h2 == T_29096 ? T_38110_2_xcpt_if : _GEN_18550; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18629 = 5'h2 == T_29096 ? T_38110_2_replay_if : _GEN_18551; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18631 = 5'h2 == T_29096 ? T_38110_2_debug_events_fetch_seq : _GEN_18553; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18632 = 5'h3 == T_29096 ? T_38110_3_valid : _GEN_18554; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18633 = 5'h3 == T_29096 ? T_38110_3_iw_state : _GEN_18555; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18634 = 5'h3 == T_29096 ? T_38110_3_uopc : _GEN_18556; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18635 = 5'h3 == T_29096 ? T_38110_3_inst : _GEN_18557; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18636 = 5'h3 == T_29096 ? T_38110_3_pc : _GEN_18558; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18637 = 5'h3 == T_29096 ? T_38110_3_fu_code : _GEN_18559; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18638 = 5'h3 == T_29096 ? T_38110_3_ctrl_br_type : _GEN_18560; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18639 = 5'h3 == T_29096 ? T_38110_3_ctrl_op1_sel : _GEN_18561; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18640 = 5'h3 == T_29096 ? T_38110_3_ctrl_op2_sel : _GEN_18562; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18641 = 5'h3 == T_29096 ? T_38110_3_ctrl_imm_sel : _GEN_18563; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18642 = 5'h3 == T_29096 ? T_38110_3_ctrl_op_fcn : _GEN_18564; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18643 = 5'h3 == T_29096 ? T_38110_3_ctrl_fcn_dw : _GEN_18565; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18644 = 5'h3 == T_29096 ? T_38110_3_ctrl_rf_wen : _GEN_18566; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18645 = 5'h3 == T_29096 ? T_38110_3_ctrl_csr_cmd : _GEN_18567; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18646 = 5'h3 == T_29096 ? T_38110_3_ctrl_is_load : _GEN_18568; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18647 = 5'h3 == T_29096 ? T_38110_3_ctrl_is_sta : _GEN_18569; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18648 = 5'h3 == T_29096 ? T_38110_3_ctrl_is_std : _GEN_18570; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18649 = 5'h3 == T_29096 ? T_38110_3_wakeup_delay : _GEN_18571; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18650 = 5'h3 == T_29096 ? T_38110_3_allocate_brtag : _GEN_18572; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18651 = 5'h3 == T_29096 ? T_38110_3_is_br_or_jmp : _GEN_18573; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18652 = 5'h3 == T_29096 ? T_38110_3_is_jump : _GEN_18574; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18653 = 5'h3 == T_29096 ? T_38110_3_is_jal : _GEN_18575; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18654 = 5'h3 == T_29096 ? T_38110_3_is_ret : _GEN_18576; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18655 = 5'h3 == T_29096 ? T_38110_3_is_call : _GEN_18577; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18656 = 5'h3 == T_29096 ? T_38110_3_br_mask : _GEN_18578; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18657 = 5'h3 == T_29096 ? T_38110_3_br_tag : _GEN_18579; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18658 = 5'h3 == T_29096 ? T_38110_3_br_prediction_bpd_predict_val : _GEN_18580; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18659 = 5'h3 == T_29096 ? T_38110_3_br_prediction_bpd_predict_taken : _GEN_18581; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18660 = 5'h3 == T_29096 ? T_38110_3_br_prediction_btb_hit : _GEN_18582; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18661 = 5'h3 == T_29096 ? T_38110_3_br_prediction_btb_predicted : _GEN_18583; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18662 = 5'h3 == T_29096 ? T_38110_3_br_prediction_is_br_or_jalr : _GEN_18584; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18663 = 5'h3 == T_29096 ? T_38110_3_stat_brjmp_mispredicted : _GEN_18585; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18664 = 5'h3 == T_29096 ? T_38110_3_stat_btb_made_pred : _GEN_18586; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18665 = 5'h3 == T_29096 ? T_38110_3_stat_btb_mispredicted : _GEN_18587; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18666 = 5'h3 == T_29096 ? T_38110_3_stat_bpd_made_pred : _GEN_18588; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18667 = 5'h3 == T_29096 ? T_38110_3_stat_bpd_mispredicted : _GEN_18589; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18668 = 5'h3 == T_29096 ? T_38110_3_fetch_pc_lob : _GEN_18590; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18669 = 5'h3 == T_29096 ? T_38110_3_imm_packed : _GEN_18591; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18670 = 5'h3 == T_29096 ? T_38110_3_csr_addr : _GEN_18592; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18671 = 5'h3 == T_29096 ? T_38110_3_rob_idx : _GEN_18593; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18672 = 5'h3 == T_29096 ? T_38110_3_ldq_idx : _GEN_18594; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18673 = 5'h3 == T_29096 ? T_38110_3_stq_idx : _GEN_18595; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18674 = 5'h3 == T_29096 ? T_38110_3_brob_idx : _GEN_18596; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18675 = 5'h3 == T_29096 ? T_38110_3_pdst : _GEN_18597; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18676 = 5'h3 == T_29096 ? T_38110_3_pop1 : _GEN_18598; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18677 = 5'h3 == T_29096 ? T_38110_3_pop2 : _GEN_18599; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18678 = 5'h3 == T_29096 ? T_38110_3_pop3 : _GEN_18600; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18679 = 5'h3 == T_29096 ? T_38110_3_prs1_busy : _GEN_18601; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18680 = 5'h3 == T_29096 ? T_38110_3_prs2_busy : _GEN_18602; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18681 = 5'h3 == T_29096 ? T_38110_3_prs3_busy : _GEN_18603; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18682 = 5'h3 == T_29096 ? T_38110_3_stale_pdst : _GEN_18604; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18683 = 5'h3 == T_29096 ? T_38110_3_exception : _GEN_18605; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18684 = 5'h3 == T_29096 ? T_38110_3_exc_cause : _GEN_18606; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18685 = 5'h3 == T_29096 ? T_38110_3_bypassable : _GEN_18607; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18686 = 5'h3 == T_29096 ? T_38110_3_mem_cmd : _GEN_18608; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18687 = 5'h3 == T_29096 ? T_38110_3_mem_typ : _GEN_18609; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18688 = 5'h3 == T_29096 ? T_38110_3_is_fence : _GEN_18610; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18689 = 5'h3 == T_29096 ? T_38110_3_is_fencei : _GEN_18611; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18690 = 5'h3 == T_29096 ? T_38110_3_is_store : _GEN_18612; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18691 = 5'h3 == T_29096 ? T_38110_3_is_amo : _GEN_18613; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18692 = 5'h3 == T_29096 ? T_38110_3_is_load : _GEN_18614; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18693 = 5'h3 == T_29096 ? T_38110_3_is_unique : _GEN_18615; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18694 = 5'h3 == T_29096 ? T_38110_3_flush_on_commit : _GEN_18616; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18695 = 5'h3 == T_29096 ? T_38110_3_ldst : _GEN_18617; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18696 = 5'h3 == T_29096 ? T_38110_3_lrs1 : _GEN_18618; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18697 = 5'h3 == T_29096 ? T_38110_3_lrs2 : _GEN_18619; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18698 = 5'h3 == T_29096 ? T_38110_3_lrs3 : _GEN_18620; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18699 = 5'h3 == T_29096 ? T_38110_3_ldst_val : _GEN_18621; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18700 = 5'h3 == T_29096 ? T_38110_3_dst_rtype : _GEN_18622; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18701 = 5'h3 == T_29096 ? T_38110_3_lrs1_rtype : _GEN_18623; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18702 = 5'h3 == T_29096 ? T_38110_3_lrs2_rtype : _GEN_18624; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18703 = 5'h3 == T_29096 ? T_38110_3_frs3_en : _GEN_18625; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18704 = 5'h3 == T_29096 ? T_38110_3_fp_val : _GEN_18626; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18705 = 5'h3 == T_29096 ? T_38110_3_fp_single : _GEN_18627; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18706 = 5'h3 == T_29096 ? T_38110_3_xcpt_if : _GEN_18628; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18707 = 5'h3 == T_29096 ? T_38110_3_replay_if : _GEN_18629; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18709 = 5'h3 == T_29096 ? T_38110_3_debug_events_fetch_seq : _GEN_18631; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18710 = 5'h4 == T_29096 ? T_38110_4_valid : _GEN_18632; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18711 = 5'h4 == T_29096 ? T_38110_4_iw_state : _GEN_18633; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18712 = 5'h4 == T_29096 ? T_38110_4_uopc : _GEN_18634; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18713 = 5'h4 == T_29096 ? T_38110_4_inst : _GEN_18635; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18714 = 5'h4 == T_29096 ? T_38110_4_pc : _GEN_18636; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18715 = 5'h4 == T_29096 ? T_38110_4_fu_code : _GEN_18637; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18716 = 5'h4 == T_29096 ? T_38110_4_ctrl_br_type : _GEN_18638; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18717 = 5'h4 == T_29096 ? T_38110_4_ctrl_op1_sel : _GEN_18639; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18718 = 5'h4 == T_29096 ? T_38110_4_ctrl_op2_sel : _GEN_18640; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18719 = 5'h4 == T_29096 ? T_38110_4_ctrl_imm_sel : _GEN_18641; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18720 = 5'h4 == T_29096 ? T_38110_4_ctrl_op_fcn : _GEN_18642; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18721 = 5'h4 == T_29096 ? T_38110_4_ctrl_fcn_dw : _GEN_18643; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18722 = 5'h4 == T_29096 ? T_38110_4_ctrl_rf_wen : _GEN_18644; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18723 = 5'h4 == T_29096 ? T_38110_4_ctrl_csr_cmd : _GEN_18645; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18724 = 5'h4 == T_29096 ? T_38110_4_ctrl_is_load : _GEN_18646; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18725 = 5'h4 == T_29096 ? T_38110_4_ctrl_is_sta : _GEN_18647; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18726 = 5'h4 == T_29096 ? T_38110_4_ctrl_is_std : _GEN_18648; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18727 = 5'h4 == T_29096 ? T_38110_4_wakeup_delay : _GEN_18649; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18728 = 5'h4 == T_29096 ? T_38110_4_allocate_brtag : _GEN_18650; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18729 = 5'h4 == T_29096 ? T_38110_4_is_br_or_jmp : _GEN_18651; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18730 = 5'h4 == T_29096 ? T_38110_4_is_jump : _GEN_18652; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18731 = 5'h4 == T_29096 ? T_38110_4_is_jal : _GEN_18653; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18732 = 5'h4 == T_29096 ? T_38110_4_is_ret : _GEN_18654; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18733 = 5'h4 == T_29096 ? T_38110_4_is_call : _GEN_18655; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18734 = 5'h4 == T_29096 ? T_38110_4_br_mask : _GEN_18656; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18735 = 5'h4 == T_29096 ? T_38110_4_br_tag : _GEN_18657; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18736 = 5'h4 == T_29096 ? T_38110_4_br_prediction_bpd_predict_val : _GEN_18658; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18737 = 5'h4 == T_29096 ? T_38110_4_br_prediction_bpd_predict_taken : _GEN_18659; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18738 = 5'h4 == T_29096 ? T_38110_4_br_prediction_btb_hit : _GEN_18660; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18739 = 5'h4 == T_29096 ? T_38110_4_br_prediction_btb_predicted : _GEN_18661; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18740 = 5'h4 == T_29096 ? T_38110_4_br_prediction_is_br_or_jalr : _GEN_18662; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18741 = 5'h4 == T_29096 ? T_38110_4_stat_brjmp_mispredicted : _GEN_18663; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18742 = 5'h4 == T_29096 ? T_38110_4_stat_btb_made_pred : _GEN_18664; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18743 = 5'h4 == T_29096 ? T_38110_4_stat_btb_mispredicted : _GEN_18665; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18744 = 5'h4 == T_29096 ? T_38110_4_stat_bpd_made_pred : _GEN_18666; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18745 = 5'h4 == T_29096 ? T_38110_4_stat_bpd_mispredicted : _GEN_18667; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18746 = 5'h4 == T_29096 ? T_38110_4_fetch_pc_lob : _GEN_18668; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18747 = 5'h4 == T_29096 ? T_38110_4_imm_packed : _GEN_18669; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18748 = 5'h4 == T_29096 ? T_38110_4_csr_addr : _GEN_18670; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18749 = 5'h4 == T_29096 ? T_38110_4_rob_idx : _GEN_18671; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18750 = 5'h4 == T_29096 ? T_38110_4_ldq_idx : _GEN_18672; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18751 = 5'h4 == T_29096 ? T_38110_4_stq_idx : _GEN_18673; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18752 = 5'h4 == T_29096 ? T_38110_4_brob_idx : _GEN_18674; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18753 = 5'h4 == T_29096 ? T_38110_4_pdst : _GEN_18675; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18754 = 5'h4 == T_29096 ? T_38110_4_pop1 : _GEN_18676; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18755 = 5'h4 == T_29096 ? T_38110_4_pop2 : _GEN_18677; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18756 = 5'h4 == T_29096 ? T_38110_4_pop3 : _GEN_18678; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18757 = 5'h4 == T_29096 ? T_38110_4_prs1_busy : _GEN_18679; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18758 = 5'h4 == T_29096 ? T_38110_4_prs2_busy : _GEN_18680; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18759 = 5'h4 == T_29096 ? T_38110_4_prs3_busy : _GEN_18681; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18760 = 5'h4 == T_29096 ? T_38110_4_stale_pdst : _GEN_18682; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18761 = 5'h4 == T_29096 ? T_38110_4_exception : _GEN_18683; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18762 = 5'h4 == T_29096 ? T_38110_4_exc_cause : _GEN_18684; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18763 = 5'h4 == T_29096 ? T_38110_4_bypassable : _GEN_18685; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18764 = 5'h4 == T_29096 ? T_38110_4_mem_cmd : _GEN_18686; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18765 = 5'h4 == T_29096 ? T_38110_4_mem_typ : _GEN_18687; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18766 = 5'h4 == T_29096 ? T_38110_4_is_fence : _GEN_18688; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18767 = 5'h4 == T_29096 ? T_38110_4_is_fencei : _GEN_18689; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18768 = 5'h4 == T_29096 ? T_38110_4_is_store : _GEN_18690; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18769 = 5'h4 == T_29096 ? T_38110_4_is_amo : _GEN_18691; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18770 = 5'h4 == T_29096 ? T_38110_4_is_load : _GEN_18692; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18771 = 5'h4 == T_29096 ? T_38110_4_is_unique : _GEN_18693; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18772 = 5'h4 == T_29096 ? T_38110_4_flush_on_commit : _GEN_18694; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18773 = 5'h4 == T_29096 ? T_38110_4_ldst : _GEN_18695; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18774 = 5'h4 == T_29096 ? T_38110_4_lrs1 : _GEN_18696; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18775 = 5'h4 == T_29096 ? T_38110_4_lrs2 : _GEN_18697; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18776 = 5'h4 == T_29096 ? T_38110_4_lrs3 : _GEN_18698; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18777 = 5'h4 == T_29096 ? T_38110_4_ldst_val : _GEN_18699; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18778 = 5'h4 == T_29096 ? T_38110_4_dst_rtype : _GEN_18700; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18779 = 5'h4 == T_29096 ? T_38110_4_lrs1_rtype : _GEN_18701; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18780 = 5'h4 == T_29096 ? T_38110_4_lrs2_rtype : _GEN_18702; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18781 = 5'h4 == T_29096 ? T_38110_4_frs3_en : _GEN_18703; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18782 = 5'h4 == T_29096 ? T_38110_4_fp_val : _GEN_18704; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18783 = 5'h4 == T_29096 ? T_38110_4_fp_single : _GEN_18705; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18784 = 5'h4 == T_29096 ? T_38110_4_xcpt_if : _GEN_18706; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18785 = 5'h4 == T_29096 ? T_38110_4_replay_if : _GEN_18707; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18787 = 5'h4 == T_29096 ? T_38110_4_debug_events_fetch_seq : _GEN_18709; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18788 = 5'h5 == T_29096 ? T_38110_5_valid : _GEN_18710; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18789 = 5'h5 == T_29096 ? T_38110_5_iw_state : _GEN_18711; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18790 = 5'h5 == T_29096 ? T_38110_5_uopc : _GEN_18712; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18791 = 5'h5 == T_29096 ? T_38110_5_inst : _GEN_18713; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18792 = 5'h5 == T_29096 ? T_38110_5_pc : _GEN_18714; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18793 = 5'h5 == T_29096 ? T_38110_5_fu_code : _GEN_18715; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18794 = 5'h5 == T_29096 ? T_38110_5_ctrl_br_type : _GEN_18716; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18795 = 5'h5 == T_29096 ? T_38110_5_ctrl_op1_sel : _GEN_18717; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18796 = 5'h5 == T_29096 ? T_38110_5_ctrl_op2_sel : _GEN_18718; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18797 = 5'h5 == T_29096 ? T_38110_5_ctrl_imm_sel : _GEN_18719; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18798 = 5'h5 == T_29096 ? T_38110_5_ctrl_op_fcn : _GEN_18720; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18799 = 5'h5 == T_29096 ? T_38110_5_ctrl_fcn_dw : _GEN_18721; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18800 = 5'h5 == T_29096 ? T_38110_5_ctrl_rf_wen : _GEN_18722; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18801 = 5'h5 == T_29096 ? T_38110_5_ctrl_csr_cmd : _GEN_18723; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18802 = 5'h5 == T_29096 ? T_38110_5_ctrl_is_load : _GEN_18724; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18803 = 5'h5 == T_29096 ? T_38110_5_ctrl_is_sta : _GEN_18725; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18804 = 5'h5 == T_29096 ? T_38110_5_ctrl_is_std : _GEN_18726; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18805 = 5'h5 == T_29096 ? T_38110_5_wakeup_delay : _GEN_18727; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18806 = 5'h5 == T_29096 ? T_38110_5_allocate_brtag : _GEN_18728; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18807 = 5'h5 == T_29096 ? T_38110_5_is_br_or_jmp : _GEN_18729; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18808 = 5'h5 == T_29096 ? T_38110_5_is_jump : _GEN_18730; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18809 = 5'h5 == T_29096 ? T_38110_5_is_jal : _GEN_18731; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18810 = 5'h5 == T_29096 ? T_38110_5_is_ret : _GEN_18732; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18811 = 5'h5 == T_29096 ? T_38110_5_is_call : _GEN_18733; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18812 = 5'h5 == T_29096 ? T_38110_5_br_mask : _GEN_18734; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18813 = 5'h5 == T_29096 ? T_38110_5_br_tag : _GEN_18735; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18814 = 5'h5 == T_29096 ? T_38110_5_br_prediction_bpd_predict_val : _GEN_18736; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18815 = 5'h5 == T_29096 ? T_38110_5_br_prediction_bpd_predict_taken : _GEN_18737; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18816 = 5'h5 == T_29096 ? T_38110_5_br_prediction_btb_hit : _GEN_18738; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18817 = 5'h5 == T_29096 ? T_38110_5_br_prediction_btb_predicted : _GEN_18739; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18818 = 5'h5 == T_29096 ? T_38110_5_br_prediction_is_br_or_jalr : _GEN_18740; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18819 = 5'h5 == T_29096 ? T_38110_5_stat_brjmp_mispredicted : _GEN_18741; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18820 = 5'h5 == T_29096 ? T_38110_5_stat_btb_made_pred : _GEN_18742; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18821 = 5'h5 == T_29096 ? T_38110_5_stat_btb_mispredicted : _GEN_18743; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18822 = 5'h5 == T_29096 ? T_38110_5_stat_bpd_made_pred : _GEN_18744; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18823 = 5'h5 == T_29096 ? T_38110_5_stat_bpd_mispredicted : _GEN_18745; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18824 = 5'h5 == T_29096 ? T_38110_5_fetch_pc_lob : _GEN_18746; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18825 = 5'h5 == T_29096 ? T_38110_5_imm_packed : _GEN_18747; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18826 = 5'h5 == T_29096 ? T_38110_5_csr_addr : _GEN_18748; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18827 = 5'h5 == T_29096 ? T_38110_5_rob_idx : _GEN_18749; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18828 = 5'h5 == T_29096 ? T_38110_5_ldq_idx : _GEN_18750; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18829 = 5'h5 == T_29096 ? T_38110_5_stq_idx : _GEN_18751; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18830 = 5'h5 == T_29096 ? T_38110_5_brob_idx : _GEN_18752; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18831 = 5'h5 == T_29096 ? T_38110_5_pdst : _GEN_18753; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18832 = 5'h5 == T_29096 ? T_38110_5_pop1 : _GEN_18754; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18833 = 5'h5 == T_29096 ? T_38110_5_pop2 : _GEN_18755; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18834 = 5'h5 == T_29096 ? T_38110_5_pop3 : _GEN_18756; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18835 = 5'h5 == T_29096 ? T_38110_5_prs1_busy : _GEN_18757; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18836 = 5'h5 == T_29096 ? T_38110_5_prs2_busy : _GEN_18758; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18837 = 5'h5 == T_29096 ? T_38110_5_prs3_busy : _GEN_18759; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18838 = 5'h5 == T_29096 ? T_38110_5_stale_pdst : _GEN_18760; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18839 = 5'h5 == T_29096 ? T_38110_5_exception : _GEN_18761; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18840 = 5'h5 == T_29096 ? T_38110_5_exc_cause : _GEN_18762; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18841 = 5'h5 == T_29096 ? T_38110_5_bypassable : _GEN_18763; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18842 = 5'h5 == T_29096 ? T_38110_5_mem_cmd : _GEN_18764; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18843 = 5'h5 == T_29096 ? T_38110_5_mem_typ : _GEN_18765; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18844 = 5'h5 == T_29096 ? T_38110_5_is_fence : _GEN_18766; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18845 = 5'h5 == T_29096 ? T_38110_5_is_fencei : _GEN_18767; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18846 = 5'h5 == T_29096 ? T_38110_5_is_store : _GEN_18768; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18847 = 5'h5 == T_29096 ? T_38110_5_is_amo : _GEN_18769; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18848 = 5'h5 == T_29096 ? T_38110_5_is_load : _GEN_18770; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18849 = 5'h5 == T_29096 ? T_38110_5_is_unique : _GEN_18771; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18850 = 5'h5 == T_29096 ? T_38110_5_flush_on_commit : _GEN_18772; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18851 = 5'h5 == T_29096 ? T_38110_5_ldst : _GEN_18773; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18852 = 5'h5 == T_29096 ? T_38110_5_lrs1 : _GEN_18774; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18853 = 5'h5 == T_29096 ? T_38110_5_lrs2 : _GEN_18775; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18854 = 5'h5 == T_29096 ? T_38110_5_lrs3 : _GEN_18776; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18855 = 5'h5 == T_29096 ? T_38110_5_ldst_val : _GEN_18777; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18856 = 5'h5 == T_29096 ? T_38110_5_dst_rtype : _GEN_18778; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18857 = 5'h5 == T_29096 ? T_38110_5_lrs1_rtype : _GEN_18779; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18858 = 5'h5 == T_29096 ? T_38110_5_lrs2_rtype : _GEN_18780; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18859 = 5'h5 == T_29096 ? T_38110_5_frs3_en : _GEN_18781; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18860 = 5'h5 == T_29096 ? T_38110_5_fp_val : _GEN_18782; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18861 = 5'h5 == T_29096 ? T_38110_5_fp_single : _GEN_18783; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18862 = 5'h5 == T_29096 ? T_38110_5_xcpt_if : _GEN_18784; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18863 = 5'h5 == T_29096 ? T_38110_5_replay_if : _GEN_18785; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18865 = 5'h5 == T_29096 ? T_38110_5_debug_events_fetch_seq : _GEN_18787; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18866 = 5'h6 == T_29096 ? T_38110_6_valid : _GEN_18788; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18867 = 5'h6 == T_29096 ? T_38110_6_iw_state : _GEN_18789; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18868 = 5'h6 == T_29096 ? T_38110_6_uopc : _GEN_18790; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18869 = 5'h6 == T_29096 ? T_38110_6_inst : _GEN_18791; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18870 = 5'h6 == T_29096 ? T_38110_6_pc : _GEN_18792; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18871 = 5'h6 == T_29096 ? T_38110_6_fu_code : _GEN_18793; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18872 = 5'h6 == T_29096 ? T_38110_6_ctrl_br_type : _GEN_18794; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18873 = 5'h6 == T_29096 ? T_38110_6_ctrl_op1_sel : _GEN_18795; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18874 = 5'h6 == T_29096 ? T_38110_6_ctrl_op2_sel : _GEN_18796; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18875 = 5'h6 == T_29096 ? T_38110_6_ctrl_imm_sel : _GEN_18797; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18876 = 5'h6 == T_29096 ? T_38110_6_ctrl_op_fcn : _GEN_18798; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18877 = 5'h6 == T_29096 ? T_38110_6_ctrl_fcn_dw : _GEN_18799; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18878 = 5'h6 == T_29096 ? T_38110_6_ctrl_rf_wen : _GEN_18800; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18879 = 5'h6 == T_29096 ? T_38110_6_ctrl_csr_cmd : _GEN_18801; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18880 = 5'h6 == T_29096 ? T_38110_6_ctrl_is_load : _GEN_18802; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18881 = 5'h6 == T_29096 ? T_38110_6_ctrl_is_sta : _GEN_18803; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18882 = 5'h6 == T_29096 ? T_38110_6_ctrl_is_std : _GEN_18804; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18883 = 5'h6 == T_29096 ? T_38110_6_wakeup_delay : _GEN_18805; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18884 = 5'h6 == T_29096 ? T_38110_6_allocate_brtag : _GEN_18806; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18885 = 5'h6 == T_29096 ? T_38110_6_is_br_or_jmp : _GEN_18807; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18886 = 5'h6 == T_29096 ? T_38110_6_is_jump : _GEN_18808; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18887 = 5'h6 == T_29096 ? T_38110_6_is_jal : _GEN_18809; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18888 = 5'h6 == T_29096 ? T_38110_6_is_ret : _GEN_18810; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18889 = 5'h6 == T_29096 ? T_38110_6_is_call : _GEN_18811; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18890 = 5'h6 == T_29096 ? T_38110_6_br_mask : _GEN_18812; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18891 = 5'h6 == T_29096 ? T_38110_6_br_tag : _GEN_18813; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18892 = 5'h6 == T_29096 ? T_38110_6_br_prediction_bpd_predict_val : _GEN_18814; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18893 = 5'h6 == T_29096 ? T_38110_6_br_prediction_bpd_predict_taken : _GEN_18815; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18894 = 5'h6 == T_29096 ? T_38110_6_br_prediction_btb_hit : _GEN_18816; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18895 = 5'h6 == T_29096 ? T_38110_6_br_prediction_btb_predicted : _GEN_18817; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18896 = 5'h6 == T_29096 ? T_38110_6_br_prediction_is_br_or_jalr : _GEN_18818; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18897 = 5'h6 == T_29096 ? T_38110_6_stat_brjmp_mispredicted : _GEN_18819; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18898 = 5'h6 == T_29096 ? T_38110_6_stat_btb_made_pred : _GEN_18820; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18899 = 5'h6 == T_29096 ? T_38110_6_stat_btb_mispredicted : _GEN_18821; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18900 = 5'h6 == T_29096 ? T_38110_6_stat_bpd_made_pred : _GEN_18822; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18901 = 5'h6 == T_29096 ? T_38110_6_stat_bpd_mispredicted : _GEN_18823; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18902 = 5'h6 == T_29096 ? T_38110_6_fetch_pc_lob : _GEN_18824; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18903 = 5'h6 == T_29096 ? T_38110_6_imm_packed : _GEN_18825; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18904 = 5'h6 == T_29096 ? T_38110_6_csr_addr : _GEN_18826; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18905 = 5'h6 == T_29096 ? T_38110_6_rob_idx : _GEN_18827; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18906 = 5'h6 == T_29096 ? T_38110_6_ldq_idx : _GEN_18828; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18907 = 5'h6 == T_29096 ? T_38110_6_stq_idx : _GEN_18829; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18908 = 5'h6 == T_29096 ? T_38110_6_brob_idx : _GEN_18830; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18909 = 5'h6 == T_29096 ? T_38110_6_pdst : _GEN_18831; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18910 = 5'h6 == T_29096 ? T_38110_6_pop1 : _GEN_18832; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18911 = 5'h6 == T_29096 ? T_38110_6_pop2 : _GEN_18833; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18912 = 5'h6 == T_29096 ? T_38110_6_pop3 : _GEN_18834; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18913 = 5'h6 == T_29096 ? T_38110_6_prs1_busy : _GEN_18835; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18914 = 5'h6 == T_29096 ? T_38110_6_prs2_busy : _GEN_18836; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18915 = 5'h6 == T_29096 ? T_38110_6_prs3_busy : _GEN_18837; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18916 = 5'h6 == T_29096 ? T_38110_6_stale_pdst : _GEN_18838; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18917 = 5'h6 == T_29096 ? T_38110_6_exception : _GEN_18839; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18918 = 5'h6 == T_29096 ? T_38110_6_exc_cause : _GEN_18840; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18919 = 5'h6 == T_29096 ? T_38110_6_bypassable : _GEN_18841; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18920 = 5'h6 == T_29096 ? T_38110_6_mem_cmd : _GEN_18842; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18921 = 5'h6 == T_29096 ? T_38110_6_mem_typ : _GEN_18843; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18922 = 5'h6 == T_29096 ? T_38110_6_is_fence : _GEN_18844; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18923 = 5'h6 == T_29096 ? T_38110_6_is_fencei : _GEN_18845; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18924 = 5'h6 == T_29096 ? T_38110_6_is_store : _GEN_18846; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18925 = 5'h6 == T_29096 ? T_38110_6_is_amo : _GEN_18847; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18926 = 5'h6 == T_29096 ? T_38110_6_is_load : _GEN_18848; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18927 = 5'h6 == T_29096 ? T_38110_6_is_unique : _GEN_18849; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18928 = 5'h6 == T_29096 ? T_38110_6_flush_on_commit : _GEN_18850; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18929 = 5'h6 == T_29096 ? T_38110_6_ldst : _GEN_18851; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18930 = 5'h6 == T_29096 ? T_38110_6_lrs1 : _GEN_18852; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18931 = 5'h6 == T_29096 ? T_38110_6_lrs2 : _GEN_18853; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18932 = 5'h6 == T_29096 ? T_38110_6_lrs3 : _GEN_18854; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18933 = 5'h6 == T_29096 ? T_38110_6_ldst_val : _GEN_18855; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18934 = 5'h6 == T_29096 ? T_38110_6_dst_rtype : _GEN_18856; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18935 = 5'h6 == T_29096 ? T_38110_6_lrs1_rtype : _GEN_18857; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18936 = 5'h6 == T_29096 ? T_38110_6_lrs2_rtype : _GEN_18858; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18937 = 5'h6 == T_29096 ? T_38110_6_frs3_en : _GEN_18859; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18938 = 5'h6 == T_29096 ? T_38110_6_fp_val : _GEN_18860; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18939 = 5'h6 == T_29096 ? T_38110_6_fp_single : _GEN_18861; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18940 = 5'h6 == T_29096 ? T_38110_6_xcpt_if : _GEN_18862; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18941 = 5'h6 == T_29096 ? T_38110_6_replay_if : _GEN_18863; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18943 = 5'h6 == T_29096 ? T_38110_6_debug_events_fetch_seq : _GEN_18865; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18944 = 5'h7 == T_29096 ? T_38110_7_valid : _GEN_18866; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18945 = 5'h7 == T_29096 ? T_38110_7_iw_state : _GEN_18867; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_18946 = 5'h7 == T_29096 ? T_38110_7_uopc : _GEN_18868; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_18947 = 5'h7 == T_29096 ? T_38110_7_inst : _GEN_18869; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_18948 = 5'h7 == T_29096 ? T_38110_7_pc : _GEN_18870; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18949 = 5'h7 == T_29096 ? T_38110_7_fu_code : _GEN_18871; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18950 = 5'h7 == T_29096 ? T_38110_7_ctrl_br_type : _GEN_18872; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18951 = 5'h7 == T_29096 ? T_38110_7_ctrl_op1_sel : _GEN_18873; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18952 = 5'h7 == T_29096 ? T_38110_7_ctrl_op2_sel : _GEN_18874; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18953 = 5'h7 == T_29096 ? T_38110_7_ctrl_imm_sel : _GEN_18875; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18954 = 5'h7 == T_29096 ? T_38110_7_ctrl_op_fcn : _GEN_18876; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18955 = 5'h7 == T_29096 ? T_38110_7_ctrl_fcn_dw : _GEN_18877; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18956 = 5'h7 == T_29096 ? T_38110_7_ctrl_rf_wen : _GEN_18878; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18957 = 5'h7 == T_29096 ? T_38110_7_ctrl_csr_cmd : _GEN_18879; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18958 = 5'h7 == T_29096 ? T_38110_7_ctrl_is_load : _GEN_18880; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18959 = 5'h7 == T_29096 ? T_38110_7_ctrl_is_sta : _GEN_18881; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18960 = 5'h7 == T_29096 ? T_38110_7_ctrl_is_std : _GEN_18882; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_18961 = 5'h7 == T_29096 ? T_38110_7_wakeup_delay : _GEN_18883; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18962 = 5'h7 == T_29096 ? T_38110_7_allocate_brtag : _GEN_18884; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18963 = 5'h7 == T_29096 ? T_38110_7_is_br_or_jmp : _GEN_18885; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18964 = 5'h7 == T_29096 ? T_38110_7_is_jump : _GEN_18886; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18965 = 5'h7 == T_29096 ? T_38110_7_is_jal : _GEN_18887; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18966 = 5'h7 == T_29096 ? T_38110_7_is_ret : _GEN_18888; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18967 = 5'h7 == T_29096 ? T_38110_7_is_call : _GEN_18889; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_18968 = 5'h7 == T_29096 ? T_38110_7_br_mask : _GEN_18890; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18969 = 5'h7 == T_29096 ? T_38110_7_br_tag : _GEN_18891; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18970 = 5'h7 == T_29096 ? T_38110_7_br_prediction_bpd_predict_val : _GEN_18892; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18971 = 5'h7 == T_29096 ? T_38110_7_br_prediction_bpd_predict_taken : _GEN_18893; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18972 = 5'h7 == T_29096 ? T_38110_7_br_prediction_btb_hit : _GEN_18894; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18973 = 5'h7 == T_29096 ? T_38110_7_br_prediction_btb_predicted : _GEN_18895; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18974 = 5'h7 == T_29096 ? T_38110_7_br_prediction_is_br_or_jalr : _GEN_18896; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18975 = 5'h7 == T_29096 ? T_38110_7_stat_brjmp_mispredicted : _GEN_18897; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18976 = 5'h7 == T_29096 ? T_38110_7_stat_btb_made_pred : _GEN_18898; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18977 = 5'h7 == T_29096 ? T_38110_7_stat_btb_mispredicted : _GEN_18899; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18978 = 5'h7 == T_29096 ? T_38110_7_stat_bpd_made_pred : _GEN_18900; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18979 = 5'h7 == T_29096 ? T_38110_7_stat_bpd_mispredicted : _GEN_18901; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18980 = 5'h7 == T_29096 ? T_38110_7_fetch_pc_lob : _GEN_18902; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_18981 = 5'h7 == T_29096 ? T_38110_7_imm_packed : _GEN_18903; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_18982 = 5'h7 == T_29096 ? T_38110_7_csr_addr : _GEN_18904; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_18983 = 5'h7 == T_29096 ? T_38110_7_rob_idx : _GEN_18905; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18984 = 5'h7 == T_29096 ? T_38110_7_ldq_idx : _GEN_18906; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18985 = 5'h7 == T_29096 ? T_38110_7_stq_idx : _GEN_18907; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_18986 = 5'h7 == T_29096 ? T_38110_7_brob_idx : _GEN_18908; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18987 = 5'h7 == T_29096 ? T_38110_7_pdst : _GEN_18909; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18988 = 5'h7 == T_29096 ? T_38110_7_pop1 : _GEN_18910; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18989 = 5'h7 == T_29096 ? T_38110_7_pop2 : _GEN_18911; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18990 = 5'h7 == T_29096 ? T_38110_7_pop3 : _GEN_18912; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18991 = 5'h7 == T_29096 ? T_38110_7_prs1_busy : _GEN_18913; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18992 = 5'h7 == T_29096 ? T_38110_7_prs2_busy : _GEN_18914; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18993 = 5'h7 == T_29096 ? T_38110_7_prs3_busy : _GEN_18915; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_18994 = 5'h7 == T_29096 ? T_38110_7_stale_pdst : _GEN_18916; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18995 = 5'h7 == T_29096 ? T_38110_7_exception : _GEN_18917; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_18996 = 5'h7 == T_29096 ? T_38110_7_exc_cause : _GEN_18918; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_18997 = 5'h7 == T_29096 ? T_38110_7_bypassable : _GEN_18919; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_18998 = 5'h7 == T_29096 ? T_38110_7_mem_cmd : _GEN_18920; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_18999 = 5'h7 == T_29096 ? T_38110_7_mem_typ : _GEN_18921; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19000 = 5'h7 == T_29096 ? T_38110_7_is_fence : _GEN_18922; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19001 = 5'h7 == T_29096 ? T_38110_7_is_fencei : _GEN_18923; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19002 = 5'h7 == T_29096 ? T_38110_7_is_store : _GEN_18924; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19003 = 5'h7 == T_29096 ? T_38110_7_is_amo : _GEN_18925; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19004 = 5'h7 == T_29096 ? T_38110_7_is_load : _GEN_18926; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19005 = 5'h7 == T_29096 ? T_38110_7_is_unique : _GEN_18927; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19006 = 5'h7 == T_29096 ? T_38110_7_flush_on_commit : _GEN_18928; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19007 = 5'h7 == T_29096 ? T_38110_7_ldst : _GEN_18929; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19008 = 5'h7 == T_29096 ? T_38110_7_lrs1 : _GEN_18930; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19009 = 5'h7 == T_29096 ? T_38110_7_lrs2 : _GEN_18931; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19010 = 5'h7 == T_29096 ? T_38110_7_lrs3 : _GEN_18932; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19011 = 5'h7 == T_29096 ? T_38110_7_ldst_val : _GEN_18933; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19012 = 5'h7 == T_29096 ? T_38110_7_dst_rtype : _GEN_18934; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19013 = 5'h7 == T_29096 ? T_38110_7_lrs1_rtype : _GEN_18935; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19014 = 5'h7 == T_29096 ? T_38110_7_lrs2_rtype : _GEN_18936; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19015 = 5'h7 == T_29096 ? T_38110_7_frs3_en : _GEN_18937; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19016 = 5'h7 == T_29096 ? T_38110_7_fp_val : _GEN_18938; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19017 = 5'h7 == T_29096 ? T_38110_7_fp_single : _GEN_18939; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19018 = 5'h7 == T_29096 ? T_38110_7_xcpt_if : _GEN_18940; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19019 = 5'h7 == T_29096 ? T_38110_7_replay_if : _GEN_18941; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19021 = 5'h7 == T_29096 ? T_38110_7_debug_events_fetch_seq : _GEN_18943; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19022 = 5'h8 == T_29096 ? T_38110_8_valid : _GEN_18944; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19023 = 5'h8 == T_29096 ? T_38110_8_iw_state : _GEN_18945; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19024 = 5'h8 == T_29096 ? T_38110_8_uopc : _GEN_18946; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19025 = 5'h8 == T_29096 ? T_38110_8_inst : _GEN_18947; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19026 = 5'h8 == T_29096 ? T_38110_8_pc : _GEN_18948; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19027 = 5'h8 == T_29096 ? T_38110_8_fu_code : _GEN_18949; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19028 = 5'h8 == T_29096 ? T_38110_8_ctrl_br_type : _GEN_18950; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19029 = 5'h8 == T_29096 ? T_38110_8_ctrl_op1_sel : _GEN_18951; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19030 = 5'h8 == T_29096 ? T_38110_8_ctrl_op2_sel : _GEN_18952; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19031 = 5'h8 == T_29096 ? T_38110_8_ctrl_imm_sel : _GEN_18953; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19032 = 5'h8 == T_29096 ? T_38110_8_ctrl_op_fcn : _GEN_18954; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19033 = 5'h8 == T_29096 ? T_38110_8_ctrl_fcn_dw : _GEN_18955; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19034 = 5'h8 == T_29096 ? T_38110_8_ctrl_rf_wen : _GEN_18956; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19035 = 5'h8 == T_29096 ? T_38110_8_ctrl_csr_cmd : _GEN_18957; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19036 = 5'h8 == T_29096 ? T_38110_8_ctrl_is_load : _GEN_18958; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19037 = 5'h8 == T_29096 ? T_38110_8_ctrl_is_sta : _GEN_18959; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19038 = 5'h8 == T_29096 ? T_38110_8_ctrl_is_std : _GEN_18960; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19039 = 5'h8 == T_29096 ? T_38110_8_wakeup_delay : _GEN_18961; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19040 = 5'h8 == T_29096 ? T_38110_8_allocate_brtag : _GEN_18962; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19041 = 5'h8 == T_29096 ? T_38110_8_is_br_or_jmp : _GEN_18963; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19042 = 5'h8 == T_29096 ? T_38110_8_is_jump : _GEN_18964; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19043 = 5'h8 == T_29096 ? T_38110_8_is_jal : _GEN_18965; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19044 = 5'h8 == T_29096 ? T_38110_8_is_ret : _GEN_18966; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19045 = 5'h8 == T_29096 ? T_38110_8_is_call : _GEN_18967; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19046 = 5'h8 == T_29096 ? T_38110_8_br_mask : _GEN_18968; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19047 = 5'h8 == T_29096 ? T_38110_8_br_tag : _GEN_18969; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19048 = 5'h8 == T_29096 ? T_38110_8_br_prediction_bpd_predict_val : _GEN_18970; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19049 = 5'h8 == T_29096 ? T_38110_8_br_prediction_bpd_predict_taken : _GEN_18971; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19050 = 5'h8 == T_29096 ? T_38110_8_br_prediction_btb_hit : _GEN_18972; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19051 = 5'h8 == T_29096 ? T_38110_8_br_prediction_btb_predicted : _GEN_18973; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19052 = 5'h8 == T_29096 ? T_38110_8_br_prediction_is_br_or_jalr : _GEN_18974; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19053 = 5'h8 == T_29096 ? T_38110_8_stat_brjmp_mispredicted : _GEN_18975; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19054 = 5'h8 == T_29096 ? T_38110_8_stat_btb_made_pred : _GEN_18976; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19055 = 5'h8 == T_29096 ? T_38110_8_stat_btb_mispredicted : _GEN_18977; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19056 = 5'h8 == T_29096 ? T_38110_8_stat_bpd_made_pred : _GEN_18978; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19057 = 5'h8 == T_29096 ? T_38110_8_stat_bpd_mispredicted : _GEN_18979; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19058 = 5'h8 == T_29096 ? T_38110_8_fetch_pc_lob : _GEN_18980; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19059 = 5'h8 == T_29096 ? T_38110_8_imm_packed : _GEN_18981; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19060 = 5'h8 == T_29096 ? T_38110_8_csr_addr : _GEN_18982; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19061 = 5'h8 == T_29096 ? T_38110_8_rob_idx : _GEN_18983; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19062 = 5'h8 == T_29096 ? T_38110_8_ldq_idx : _GEN_18984; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19063 = 5'h8 == T_29096 ? T_38110_8_stq_idx : _GEN_18985; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19064 = 5'h8 == T_29096 ? T_38110_8_brob_idx : _GEN_18986; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19065 = 5'h8 == T_29096 ? T_38110_8_pdst : _GEN_18987; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19066 = 5'h8 == T_29096 ? T_38110_8_pop1 : _GEN_18988; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19067 = 5'h8 == T_29096 ? T_38110_8_pop2 : _GEN_18989; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19068 = 5'h8 == T_29096 ? T_38110_8_pop3 : _GEN_18990; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19069 = 5'h8 == T_29096 ? T_38110_8_prs1_busy : _GEN_18991; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19070 = 5'h8 == T_29096 ? T_38110_8_prs2_busy : _GEN_18992; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19071 = 5'h8 == T_29096 ? T_38110_8_prs3_busy : _GEN_18993; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19072 = 5'h8 == T_29096 ? T_38110_8_stale_pdst : _GEN_18994; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19073 = 5'h8 == T_29096 ? T_38110_8_exception : _GEN_18995; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19074 = 5'h8 == T_29096 ? T_38110_8_exc_cause : _GEN_18996; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19075 = 5'h8 == T_29096 ? T_38110_8_bypassable : _GEN_18997; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19076 = 5'h8 == T_29096 ? T_38110_8_mem_cmd : _GEN_18998; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19077 = 5'h8 == T_29096 ? T_38110_8_mem_typ : _GEN_18999; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19078 = 5'h8 == T_29096 ? T_38110_8_is_fence : _GEN_19000; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19079 = 5'h8 == T_29096 ? T_38110_8_is_fencei : _GEN_19001; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19080 = 5'h8 == T_29096 ? T_38110_8_is_store : _GEN_19002; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19081 = 5'h8 == T_29096 ? T_38110_8_is_amo : _GEN_19003; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19082 = 5'h8 == T_29096 ? T_38110_8_is_load : _GEN_19004; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19083 = 5'h8 == T_29096 ? T_38110_8_is_unique : _GEN_19005; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19084 = 5'h8 == T_29096 ? T_38110_8_flush_on_commit : _GEN_19006; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19085 = 5'h8 == T_29096 ? T_38110_8_ldst : _GEN_19007; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19086 = 5'h8 == T_29096 ? T_38110_8_lrs1 : _GEN_19008; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19087 = 5'h8 == T_29096 ? T_38110_8_lrs2 : _GEN_19009; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19088 = 5'h8 == T_29096 ? T_38110_8_lrs3 : _GEN_19010; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19089 = 5'h8 == T_29096 ? T_38110_8_ldst_val : _GEN_19011; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19090 = 5'h8 == T_29096 ? T_38110_8_dst_rtype : _GEN_19012; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19091 = 5'h8 == T_29096 ? T_38110_8_lrs1_rtype : _GEN_19013; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19092 = 5'h8 == T_29096 ? T_38110_8_lrs2_rtype : _GEN_19014; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19093 = 5'h8 == T_29096 ? T_38110_8_frs3_en : _GEN_19015; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19094 = 5'h8 == T_29096 ? T_38110_8_fp_val : _GEN_19016; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19095 = 5'h8 == T_29096 ? T_38110_8_fp_single : _GEN_19017; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19096 = 5'h8 == T_29096 ? T_38110_8_xcpt_if : _GEN_19018; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19097 = 5'h8 == T_29096 ? T_38110_8_replay_if : _GEN_19019; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19099 = 5'h8 == T_29096 ? T_38110_8_debug_events_fetch_seq : _GEN_19021; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19100 = 5'h9 == T_29096 ? T_38110_9_valid : _GEN_19022; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19101 = 5'h9 == T_29096 ? T_38110_9_iw_state : _GEN_19023; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19102 = 5'h9 == T_29096 ? T_38110_9_uopc : _GEN_19024; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19103 = 5'h9 == T_29096 ? T_38110_9_inst : _GEN_19025; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19104 = 5'h9 == T_29096 ? T_38110_9_pc : _GEN_19026; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19105 = 5'h9 == T_29096 ? T_38110_9_fu_code : _GEN_19027; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19106 = 5'h9 == T_29096 ? T_38110_9_ctrl_br_type : _GEN_19028; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19107 = 5'h9 == T_29096 ? T_38110_9_ctrl_op1_sel : _GEN_19029; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19108 = 5'h9 == T_29096 ? T_38110_9_ctrl_op2_sel : _GEN_19030; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19109 = 5'h9 == T_29096 ? T_38110_9_ctrl_imm_sel : _GEN_19031; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19110 = 5'h9 == T_29096 ? T_38110_9_ctrl_op_fcn : _GEN_19032; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19111 = 5'h9 == T_29096 ? T_38110_9_ctrl_fcn_dw : _GEN_19033; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19112 = 5'h9 == T_29096 ? T_38110_9_ctrl_rf_wen : _GEN_19034; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19113 = 5'h9 == T_29096 ? T_38110_9_ctrl_csr_cmd : _GEN_19035; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19114 = 5'h9 == T_29096 ? T_38110_9_ctrl_is_load : _GEN_19036; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19115 = 5'h9 == T_29096 ? T_38110_9_ctrl_is_sta : _GEN_19037; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19116 = 5'h9 == T_29096 ? T_38110_9_ctrl_is_std : _GEN_19038; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19117 = 5'h9 == T_29096 ? T_38110_9_wakeup_delay : _GEN_19039; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19118 = 5'h9 == T_29096 ? T_38110_9_allocate_brtag : _GEN_19040; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19119 = 5'h9 == T_29096 ? T_38110_9_is_br_or_jmp : _GEN_19041; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19120 = 5'h9 == T_29096 ? T_38110_9_is_jump : _GEN_19042; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19121 = 5'h9 == T_29096 ? T_38110_9_is_jal : _GEN_19043; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19122 = 5'h9 == T_29096 ? T_38110_9_is_ret : _GEN_19044; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19123 = 5'h9 == T_29096 ? T_38110_9_is_call : _GEN_19045; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19124 = 5'h9 == T_29096 ? T_38110_9_br_mask : _GEN_19046; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19125 = 5'h9 == T_29096 ? T_38110_9_br_tag : _GEN_19047; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19126 = 5'h9 == T_29096 ? T_38110_9_br_prediction_bpd_predict_val : _GEN_19048; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19127 = 5'h9 == T_29096 ? T_38110_9_br_prediction_bpd_predict_taken : _GEN_19049; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19128 = 5'h9 == T_29096 ? T_38110_9_br_prediction_btb_hit : _GEN_19050; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19129 = 5'h9 == T_29096 ? T_38110_9_br_prediction_btb_predicted : _GEN_19051; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19130 = 5'h9 == T_29096 ? T_38110_9_br_prediction_is_br_or_jalr : _GEN_19052; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19131 = 5'h9 == T_29096 ? T_38110_9_stat_brjmp_mispredicted : _GEN_19053; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19132 = 5'h9 == T_29096 ? T_38110_9_stat_btb_made_pred : _GEN_19054; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19133 = 5'h9 == T_29096 ? T_38110_9_stat_btb_mispredicted : _GEN_19055; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19134 = 5'h9 == T_29096 ? T_38110_9_stat_bpd_made_pred : _GEN_19056; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19135 = 5'h9 == T_29096 ? T_38110_9_stat_bpd_mispredicted : _GEN_19057; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19136 = 5'h9 == T_29096 ? T_38110_9_fetch_pc_lob : _GEN_19058; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19137 = 5'h9 == T_29096 ? T_38110_9_imm_packed : _GEN_19059; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19138 = 5'h9 == T_29096 ? T_38110_9_csr_addr : _GEN_19060; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19139 = 5'h9 == T_29096 ? T_38110_9_rob_idx : _GEN_19061; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19140 = 5'h9 == T_29096 ? T_38110_9_ldq_idx : _GEN_19062; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19141 = 5'h9 == T_29096 ? T_38110_9_stq_idx : _GEN_19063; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19142 = 5'h9 == T_29096 ? T_38110_9_brob_idx : _GEN_19064; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19143 = 5'h9 == T_29096 ? T_38110_9_pdst : _GEN_19065; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19144 = 5'h9 == T_29096 ? T_38110_9_pop1 : _GEN_19066; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19145 = 5'h9 == T_29096 ? T_38110_9_pop2 : _GEN_19067; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19146 = 5'h9 == T_29096 ? T_38110_9_pop3 : _GEN_19068; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19147 = 5'h9 == T_29096 ? T_38110_9_prs1_busy : _GEN_19069; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19148 = 5'h9 == T_29096 ? T_38110_9_prs2_busy : _GEN_19070; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19149 = 5'h9 == T_29096 ? T_38110_9_prs3_busy : _GEN_19071; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19150 = 5'h9 == T_29096 ? T_38110_9_stale_pdst : _GEN_19072; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19151 = 5'h9 == T_29096 ? T_38110_9_exception : _GEN_19073; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19152 = 5'h9 == T_29096 ? T_38110_9_exc_cause : _GEN_19074; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19153 = 5'h9 == T_29096 ? T_38110_9_bypassable : _GEN_19075; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19154 = 5'h9 == T_29096 ? T_38110_9_mem_cmd : _GEN_19076; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19155 = 5'h9 == T_29096 ? T_38110_9_mem_typ : _GEN_19077; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19156 = 5'h9 == T_29096 ? T_38110_9_is_fence : _GEN_19078; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19157 = 5'h9 == T_29096 ? T_38110_9_is_fencei : _GEN_19079; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19158 = 5'h9 == T_29096 ? T_38110_9_is_store : _GEN_19080; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19159 = 5'h9 == T_29096 ? T_38110_9_is_amo : _GEN_19081; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19160 = 5'h9 == T_29096 ? T_38110_9_is_load : _GEN_19082; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19161 = 5'h9 == T_29096 ? T_38110_9_is_unique : _GEN_19083; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19162 = 5'h9 == T_29096 ? T_38110_9_flush_on_commit : _GEN_19084; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19163 = 5'h9 == T_29096 ? T_38110_9_ldst : _GEN_19085; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19164 = 5'h9 == T_29096 ? T_38110_9_lrs1 : _GEN_19086; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19165 = 5'h9 == T_29096 ? T_38110_9_lrs2 : _GEN_19087; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19166 = 5'h9 == T_29096 ? T_38110_9_lrs3 : _GEN_19088; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19167 = 5'h9 == T_29096 ? T_38110_9_ldst_val : _GEN_19089; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19168 = 5'h9 == T_29096 ? T_38110_9_dst_rtype : _GEN_19090; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19169 = 5'h9 == T_29096 ? T_38110_9_lrs1_rtype : _GEN_19091; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19170 = 5'h9 == T_29096 ? T_38110_9_lrs2_rtype : _GEN_19092; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19171 = 5'h9 == T_29096 ? T_38110_9_frs3_en : _GEN_19093; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19172 = 5'h9 == T_29096 ? T_38110_9_fp_val : _GEN_19094; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19173 = 5'h9 == T_29096 ? T_38110_9_fp_single : _GEN_19095; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19174 = 5'h9 == T_29096 ? T_38110_9_xcpt_if : _GEN_19096; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19175 = 5'h9 == T_29096 ? T_38110_9_replay_if : _GEN_19097; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19177 = 5'h9 == T_29096 ? T_38110_9_debug_events_fetch_seq : _GEN_19099; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19178 = 5'ha == T_29096 ? T_38110_10_valid : _GEN_19100; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19179 = 5'ha == T_29096 ? T_38110_10_iw_state : _GEN_19101; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19180 = 5'ha == T_29096 ? T_38110_10_uopc : _GEN_19102; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19181 = 5'ha == T_29096 ? T_38110_10_inst : _GEN_19103; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19182 = 5'ha == T_29096 ? T_38110_10_pc : _GEN_19104; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19183 = 5'ha == T_29096 ? T_38110_10_fu_code : _GEN_19105; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19184 = 5'ha == T_29096 ? T_38110_10_ctrl_br_type : _GEN_19106; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19185 = 5'ha == T_29096 ? T_38110_10_ctrl_op1_sel : _GEN_19107; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19186 = 5'ha == T_29096 ? T_38110_10_ctrl_op2_sel : _GEN_19108; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19187 = 5'ha == T_29096 ? T_38110_10_ctrl_imm_sel : _GEN_19109; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19188 = 5'ha == T_29096 ? T_38110_10_ctrl_op_fcn : _GEN_19110; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19189 = 5'ha == T_29096 ? T_38110_10_ctrl_fcn_dw : _GEN_19111; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19190 = 5'ha == T_29096 ? T_38110_10_ctrl_rf_wen : _GEN_19112; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19191 = 5'ha == T_29096 ? T_38110_10_ctrl_csr_cmd : _GEN_19113; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19192 = 5'ha == T_29096 ? T_38110_10_ctrl_is_load : _GEN_19114; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19193 = 5'ha == T_29096 ? T_38110_10_ctrl_is_sta : _GEN_19115; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19194 = 5'ha == T_29096 ? T_38110_10_ctrl_is_std : _GEN_19116; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19195 = 5'ha == T_29096 ? T_38110_10_wakeup_delay : _GEN_19117; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19196 = 5'ha == T_29096 ? T_38110_10_allocate_brtag : _GEN_19118; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19197 = 5'ha == T_29096 ? T_38110_10_is_br_or_jmp : _GEN_19119; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19198 = 5'ha == T_29096 ? T_38110_10_is_jump : _GEN_19120; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19199 = 5'ha == T_29096 ? T_38110_10_is_jal : _GEN_19121; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19200 = 5'ha == T_29096 ? T_38110_10_is_ret : _GEN_19122; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19201 = 5'ha == T_29096 ? T_38110_10_is_call : _GEN_19123; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19202 = 5'ha == T_29096 ? T_38110_10_br_mask : _GEN_19124; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19203 = 5'ha == T_29096 ? T_38110_10_br_tag : _GEN_19125; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19204 = 5'ha == T_29096 ? T_38110_10_br_prediction_bpd_predict_val : _GEN_19126; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19205 = 5'ha == T_29096 ? T_38110_10_br_prediction_bpd_predict_taken : _GEN_19127; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19206 = 5'ha == T_29096 ? T_38110_10_br_prediction_btb_hit : _GEN_19128; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19207 = 5'ha == T_29096 ? T_38110_10_br_prediction_btb_predicted : _GEN_19129; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19208 = 5'ha == T_29096 ? T_38110_10_br_prediction_is_br_or_jalr : _GEN_19130; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19209 = 5'ha == T_29096 ? T_38110_10_stat_brjmp_mispredicted : _GEN_19131; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19210 = 5'ha == T_29096 ? T_38110_10_stat_btb_made_pred : _GEN_19132; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19211 = 5'ha == T_29096 ? T_38110_10_stat_btb_mispredicted : _GEN_19133; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19212 = 5'ha == T_29096 ? T_38110_10_stat_bpd_made_pred : _GEN_19134; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19213 = 5'ha == T_29096 ? T_38110_10_stat_bpd_mispredicted : _GEN_19135; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19214 = 5'ha == T_29096 ? T_38110_10_fetch_pc_lob : _GEN_19136; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19215 = 5'ha == T_29096 ? T_38110_10_imm_packed : _GEN_19137; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19216 = 5'ha == T_29096 ? T_38110_10_csr_addr : _GEN_19138; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19217 = 5'ha == T_29096 ? T_38110_10_rob_idx : _GEN_19139; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19218 = 5'ha == T_29096 ? T_38110_10_ldq_idx : _GEN_19140; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19219 = 5'ha == T_29096 ? T_38110_10_stq_idx : _GEN_19141; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19220 = 5'ha == T_29096 ? T_38110_10_brob_idx : _GEN_19142; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19221 = 5'ha == T_29096 ? T_38110_10_pdst : _GEN_19143; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19222 = 5'ha == T_29096 ? T_38110_10_pop1 : _GEN_19144; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19223 = 5'ha == T_29096 ? T_38110_10_pop2 : _GEN_19145; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19224 = 5'ha == T_29096 ? T_38110_10_pop3 : _GEN_19146; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19225 = 5'ha == T_29096 ? T_38110_10_prs1_busy : _GEN_19147; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19226 = 5'ha == T_29096 ? T_38110_10_prs2_busy : _GEN_19148; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19227 = 5'ha == T_29096 ? T_38110_10_prs3_busy : _GEN_19149; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19228 = 5'ha == T_29096 ? T_38110_10_stale_pdst : _GEN_19150; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19229 = 5'ha == T_29096 ? T_38110_10_exception : _GEN_19151; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19230 = 5'ha == T_29096 ? T_38110_10_exc_cause : _GEN_19152; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19231 = 5'ha == T_29096 ? T_38110_10_bypassable : _GEN_19153; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19232 = 5'ha == T_29096 ? T_38110_10_mem_cmd : _GEN_19154; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19233 = 5'ha == T_29096 ? T_38110_10_mem_typ : _GEN_19155; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19234 = 5'ha == T_29096 ? T_38110_10_is_fence : _GEN_19156; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19235 = 5'ha == T_29096 ? T_38110_10_is_fencei : _GEN_19157; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19236 = 5'ha == T_29096 ? T_38110_10_is_store : _GEN_19158; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19237 = 5'ha == T_29096 ? T_38110_10_is_amo : _GEN_19159; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19238 = 5'ha == T_29096 ? T_38110_10_is_load : _GEN_19160; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19239 = 5'ha == T_29096 ? T_38110_10_is_unique : _GEN_19161; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19240 = 5'ha == T_29096 ? T_38110_10_flush_on_commit : _GEN_19162; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19241 = 5'ha == T_29096 ? T_38110_10_ldst : _GEN_19163; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19242 = 5'ha == T_29096 ? T_38110_10_lrs1 : _GEN_19164; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19243 = 5'ha == T_29096 ? T_38110_10_lrs2 : _GEN_19165; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19244 = 5'ha == T_29096 ? T_38110_10_lrs3 : _GEN_19166; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19245 = 5'ha == T_29096 ? T_38110_10_ldst_val : _GEN_19167; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19246 = 5'ha == T_29096 ? T_38110_10_dst_rtype : _GEN_19168; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19247 = 5'ha == T_29096 ? T_38110_10_lrs1_rtype : _GEN_19169; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19248 = 5'ha == T_29096 ? T_38110_10_lrs2_rtype : _GEN_19170; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19249 = 5'ha == T_29096 ? T_38110_10_frs3_en : _GEN_19171; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19250 = 5'ha == T_29096 ? T_38110_10_fp_val : _GEN_19172; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19251 = 5'ha == T_29096 ? T_38110_10_fp_single : _GEN_19173; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19252 = 5'ha == T_29096 ? T_38110_10_xcpt_if : _GEN_19174; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19253 = 5'ha == T_29096 ? T_38110_10_replay_if : _GEN_19175; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19255 = 5'ha == T_29096 ? T_38110_10_debug_events_fetch_seq : _GEN_19177; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19256 = 5'hb == T_29096 ? T_38110_11_valid : _GEN_19178; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19257 = 5'hb == T_29096 ? T_38110_11_iw_state : _GEN_19179; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19258 = 5'hb == T_29096 ? T_38110_11_uopc : _GEN_19180; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19259 = 5'hb == T_29096 ? T_38110_11_inst : _GEN_19181; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19260 = 5'hb == T_29096 ? T_38110_11_pc : _GEN_19182; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19261 = 5'hb == T_29096 ? T_38110_11_fu_code : _GEN_19183; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19262 = 5'hb == T_29096 ? T_38110_11_ctrl_br_type : _GEN_19184; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19263 = 5'hb == T_29096 ? T_38110_11_ctrl_op1_sel : _GEN_19185; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19264 = 5'hb == T_29096 ? T_38110_11_ctrl_op2_sel : _GEN_19186; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19265 = 5'hb == T_29096 ? T_38110_11_ctrl_imm_sel : _GEN_19187; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19266 = 5'hb == T_29096 ? T_38110_11_ctrl_op_fcn : _GEN_19188; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19267 = 5'hb == T_29096 ? T_38110_11_ctrl_fcn_dw : _GEN_19189; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19268 = 5'hb == T_29096 ? T_38110_11_ctrl_rf_wen : _GEN_19190; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19269 = 5'hb == T_29096 ? T_38110_11_ctrl_csr_cmd : _GEN_19191; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19270 = 5'hb == T_29096 ? T_38110_11_ctrl_is_load : _GEN_19192; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19271 = 5'hb == T_29096 ? T_38110_11_ctrl_is_sta : _GEN_19193; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19272 = 5'hb == T_29096 ? T_38110_11_ctrl_is_std : _GEN_19194; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19273 = 5'hb == T_29096 ? T_38110_11_wakeup_delay : _GEN_19195; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19274 = 5'hb == T_29096 ? T_38110_11_allocate_brtag : _GEN_19196; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19275 = 5'hb == T_29096 ? T_38110_11_is_br_or_jmp : _GEN_19197; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19276 = 5'hb == T_29096 ? T_38110_11_is_jump : _GEN_19198; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19277 = 5'hb == T_29096 ? T_38110_11_is_jal : _GEN_19199; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19278 = 5'hb == T_29096 ? T_38110_11_is_ret : _GEN_19200; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19279 = 5'hb == T_29096 ? T_38110_11_is_call : _GEN_19201; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19280 = 5'hb == T_29096 ? T_38110_11_br_mask : _GEN_19202; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19281 = 5'hb == T_29096 ? T_38110_11_br_tag : _GEN_19203; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19282 = 5'hb == T_29096 ? T_38110_11_br_prediction_bpd_predict_val : _GEN_19204; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19283 = 5'hb == T_29096 ? T_38110_11_br_prediction_bpd_predict_taken : _GEN_19205; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19284 = 5'hb == T_29096 ? T_38110_11_br_prediction_btb_hit : _GEN_19206; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19285 = 5'hb == T_29096 ? T_38110_11_br_prediction_btb_predicted : _GEN_19207; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19286 = 5'hb == T_29096 ? T_38110_11_br_prediction_is_br_or_jalr : _GEN_19208; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19287 = 5'hb == T_29096 ? T_38110_11_stat_brjmp_mispredicted : _GEN_19209; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19288 = 5'hb == T_29096 ? T_38110_11_stat_btb_made_pred : _GEN_19210; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19289 = 5'hb == T_29096 ? T_38110_11_stat_btb_mispredicted : _GEN_19211; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19290 = 5'hb == T_29096 ? T_38110_11_stat_bpd_made_pred : _GEN_19212; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19291 = 5'hb == T_29096 ? T_38110_11_stat_bpd_mispredicted : _GEN_19213; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19292 = 5'hb == T_29096 ? T_38110_11_fetch_pc_lob : _GEN_19214; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19293 = 5'hb == T_29096 ? T_38110_11_imm_packed : _GEN_19215; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19294 = 5'hb == T_29096 ? T_38110_11_csr_addr : _GEN_19216; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19295 = 5'hb == T_29096 ? T_38110_11_rob_idx : _GEN_19217; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19296 = 5'hb == T_29096 ? T_38110_11_ldq_idx : _GEN_19218; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19297 = 5'hb == T_29096 ? T_38110_11_stq_idx : _GEN_19219; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19298 = 5'hb == T_29096 ? T_38110_11_brob_idx : _GEN_19220; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19299 = 5'hb == T_29096 ? T_38110_11_pdst : _GEN_19221; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19300 = 5'hb == T_29096 ? T_38110_11_pop1 : _GEN_19222; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19301 = 5'hb == T_29096 ? T_38110_11_pop2 : _GEN_19223; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19302 = 5'hb == T_29096 ? T_38110_11_pop3 : _GEN_19224; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19303 = 5'hb == T_29096 ? T_38110_11_prs1_busy : _GEN_19225; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19304 = 5'hb == T_29096 ? T_38110_11_prs2_busy : _GEN_19226; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19305 = 5'hb == T_29096 ? T_38110_11_prs3_busy : _GEN_19227; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19306 = 5'hb == T_29096 ? T_38110_11_stale_pdst : _GEN_19228; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19307 = 5'hb == T_29096 ? T_38110_11_exception : _GEN_19229; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19308 = 5'hb == T_29096 ? T_38110_11_exc_cause : _GEN_19230; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19309 = 5'hb == T_29096 ? T_38110_11_bypassable : _GEN_19231; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19310 = 5'hb == T_29096 ? T_38110_11_mem_cmd : _GEN_19232; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19311 = 5'hb == T_29096 ? T_38110_11_mem_typ : _GEN_19233; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19312 = 5'hb == T_29096 ? T_38110_11_is_fence : _GEN_19234; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19313 = 5'hb == T_29096 ? T_38110_11_is_fencei : _GEN_19235; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19314 = 5'hb == T_29096 ? T_38110_11_is_store : _GEN_19236; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19315 = 5'hb == T_29096 ? T_38110_11_is_amo : _GEN_19237; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19316 = 5'hb == T_29096 ? T_38110_11_is_load : _GEN_19238; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19317 = 5'hb == T_29096 ? T_38110_11_is_unique : _GEN_19239; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19318 = 5'hb == T_29096 ? T_38110_11_flush_on_commit : _GEN_19240; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19319 = 5'hb == T_29096 ? T_38110_11_ldst : _GEN_19241; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19320 = 5'hb == T_29096 ? T_38110_11_lrs1 : _GEN_19242; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19321 = 5'hb == T_29096 ? T_38110_11_lrs2 : _GEN_19243; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19322 = 5'hb == T_29096 ? T_38110_11_lrs3 : _GEN_19244; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19323 = 5'hb == T_29096 ? T_38110_11_ldst_val : _GEN_19245; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19324 = 5'hb == T_29096 ? T_38110_11_dst_rtype : _GEN_19246; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19325 = 5'hb == T_29096 ? T_38110_11_lrs1_rtype : _GEN_19247; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19326 = 5'hb == T_29096 ? T_38110_11_lrs2_rtype : _GEN_19248; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19327 = 5'hb == T_29096 ? T_38110_11_frs3_en : _GEN_19249; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19328 = 5'hb == T_29096 ? T_38110_11_fp_val : _GEN_19250; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19329 = 5'hb == T_29096 ? T_38110_11_fp_single : _GEN_19251; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19330 = 5'hb == T_29096 ? T_38110_11_xcpt_if : _GEN_19252; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19331 = 5'hb == T_29096 ? T_38110_11_replay_if : _GEN_19253; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19333 = 5'hb == T_29096 ? T_38110_11_debug_events_fetch_seq : _GEN_19255; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19334 = 5'hc == T_29096 ? T_38110_12_valid : _GEN_19256; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19335 = 5'hc == T_29096 ? T_38110_12_iw_state : _GEN_19257; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19336 = 5'hc == T_29096 ? T_38110_12_uopc : _GEN_19258; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19337 = 5'hc == T_29096 ? T_38110_12_inst : _GEN_19259; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19338 = 5'hc == T_29096 ? T_38110_12_pc : _GEN_19260; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19339 = 5'hc == T_29096 ? T_38110_12_fu_code : _GEN_19261; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19340 = 5'hc == T_29096 ? T_38110_12_ctrl_br_type : _GEN_19262; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19341 = 5'hc == T_29096 ? T_38110_12_ctrl_op1_sel : _GEN_19263; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19342 = 5'hc == T_29096 ? T_38110_12_ctrl_op2_sel : _GEN_19264; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19343 = 5'hc == T_29096 ? T_38110_12_ctrl_imm_sel : _GEN_19265; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19344 = 5'hc == T_29096 ? T_38110_12_ctrl_op_fcn : _GEN_19266; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19345 = 5'hc == T_29096 ? T_38110_12_ctrl_fcn_dw : _GEN_19267; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19346 = 5'hc == T_29096 ? T_38110_12_ctrl_rf_wen : _GEN_19268; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19347 = 5'hc == T_29096 ? T_38110_12_ctrl_csr_cmd : _GEN_19269; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19348 = 5'hc == T_29096 ? T_38110_12_ctrl_is_load : _GEN_19270; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19349 = 5'hc == T_29096 ? T_38110_12_ctrl_is_sta : _GEN_19271; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19350 = 5'hc == T_29096 ? T_38110_12_ctrl_is_std : _GEN_19272; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19351 = 5'hc == T_29096 ? T_38110_12_wakeup_delay : _GEN_19273; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19352 = 5'hc == T_29096 ? T_38110_12_allocate_brtag : _GEN_19274; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19353 = 5'hc == T_29096 ? T_38110_12_is_br_or_jmp : _GEN_19275; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19354 = 5'hc == T_29096 ? T_38110_12_is_jump : _GEN_19276; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19355 = 5'hc == T_29096 ? T_38110_12_is_jal : _GEN_19277; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19356 = 5'hc == T_29096 ? T_38110_12_is_ret : _GEN_19278; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19357 = 5'hc == T_29096 ? T_38110_12_is_call : _GEN_19279; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19358 = 5'hc == T_29096 ? T_38110_12_br_mask : _GEN_19280; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19359 = 5'hc == T_29096 ? T_38110_12_br_tag : _GEN_19281; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19360 = 5'hc == T_29096 ? T_38110_12_br_prediction_bpd_predict_val : _GEN_19282; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19361 = 5'hc == T_29096 ? T_38110_12_br_prediction_bpd_predict_taken : _GEN_19283; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19362 = 5'hc == T_29096 ? T_38110_12_br_prediction_btb_hit : _GEN_19284; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19363 = 5'hc == T_29096 ? T_38110_12_br_prediction_btb_predicted : _GEN_19285; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19364 = 5'hc == T_29096 ? T_38110_12_br_prediction_is_br_or_jalr : _GEN_19286; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19365 = 5'hc == T_29096 ? T_38110_12_stat_brjmp_mispredicted : _GEN_19287; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19366 = 5'hc == T_29096 ? T_38110_12_stat_btb_made_pred : _GEN_19288; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19367 = 5'hc == T_29096 ? T_38110_12_stat_btb_mispredicted : _GEN_19289; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19368 = 5'hc == T_29096 ? T_38110_12_stat_bpd_made_pred : _GEN_19290; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19369 = 5'hc == T_29096 ? T_38110_12_stat_bpd_mispredicted : _GEN_19291; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19370 = 5'hc == T_29096 ? T_38110_12_fetch_pc_lob : _GEN_19292; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19371 = 5'hc == T_29096 ? T_38110_12_imm_packed : _GEN_19293; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19372 = 5'hc == T_29096 ? T_38110_12_csr_addr : _GEN_19294; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19373 = 5'hc == T_29096 ? T_38110_12_rob_idx : _GEN_19295; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19374 = 5'hc == T_29096 ? T_38110_12_ldq_idx : _GEN_19296; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19375 = 5'hc == T_29096 ? T_38110_12_stq_idx : _GEN_19297; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19376 = 5'hc == T_29096 ? T_38110_12_brob_idx : _GEN_19298; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19377 = 5'hc == T_29096 ? T_38110_12_pdst : _GEN_19299; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19378 = 5'hc == T_29096 ? T_38110_12_pop1 : _GEN_19300; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19379 = 5'hc == T_29096 ? T_38110_12_pop2 : _GEN_19301; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19380 = 5'hc == T_29096 ? T_38110_12_pop3 : _GEN_19302; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19381 = 5'hc == T_29096 ? T_38110_12_prs1_busy : _GEN_19303; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19382 = 5'hc == T_29096 ? T_38110_12_prs2_busy : _GEN_19304; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19383 = 5'hc == T_29096 ? T_38110_12_prs3_busy : _GEN_19305; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19384 = 5'hc == T_29096 ? T_38110_12_stale_pdst : _GEN_19306; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19385 = 5'hc == T_29096 ? T_38110_12_exception : _GEN_19307; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19386 = 5'hc == T_29096 ? T_38110_12_exc_cause : _GEN_19308; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19387 = 5'hc == T_29096 ? T_38110_12_bypassable : _GEN_19309; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19388 = 5'hc == T_29096 ? T_38110_12_mem_cmd : _GEN_19310; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19389 = 5'hc == T_29096 ? T_38110_12_mem_typ : _GEN_19311; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19390 = 5'hc == T_29096 ? T_38110_12_is_fence : _GEN_19312; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19391 = 5'hc == T_29096 ? T_38110_12_is_fencei : _GEN_19313; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19392 = 5'hc == T_29096 ? T_38110_12_is_store : _GEN_19314; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19393 = 5'hc == T_29096 ? T_38110_12_is_amo : _GEN_19315; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19394 = 5'hc == T_29096 ? T_38110_12_is_load : _GEN_19316; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19395 = 5'hc == T_29096 ? T_38110_12_is_unique : _GEN_19317; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19396 = 5'hc == T_29096 ? T_38110_12_flush_on_commit : _GEN_19318; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19397 = 5'hc == T_29096 ? T_38110_12_ldst : _GEN_19319; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19398 = 5'hc == T_29096 ? T_38110_12_lrs1 : _GEN_19320; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19399 = 5'hc == T_29096 ? T_38110_12_lrs2 : _GEN_19321; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19400 = 5'hc == T_29096 ? T_38110_12_lrs3 : _GEN_19322; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19401 = 5'hc == T_29096 ? T_38110_12_ldst_val : _GEN_19323; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19402 = 5'hc == T_29096 ? T_38110_12_dst_rtype : _GEN_19324; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19403 = 5'hc == T_29096 ? T_38110_12_lrs1_rtype : _GEN_19325; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19404 = 5'hc == T_29096 ? T_38110_12_lrs2_rtype : _GEN_19326; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19405 = 5'hc == T_29096 ? T_38110_12_frs3_en : _GEN_19327; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19406 = 5'hc == T_29096 ? T_38110_12_fp_val : _GEN_19328; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19407 = 5'hc == T_29096 ? T_38110_12_fp_single : _GEN_19329; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19408 = 5'hc == T_29096 ? T_38110_12_xcpt_if : _GEN_19330; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19409 = 5'hc == T_29096 ? T_38110_12_replay_if : _GEN_19331; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19411 = 5'hc == T_29096 ? T_38110_12_debug_events_fetch_seq : _GEN_19333; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19412 = 5'hd == T_29096 ? T_38110_13_valid : _GEN_19334; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19413 = 5'hd == T_29096 ? T_38110_13_iw_state : _GEN_19335; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19414 = 5'hd == T_29096 ? T_38110_13_uopc : _GEN_19336; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19415 = 5'hd == T_29096 ? T_38110_13_inst : _GEN_19337; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19416 = 5'hd == T_29096 ? T_38110_13_pc : _GEN_19338; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19417 = 5'hd == T_29096 ? T_38110_13_fu_code : _GEN_19339; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19418 = 5'hd == T_29096 ? T_38110_13_ctrl_br_type : _GEN_19340; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19419 = 5'hd == T_29096 ? T_38110_13_ctrl_op1_sel : _GEN_19341; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19420 = 5'hd == T_29096 ? T_38110_13_ctrl_op2_sel : _GEN_19342; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19421 = 5'hd == T_29096 ? T_38110_13_ctrl_imm_sel : _GEN_19343; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19422 = 5'hd == T_29096 ? T_38110_13_ctrl_op_fcn : _GEN_19344; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19423 = 5'hd == T_29096 ? T_38110_13_ctrl_fcn_dw : _GEN_19345; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19424 = 5'hd == T_29096 ? T_38110_13_ctrl_rf_wen : _GEN_19346; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19425 = 5'hd == T_29096 ? T_38110_13_ctrl_csr_cmd : _GEN_19347; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19426 = 5'hd == T_29096 ? T_38110_13_ctrl_is_load : _GEN_19348; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19427 = 5'hd == T_29096 ? T_38110_13_ctrl_is_sta : _GEN_19349; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19428 = 5'hd == T_29096 ? T_38110_13_ctrl_is_std : _GEN_19350; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19429 = 5'hd == T_29096 ? T_38110_13_wakeup_delay : _GEN_19351; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19430 = 5'hd == T_29096 ? T_38110_13_allocate_brtag : _GEN_19352; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19431 = 5'hd == T_29096 ? T_38110_13_is_br_or_jmp : _GEN_19353; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19432 = 5'hd == T_29096 ? T_38110_13_is_jump : _GEN_19354; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19433 = 5'hd == T_29096 ? T_38110_13_is_jal : _GEN_19355; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19434 = 5'hd == T_29096 ? T_38110_13_is_ret : _GEN_19356; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19435 = 5'hd == T_29096 ? T_38110_13_is_call : _GEN_19357; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19436 = 5'hd == T_29096 ? T_38110_13_br_mask : _GEN_19358; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19437 = 5'hd == T_29096 ? T_38110_13_br_tag : _GEN_19359; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19438 = 5'hd == T_29096 ? T_38110_13_br_prediction_bpd_predict_val : _GEN_19360; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19439 = 5'hd == T_29096 ? T_38110_13_br_prediction_bpd_predict_taken : _GEN_19361; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19440 = 5'hd == T_29096 ? T_38110_13_br_prediction_btb_hit : _GEN_19362; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19441 = 5'hd == T_29096 ? T_38110_13_br_prediction_btb_predicted : _GEN_19363; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19442 = 5'hd == T_29096 ? T_38110_13_br_prediction_is_br_or_jalr : _GEN_19364; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19443 = 5'hd == T_29096 ? T_38110_13_stat_brjmp_mispredicted : _GEN_19365; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19444 = 5'hd == T_29096 ? T_38110_13_stat_btb_made_pred : _GEN_19366; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19445 = 5'hd == T_29096 ? T_38110_13_stat_btb_mispredicted : _GEN_19367; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19446 = 5'hd == T_29096 ? T_38110_13_stat_bpd_made_pred : _GEN_19368; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19447 = 5'hd == T_29096 ? T_38110_13_stat_bpd_mispredicted : _GEN_19369; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19448 = 5'hd == T_29096 ? T_38110_13_fetch_pc_lob : _GEN_19370; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19449 = 5'hd == T_29096 ? T_38110_13_imm_packed : _GEN_19371; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19450 = 5'hd == T_29096 ? T_38110_13_csr_addr : _GEN_19372; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19451 = 5'hd == T_29096 ? T_38110_13_rob_idx : _GEN_19373; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19452 = 5'hd == T_29096 ? T_38110_13_ldq_idx : _GEN_19374; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19453 = 5'hd == T_29096 ? T_38110_13_stq_idx : _GEN_19375; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19454 = 5'hd == T_29096 ? T_38110_13_brob_idx : _GEN_19376; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19455 = 5'hd == T_29096 ? T_38110_13_pdst : _GEN_19377; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19456 = 5'hd == T_29096 ? T_38110_13_pop1 : _GEN_19378; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19457 = 5'hd == T_29096 ? T_38110_13_pop2 : _GEN_19379; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19458 = 5'hd == T_29096 ? T_38110_13_pop3 : _GEN_19380; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19459 = 5'hd == T_29096 ? T_38110_13_prs1_busy : _GEN_19381; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19460 = 5'hd == T_29096 ? T_38110_13_prs2_busy : _GEN_19382; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19461 = 5'hd == T_29096 ? T_38110_13_prs3_busy : _GEN_19383; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19462 = 5'hd == T_29096 ? T_38110_13_stale_pdst : _GEN_19384; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19463 = 5'hd == T_29096 ? T_38110_13_exception : _GEN_19385; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19464 = 5'hd == T_29096 ? T_38110_13_exc_cause : _GEN_19386; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19465 = 5'hd == T_29096 ? T_38110_13_bypassable : _GEN_19387; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19466 = 5'hd == T_29096 ? T_38110_13_mem_cmd : _GEN_19388; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19467 = 5'hd == T_29096 ? T_38110_13_mem_typ : _GEN_19389; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19468 = 5'hd == T_29096 ? T_38110_13_is_fence : _GEN_19390; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19469 = 5'hd == T_29096 ? T_38110_13_is_fencei : _GEN_19391; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19470 = 5'hd == T_29096 ? T_38110_13_is_store : _GEN_19392; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19471 = 5'hd == T_29096 ? T_38110_13_is_amo : _GEN_19393; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19472 = 5'hd == T_29096 ? T_38110_13_is_load : _GEN_19394; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19473 = 5'hd == T_29096 ? T_38110_13_is_unique : _GEN_19395; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19474 = 5'hd == T_29096 ? T_38110_13_flush_on_commit : _GEN_19396; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19475 = 5'hd == T_29096 ? T_38110_13_ldst : _GEN_19397; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19476 = 5'hd == T_29096 ? T_38110_13_lrs1 : _GEN_19398; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19477 = 5'hd == T_29096 ? T_38110_13_lrs2 : _GEN_19399; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19478 = 5'hd == T_29096 ? T_38110_13_lrs3 : _GEN_19400; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19479 = 5'hd == T_29096 ? T_38110_13_ldst_val : _GEN_19401; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19480 = 5'hd == T_29096 ? T_38110_13_dst_rtype : _GEN_19402; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19481 = 5'hd == T_29096 ? T_38110_13_lrs1_rtype : _GEN_19403; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19482 = 5'hd == T_29096 ? T_38110_13_lrs2_rtype : _GEN_19404; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19483 = 5'hd == T_29096 ? T_38110_13_frs3_en : _GEN_19405; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19484 = 5'hd == T_29096 ? T_38110_13_fp_val : _GEN_19406; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19485 = 5'hd == T_29096 ? T_38110_13_fp_single : _GEN_19407; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19486 = 5'hd == T_29096 ? T_38110_13_xcpt_if : _GEN_19408; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19487 = 5'hd == T_29096 ? T_38110_13_replay_if : _GEN_19409; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19489 = 5'hd == T_29096 ? T_38110_13_debug_events_fetch_seq : _GEN_19411; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19490 = 5'he == T_29096 ? T_38110_14_valid : _GEN_19412; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19491 = 5'he == T_29096 ? T_38110_14_iw_state : _GEN_19413; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19492 = 5'he == T_29096 ? T_38110_14_uopc : _GEN_19414; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19493 = 5'he == T_29096 ? T_38110_14_inst : _GEN_19415; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19494 = 5'he == T_29096 ? T_38110_14_pc : _GEN_19416; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19495 = 5'he == T_29096 ? T_38110_14_fu_code : _GEN_19417; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19496 = 5'he == T_29096 ? T_38110_14_ctrl_br_type : _GEN_19418; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19497 = 5'he == T_29096 ? T_38110_14_ctrl_op1_sel : _GEN_19419; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19498 = 5'he == T_29096 ? T_38110_14_ctrl_op2_sel : _GEN_19420; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19499 = 5'he == T_29096 ? T_38110_14_ctrl_imm_sel : _GEN_19421; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19500 = 5'he == T_29096 ? T_38110_14_ctrl_op_fcn : _GEN_19422; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19501 = 5'he == T_29096 ? T_38110_14_ctrl_fcn_dw : _GEN_19423; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19502 = 5'he == T_29096 ? T_38110_14_ctrl_rf_wen : _GEN_19424; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19503 = 5'he == T_29096 ? T_38110_14_ctrl_csr_cmd : _GEN_19425; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19504 = 5'he == T_29096 ? T_38110_14_ctrl_is_load : _GEN_19426; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19505 = 5'he == T_29096 ? T_38110_14_ctrl_is_sta : _GEN_19427; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19506 = 5'he == T_29096 ? T_38110_14_ctrl_is_std : _GEN_19428; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19507 = 5'he == T_29096 ? T_38110_14_wakeup_delay : _GEN_19429; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19508 = 5'he == T_29096 ? T_38110_14_allocate_brtag : _GEN_19430; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19509 = 5'he == T_29096 ? T_38110_14_is_br_or_jmp : _GEN_19431; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19510 = 5'he == T_29096 ? T_38110_14_is_jump : _GEN_19432; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19511 = 5'he == T_29096 ? T_38110_14_is_jal : _GEN_19433; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19512 = 5'he == T_29096 ? T_38110_14_is_ret : _GEN_19434; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19513 = 5'he == T_29096 ? T_38110_14_is_call : _GEN_19435; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19514 = 5'he == T_29096 ? T_38110_14_br_mask : _GEN_19436; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19515 = 5'he == T_29096 ? T_38110_14_br_tag : _GEN_19437; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19516 = 5'he == T_29096 ? T_38110_14_br_prediction_bpd_predict_val : _GEN_19438; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19517 = 5'he == T_29096 ? T_38110_14_br_prediction_bpd_predict_taken : _GEN_19439; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19518 = 5'he == T_29096 ? T_38110_14_br_prediction_btb_hit : _GEN_19440; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19519 = 5'he == T_29096 ? T_38110_14_br_prediction_btb_predicted : _GEN_19441; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19520 = 5'he == T_29096 ? T_38110_14_br_prediction_is_br_or_jalr : _GEN_19442; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19521 = 5'he == T_29096 ? T_38110_14_stat_brjmp_mispredicted : _GEN_19443; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19522 = 5'he == T_29096 ? T_38110_14_stat_btb_made_pred : _GEN_19444; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19523 = 5'he == T_29096 ? T_38110_14_stat_btb_mispredicted : _GEN_19445; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19524 = 5'he == T_29096 ? T_38110_14_stat_bpd_made_pred : _GEN_19446; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19525 = 5'he == T_29096 ? T_38110_14_stat_bpd_mispredicted : _GEN_19447; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19526 = 5'he == T_29096 ? T_38110_14_fetch_pc_lob : _GEN_19448; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19527 = 5'he == T_29096 ? T_38110_14_imm_packed : _GEN_19449; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19528 = 5'he == T_29096 ? T_38110_14_csr_addr : _GEN_19450; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19529 = 5'he == T_29096 ? T_38110_14_rob_idx : _GEN_19451; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19530 = 5'he == T_29096 ? T_38110_14_ldq_idx : _GEN_19452; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19531 = 5'he == T_29096 ? T_38110_14_stq_idx : _GEN_19453; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19532 = 5'he == T_29096 ? T_38110_14_brob_idx : _GEN_19454; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19533 = 5'he == T_29096 ? T_38110_14_pdst : _GEN_19455; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19534 = 5'he == T_29096 ? T_38110_14_pop1 : _GEN_19456; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19535 = 5'he == T_29096 ? T_38110_14_pop2 : _GEN_19457; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19536 = 5'he == T_29096 ? T_38110_14_pop3 : _GEN_19458; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19537 = 5'he == T_29096 ? T_38110_14_prs1_busy : _GEN_19459; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19538 = 5'he == T_29096 ? T_38110_14_prs2_busy : _GEN_19460; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19539 = 5'he == T_29096 ? T_38110_14_prs3_busy : _GEN_19461; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19540 = 5'he == T_29096 ? T_38110_14_stale_pdst : _GEN_19462; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19541 = 5'he == T_29096 ? T_38110_14_exception : _GEN_19463; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19542 = 5'he == T_29096 ? T_38110_14_exc_cause : _GEN_19464; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19543 = 5'he == T_29096 ? T_38110_14_bypassable : _GEN_19465; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19544 = 5'he == T_29096 ? T_38110_14_mem_cmd : _GEN_19466; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19545 = 5'he == T_29096 ? T_38110_14_mem_typ : _GEN_19467; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19546 = 5'he == T_29096 ? T_38110_14_is_fence : _GEN_19468; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19547 = 5'he == T_29096 ? T_38110_14_is_fencei : _GEN_19469; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19548 = 5'he == T_29096 ? T_38110_14_is_store : _GEN_19470; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19549 = 5'he == T_29096 ? T_38110_14_is_amo : _GEN_19471; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19550 = 5'he == T_29096 ? T_38110_14_is_load : _GEN_19472; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19551 = 5'he == T_29096 ? T_38110_14_is_unique : _GEN_19473; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19552 = 5'he == T_29096 ? T_38110_14_flush_on_commit : _GEN_19474; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19553 = 5'he == T_29096 ? T_38110_14_ldst : _GEN_19475; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19554 = 5'he == T_29096 ? T_38110_14_lrs1 : _GEN_19476; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19555 = 5'he == T_29096 ? T_38110_14_lrs2 : _GEN_19477; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19556 = 5'he == T_29096 ? T_38110_14_lrs3 : _GEN_19478; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19557 = 5'he == T_29096 ? T_38110_14_ldst_val : _GEN_19479; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19558 = 5'he == T_29096 ? T_38110_14_dst_rtype : _GEN_19480; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19559 = 5'he == T_29096 ? T_38110_14_lrs1_rtype : _GEN_19481; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19560 = 5'he == T_29096 ? T_38110_14_lrs2_rtype : _GEN_19482; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19561 = 5'he == T_29096 ? T_38110_14_frs3_en : _GEN_19483; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19562 = 5'he == T_29096 ? T_38110_14_fp_val : _GEN_19484; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19563 = 5'he == T_29096 ? T_38110_14_fp_single : _GEN_19485; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19564 = 5'he == T_29096 ? T_38110_14_xcpt_if : _GEN_19486; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19565 = 5'he == T_29096 ? T_38110_14_replay_if : _GEN_19487; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19567 = 5'he == T_29096 ? T_38110_14_debug_events_fetch_seq : _GEN_19489; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19568 = 5'hf == T_29096 ? T_38110_15_valid : _GEN_19490; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19569 = 5'hf == T_29096 ? T_38110_15_iw_state : _GEN_19491; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19570 = 5'hf == T_29096 ? T_38110_15_uopc : _GEN_19492; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19571 = 5'hf == T_29096 ? T_38110_15_inst : _GEN_19493; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19572 = 5'hf == T_29096 ? T_38110_15_pc : _GEN_19494; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19573 = 5'hf == T_29096 ? T_38110_15_fu_code : _GEN_19495; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19574 = 5'hf == T_29096 ? T_38110_15_ctrl_br_type : _GEN_19496; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19575 = 5'hf == T_29096 ? T_38110_15_ctrl_op1_sel : _GEN_19497; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19576 = 5'hf == T_29096 ? T_38110_15_ctrl_op2_sel : _GEN_19498; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19577 = 5'hf == T_29096 ? T_38110_15_ctrl_imm_sel : _GEN_19499; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19578 = 5'hf == T_29096 ? T_38110_15_ctrl_op_fcn : _GEN_19500; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19579 = 5'hf == T_29096 ? T_38110_15_ctrl_fcn_dw : _GEN_19501; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19580 = 5'hf == T_29096 ? T_38110_15_ctrl_rf_wen : _GEN_19502; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19581 = 5'hf == T_29096 ? T_38110_15_ctrl_csr_cmd : _GEN_19503; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19582 = 5'hf == T_29096 ? T_38110_15_ctrl_is_load : _GEN_19504; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19583 = 5'hf == T_29096 ? T_38110_15_ctrl_is_sta : _GEN_19505; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19584 = 5'hf == T_29096 ? T_38110_15_ctrl_is_std : _GEN_19506; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19585 = 5'hf == T_29096 ? T_38110_15_wakeup_delay : _GEN_19507; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19586 = 5'hf == T_29096 ? T_38110_15_allocate_brtag : _GEN_19508; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19587 = 5'hf == T_29096 ? T_38110_15_is_br_or_jmp : _GEN_19509; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19588 = 5'hf == T_29096 ? T_38110_15_is_jump : _GEN_19510; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19589 = 5'hf == T_29096 ? T_38110_15_is_jal : _GEN_19511; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19590 = 5'hf == T_29096 ? T_38110_15_is_ret : _GEN_19512; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19591 = 5'hf == T_29096 ? T_38110_15_is_call : _GEN_19513; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19592 = 5'hf == T_29096 ? T_38110_15_br_mask : _GEN_19514; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19593 = 5'hf == T_29096 ? T_38110_15_br_tag : _GEN_19515; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19594 = 5'hf == T_29096 ? T_38110_15_br_prediction_bpd_predict_val : _GEN_19516; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19595 = 5'hf == T_29096 ? T_38110_15_br_prediction_bpd_predict_taken : _GEN_19517; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19596 = 5'hf == T_29096 ? T_38110_15_br_prediction_btb_hit : _GEN_19518; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19597 = 5'hf == T_29096 ? T_38110_15_br_prediction_btb_predicted : _GEN_19519; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19598 = 5'hf == T_29096 ? T_38110_15_br_prediction_is_br_or_jalr : _GEN_19520; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19599 = 5'hf == T_29096 ? T_38110_15_stat_brjmp_mispredicted : _GEN_19521; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19600 = 5'hf == T_29096 ? T_38110_15_stat_btb_made_pred : _GEN_19522; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19601 = 5'hf == T_29096 ? T_38110_15_stat_btb_mispredicted : _GEN_19523; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19602 = 5'hf == T_29096 ? T_38110_15_stat_bpd_made_pred : _GEN_19524; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19603 = 5'hf == T_29096 ? T_38110_15_stat_bpd_mispredicted : _GEN_19525; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19604 = 5'hf == T_29096 ? T_38110_15_fetch_pc_lob : _GEN_19526; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19605 = 5'hf == T_29096 ? T_38110_15_imm_packed : _GEN_19527; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19606 = 5'hf == T_29096 ? T_38110_15_csr_addr : _GEN_19528; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19607 = 5'hf == T_29096 ? T_38110_15_rob_idx : _GEN_19529; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19608 = 5'hf == T_29096 ? T_38110_15_ldq_idx : _GEN_19530; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19609 = 5'hf == T_29096 ? T_38110_15_stq_idx : _GEN_19531; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19610 = 5'hf == T_29096 ? T_38110_15_brob_idx : _GEN_19532; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19611 = 5'hf == T_29096 ? T_38110_15_pdst : _GEN_19533; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19612 = 5'hf == T_29096 ? T_38110_15_pop1 : _GEN_19534; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19613 = 5'hf == T_29096 ? T_38110_15_pop2 : _GEN_19535; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19614 = 5'hf == T_29096 ? T_38110_15_pop3 : _GEN_19536; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19615 = 5'hf == T_29096 ? T_38110_15_prs1_busy : _GEN_19537; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19616 = 5'hf == T_29096 ? T_38110_15_prs2_busy : _GEN_19538; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19617 = 5'hf == T_29096 ? T_38110_15_prs3_busy : _GEN_19539; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19618 = 5'hf == T_29096 ? T_38110_15_stale_pdst : _GEN_19540; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19619 = 5'hf == T_29096 ? T_38110_15_exception : _GEN_19541; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19620 = 5'hf == T_29096 ? T_38110_15_exc_cause : _GEN_19542; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19621 = 5'hf == T_29096 ? T_38110_15_bypassable : _GEN_19543; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19622 = 5'hf == T_29096 ? T_38110_15_mem_cmd : _GEN_19544; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19623 = 5'hf == T_29096 ? T_38110_15_mem_typ : _GEN_19545; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19624 = 5'hf == T_29096 ? T_38110_15_is_fence : _GEN_19546; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19625 = 5'hf == T_29096 ? T_38110_15_is_fencei : _GEN_19547; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19626 = 5'hf == T_29096 ? T_38110_15_is_store : _GEN_19548; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19627 = 5'hf == T_29096 ? T_38110_15_is_amo : _GEN_19549; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19628 = 5'hf == T_29096 ? T_38110_15_is_load : _GEN_19550; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19629 = 5'hf == T_29096 ? T_38110_15_is_unique : _GEN_19551; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19630 = 5'hf == T_29096 ? T_38110_15_flush_on_commit : _GEN_19552; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19631 = 5'hf == T_29096 ? T_38110_15_ldst : _GEN_19553; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19632 = 5'hf == T_29096 ? T_38110_15_lrs1 : _GEN_19554; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19633 = 5'hf == T_29096 ? T_38110_15_lrs2 : _GEN_19555; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19634 = 5'hf == T_29096 ? T_38110_15_lrs3 : _GEN_19556; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19635 = 5'hf == T_29096 ? T_38110_15_ldst_val : _GEN_19557; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19636 = 5'hf == T_29096 ? T_38110_15_dst_rtype : _GEN_19558; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19637 = 5'hf == T_29096 ? T_38110_15_lrs1_rtype : _GEN_19559; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19638 = 5'hf == T_29096 ? T_38110_15_lrs2_rtype : _GEN_19560; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19639 = 5'hf == T_29096 ? T_38110_15_frs3_en : _GEN_19561; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19640 = 5'hf == T_29096 ? T_38110_15_fp_val : _GEN_19562; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19641 = 5'hf == T_29096 ? T_38110_15_fp_single : _GEN_19563; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19642 = 5'hf == T_29096 ? T_38110_15_xcpt_if : _GEN_19564; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19643 = 5'hf == T_29096 ? T_38110_15_replay_if : _GEN_19565; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19645 = 5'hf == T_29096 ? T_38110_15_debug_events_fetch_seq : _GEN_19567; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19646 = 5'h10 == T_29096 ? T_38110_16_valid : _GEN_19568; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19647 = 5'h10 == T_29096 ? T_38110_16_iw_state : _GEN_19569; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19648 = 5'h10 == T_29096 ? T_38110_16_uopc : _GEN_19570; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19649 = 5'h10 == T_29096 ? T_38110_16_inst : _GEN_19571; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19650 = 5'h10 == T_29096 ? T_38110_16_pc : _GEN_19572; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19651 = 5'h10 == T_29096 ? T_38110_16_fu_code : _GEN_19573; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19652 = 5'h10 == T_29096 ? T_38110_16_ctrl_br_type : _GEN_19574; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19653 = 5'h10 == T_29096 ? T_38110_16_ctrl_op1_sel : _GEN_19575; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19654 = 5'h10 == T_29096 ? T_38110_16_ctrl_op2_sel : _GEN_19576; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19655 = 5'h10 == T_29096 ? T_38110_16_ctrl_imm_sel : _GEN_19577; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19656 = 5'h10 == T_29096 ? T_38110_16_ctrl_op_fcn : _GEN_19578; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19657 = 5'h10 == T_29096 ? T_38110_16_ctrl_fcn_dw : _GEN_19579; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19658 = 5'h10 == T_29096 ? T_38110_16_ctrl_rf_wen : _GEN_19580; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19659 = 5'h10 == T_29096 ? T_38110_16_ctrl_csr_cmd : _GEN_19581; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19660 = 5'h10 == T_29096 ? T_38110_16_ctrl_is_load : _GEN_19582; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19661 = 5'h10 == T_29096 ? T_38110_16_ctrl_is_sta : _GEN_19583; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19662 = 5'h10 == T_29096 ? T_38110_16_ctrl_is_std : _GEN_19584; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19663 = 5'h10 == T_29096 ? T_38110_16_wakeup_delay : _GEN_19585; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19664 = 5'h10 == T_29096 ? T_38110_16_allocate_brtag : _GEN_19586; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19665 = 5'h10 == T_29096 ? T_38110_16_is_br_or_jmp : _GEN_19587; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19666 = 5'h10 == T_29096 ? T_38110_16_is_jump : _GEN_19588; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19667 = 5'h10 == T_29096 ? T_38110_16_is_jal : _GEN_19589; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19668 = 5'h10 == T_29096 ? T_38110_16_is_ret : _GEN_19590; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19669 = 5'h10 == T_29096 ? T_38110_16_is_call : _GEN_19591; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19670 = 5'h10 == T_29096 ? T_38110_16_br_mask : _GEN_19592; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19671 = 5'h10 == T_29096 ? T_38110_16_br_tag : _GEN_19593; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19672 = 5'h10 == T_29096 ? T_38110_16_br_prediction_bpd_predict_val : _GEN_19594; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19673 = 5'h10 == T_29096 ? T_38110_16_br_prediction_bpd_predict_taken : _GEN_19595; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19674 = 5'h10 == T_29096 ? T_38110_16_br_prediction_btb_hit : _GEN_19596; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19675 = 5'h10 == T_29096 ? T_38110_16_br_prediction_btb_predicted : _GEN_19597; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19676 = 5'h10 == T_29096 ? T_38110_16_br_prediction_is_br_or_jalr : _GEN_19598; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19677 = 5'h10 == T_29096 ? T_38110_16_stat_brjmp_mispredicted : _GEN_19599; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19678 = 5'h10 == T_29096 ? T_38110_16_stat_btb_made_pred : _GEN_19600; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19679 = 5'h10 == T_29096 ? T_38110_16_stat_btb_mispredicted : _GEN_19601; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19680 = 5'h10 == T_29096 ? T_38110_16_stat_bpd_made_pred : _GEN_19602; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19681 = 5'h10 == T_29096 ? T_38110_16_stat_bpd_mispredicted : _GEN_19603; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19682 = 5'h10 == T_29096 ? T_38110_16_fetch_pc_lob : _GEN_19604; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19683 = 5'h10 == T_29096 ? T_38110_16_imm_packed : _GEN_19605; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19684 = 5'h10 == T_29096 ? T_38110_16_csr_addr : _GEN_19606; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19685 = 5'h10 == T_29096 ? T_38110_16_rob_idx : _GEN_19607; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19686 = 5'h10 == T_29096 ? T_38110_16_ldq_idx : _GEN_19608; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19687 = 5'h10 == T_29096 ? T_38110_16_stq_idx : _GEN_19609; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19688 = 5'h10 == T_29096 ? T_38110_16_brob_idx : _GEN_19610; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19689 = 5'h10 == T_29096 ? T_38110_16_pdst : _GEN_19611; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19690 = 5'h10 == T_29096 ? T_38110_16_pop1 : _GEN_19612; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19691 = 5'h10 == T_29096 ? T_38110_16_pop2 : _GEN_19613; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19692 = 5'h10 == T_29096 ? T_38110_16_pop3 : _GEN_19614; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19693 = 5'h10 == T_29096 ? T_38110_16_prs1_busy : _GEN_19615; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19694 = 5'h10 == T_29096 ? T_38110_16_prs2_busy : _GEN_19616; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19695 = 5'h10 == T_29096 ? T_38110_16_prs3_busy : _GEN_19617; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19696 = 5'h10 == T_29096 ? T_38110_16_stale_pdst : _GEN_19618; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19697 = 5'h10 == T_29096 ? T_38110_16_exception : _GEN_19619; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19698 = 5'h10 == T_29096 ? T_38110_16_exc_cause : _GEN_19620; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19699 = 5'h10 == T_29096 ? T_38110_16_bypassable : _GEN_19621; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19700 = 5'h10 == T_29096 ? T_38110_16_mem_cmd : _GEN_19622; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19701 = 5'h10 == T_29096 ? T_38110_16_mem_typ : _GEN_19623; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19702 = 5'h10 == T_29096 ? T_38110_16_is_fence : _GEN_19624; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19703 = 5'h10 == T_29096 ? T_38110_16_is_fencei : _GEN_19625; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19704 = 5'h10 == T_29096 ? T_38110_16_is_store : _GEN_19626; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19705 = 5'h10 == T_29096 ? T_38110_16_is_amo : _GEN_19627; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19706 = 5'h10 == T_29096 ? T_38110_16_is_load : _GEN_19628; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19707 = 5'h10 == T_29096 ? T_38110_16_is_unique : _GEN_19629; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19708 = 5'h10 == T_29096 ? T_38110_16_flush_on_commit : _GEN_19630; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19709 = 5'h10 == T_29096 ? T_38110_16_ldst : _GEN_19631; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19710 = 5'h10 == T_29096 ? T_38110_16_lrs1 : _GEN_19632; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19711 = 5'h10 == T_29096 ? T_38110_16_lrs2 : _GEN_19633; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19712 = 5'h10 == T_29096 ? T_38110_16_lrs3 : _GEN_19634; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19713 = 5'h10 == T_29096 ? T_38110_16_ldst_val : _GEN_19635; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19714 = 5'h10 == T_29096 ? T_38110_16_dst_rtype : _GEN_19636; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19715 = 5'h10 == T_29096 ? T_38110_16_lrs1_rtype : _GEN_19637; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19716 = 5'h10 == T_29096 ? T_38110_16_lrs2_rtype : _GEN_19638; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19717 = 5'h10 == T_29096 ? T_38110_16_frs3_en : _GEN_19639; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19718 = 5'h10 == T_29096 ? T_38110_16_fp_val : _GEN_19640; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19719 = 5'h10 == T_29096 ? T_38110_16_fp_single : _GEN_19641; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19720 = 5'h10 == T_29096 ? T_38110_16_xcpt_if : _GEN_19642; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19721 = 5'h10 == T_29096 ? T_38110_16_replay_if : _GEN_19643; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19723 = 5'h10 == T_29096 ? T_38110_16_debug_events_fetch_seq : _GEN_19645; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19724 = 5'h11 == T_29096 ? T_38110_17_valid : _GEN_19646; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19725 = 5'h11 == T_29096 ? T_38110_17_iw_state : _GEN_19647; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19726 = 5'h11 == T_29096 ? T_38110_17_uopc : _GEN_19648; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19727 = 5'h11 == T_29096 ? T_38110_17_inst : _GEN_19649; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19728 = 5'h11 == T_29096 ? T_38110_17_pc : _GEN_19650; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19729 = 5'h11 == T_29096 ? T_38110_17_fu_code : _GEN_19651; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19730 = 5'h11 == T_29096 ? T_38110_17_ctrl_br_type : _GEN_19652; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19731 = 5'h11 == T_29096 ? T_38110_17_ctrl_op1_sel : _GEN_19653; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19732 = 5'h11 == T_29096 ? T_38110_17_ctrl_op2_sel : _GEN_19654; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19733 = 5'h11 == T_29096 ? T_38110_17_ctrl_imm_sel : _GEN_19655; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19734 = 5'h11 == T_29096 ? T_38110_17_ctrl_op_fcn : _GEN_19656; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19735 = 5'h11 == T_29096 ? T_38110_17_ctrl_fcn_dw : _GEN_19657; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19736 = 5'h11 == T_29096 ? T_38110_17_ctrl_rf_wen : _GEN_19658; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19737 = 5'h11 == T_29096 ? T_38110_17_ctrl_csr_cmd : _GEN_19659; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19738 = 5'h11 == T_29096 ? T_38110_17_ctrl_is_load : _GEN_19660; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19739 = 5'h11 == T_29096 ? T_38110_17_ctrl_is_sta : _GEN_19661; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19740 = 5'h11 == T_29096 ? T_38110_17_ctrl_is_std : _GEN_19662; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19741 = 5'h11 == T_29096 ? T_38110_17_wakeup_delay : _GEN_19663; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19742 = 5'h11 == T_29096 ? T_38110_17_allocate_brtag : _GEN_19664; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19743 = 5'h11 == T_29096 ? T_38110_17_is_br_or_jmp : _GEN_19665; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19744 = 5'h11 == T_29096 ? T_38110_17_is_jump : _GEN_19666; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19745 = 5'h11 == T_29096 ? T_38110_17_is_jal : _GEN_19667; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19746 = 5'h11 == T_29096 ? T_38110_17_is_ret : _GEN_19668; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19747 = 5'h11 == T_29096 ? T_38110_17_is_call : _GEN_19669; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19748 = 5'h11 == T_29096 ? T_38110_17_br_mask : _GEN_19670; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19749 = 5'h11 == T_29096 ? T_38110_17_br_tag : _GEN_19671; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19750 = 5'h11 == T_29096 ? T_38110_17_br_prediction_bpd_predict_val : _GEN_19672; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19751 = 5'h11 == T_29096 ? T_38110_17_br_prediction_bpd_predict_taken : _GEN_19673; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19752 = 5'h11 == T_29096 ? T_38110_17_br_prediction_btb_hit : _GEN_19674; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19753 = 5'h11 == T_29096 ? T_38110_17_br_prediction_btb_predicted : _GEN_19675; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19754 = 5'h11 == T_29096 ? T_38110_17_br_prediction_is_br_or_jalr : _GEN_19676; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19755 = 5'h11 == T_29096 ? T_38110_17_stat_brjmp_mispredicted : _GEN_19677; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19756 = 5'h11 == T_29096 ? T_38110_17_stat_btb_made_pred : _GEN_19678; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19757 = 5'h11 == T_29096 ? T_38110_17_stat_btb_mispredicted : _GEN_19679; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19758 = 5'h11 == T_29096 ? T_38110_17_stat_bpd_made_pred : _GEN_19680; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19759 = 5'h11 == T_29096 ? T_38110_17_stat_bpd_mispredicted : _GEN_19681; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19760 = 5'h11 == T_29096 ? T_38110_17_fetch_pc_lob : _GEN_19682; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19761 = 5'h11 == T_29096 ? T_38110_17_imm_packed : _GEN_19683; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19762 = 5'h11 == T_29096 ? T_38110_17_csr_addr : _GEN_19684; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19763 = 5'h11 == T_29096 ? T_38110_17_rob_idx : _GEN_19685; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19764 = 5'h11 == T_29096 ? T_38110_17_ldq_idx : _GEN_19686; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19765 = 5'h11 == T_29096 ? T_38110_17_stq_idx : _GEN_19687; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19766 = 5'h11 == T_29096 ? T_38110_17_brob_idx : _GEN_19688; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19767 = 5'h11 == T_29096 ? T_38110_17_pdst : _GEN_19689; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19768 = 5'h11 == T_29096 ? T_38110_17_pop1 : _GEN_19690; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19769 = 5'h11 == T_29096 ? T_38110_17_pop2 : _GEN_19691; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19770 = 5'h11 == T_29096 ? T_38110_17_pop3 : _GEN_19692; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19771 = 5'h11 == T_29096 ? T_38110_17_prs1_busy : _GEN_19693; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19772 = 5'h11 == T_29096 ? T_38110_17_prs2_busy : _GEN_19694; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19773 = 5'h11 == T_29096 ? T_38110_17_prs3_busy : _GEN_19695; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19774 = 5'h11 == T_29096 ? T_38110_17_stale_pdst : _GEN_19696; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19775 = 5'h11 == T_29096 ? T_38110_17_exception : _GEN_19697; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19776 = 5'h11 == T_29096 ? T_38110_17_exc_cause : _GEN_19698; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19777 = 5'h11 == T_29096 ? T_38110_17_bypassable : _GEN_19699; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19778 = 5'h11 == T_29096 ? T_38110_17_mem_cmd : _GEN_19700; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19779 = 5'h11 == T_29096 ? T_38110_17_mem_typ : _GEN_19701; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19780 = 5'h11 == T_29096 ? T_38110_17_is_fence : _GEN_19702; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19781 = 5'h11 == T_29096 ? T_38110_17_is_fencei : _GEN_19703; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19782 = 5'h11 == T_29096 ? T_38110_17_is_store : _GEN_19704; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19783 = 5'h11 == T_29096 ? T_38110_17_is_amo : _GEN_19705; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19784 = 5'h11 == T_29096 ? T_38110_17_is_load : _GEN_19706; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19785 = 5'h11 == T_29096 ? T_38110_17_is_unique : _GEN_19707; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19786 = 5'h11 == T_29096 ? T_38110_17_flush_on_commit : _GEN_19708; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19787 = 5'h11 == T_29096 ? T_38110_17_ldst : _GEN_19709; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19788 = 5'h11 == T_29096 ? T_38110_17_lrs1 : _GEN_19710; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19789 = 5'h11 == T_29096 ? T_38110_17_lrs2 : _GEN_19711; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19790 = 5'h11 == T_29096 ? T_38110_17_lrs3 : _GEN_19712; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19791 = 5'h11 == T_29096 ? T_38110_17_ldst_val : _GEN_19713; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19792 = 5'h11 == T_29096 ? T_38110_17_dst_rtype : _GEN_19714; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19793 = 5'h11 == T_29096 ? T_38110_17_lrs1_rtype : _GEN_19715; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19794 = 5'h11 == T_29096 ? T_38110_17_lrs2_rtype : _GEN_19716; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19795 = 5'h11 == T_29096 ? T_38110_17_frs3_en : _GEN_19717; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19796 = 5'h11 == T_29096 ? T_38110_17_fp_val : _GEN_19718; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19797 = 5'h11 == T_29096 ? T_38110_17_fp_single : _GEN_19719; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19798 = 5'h11 == T_29096 ? T_38110_17_xcpt_if : _GEN_19720; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19799 = 5'h11 == T_29096 ? T_38110_17_replay_if : _GEN_19721; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19801 = 5'h11 == T_29096 ? T_38110_17_debug_events_fetch_seq : _GEN_19723; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19802 = 5'h12 == T_29096 ? T_38110_18_valid : _GEN_19724; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19803 = 5'h12 == T_29096 ? T_38110_18_iw_state : _GEN_19725; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19804 = 5'h12 == T_29096 ? T_38110_18_uopc : _GEN_19726; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19805 = 5'h12 == T_29096 ? T_38110_18_inst : _GEN_19727; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19806 = 5'h12 == T_29096 ? T_38110_18_pc : _GEN_19728; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19807 = 5'h12 == T_29096 ? T_38110_18_fu_code : _GEN_19729; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19808 = 5'h12 == T_29096 ? T_38110_18_ctrl_br_type : _GEN_19730; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19809 = 5'h12 == T_29096 ? T_38110_18_ctrl_op1_sel : _GEN_19731; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19810 = 5'h12 == T_29096 ? T_38110_18_ctrl_op2_sel : _GEN_19732; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19811 = 5'h12 == T_29096 ? T_38110_18_ctrl_imm_sel : _GEN_19733; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19812 = 5'h12 == T_29096 ? T_38110_18_ctrl_op_fcn : _GEN_19734; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19813 = 5'h12 == T_29096 ? T_38110_18_ctrl_fcn_dw : _GEN_19735; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19814 = 5'h12 == T_29096 ? T_38110_18_ctrl_rf_wen : _GEN_19736; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19815 = 5'h12 == T_29096 ? T_38110_18_ctrl_csr_cmd : _GEN_19737; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19816 = 5'h12 == T_29096 ? T_38110_18_ctrl_is_load : _GEN_19738; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19817 = 5'h12 == T_29096 ? T_38110_18_ctrl_is_sta : _GEN_19739; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19818 = 5'h12 == T_29096 ? T_38110_18_ctrl_is_std : _GEN_19740; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19819 = 5'h12 == T_29096 ? T_38110_18_wakeup_delay : _GEN_19741; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19820 = 5'h12 == T_29096 ? T_38110_18_allocate_brtag : _GEN_19742; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19821 = 5'h12 == T_29096 ? T_38110_18_is_br_or_jmp : _GEN_19743; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19822 = 5'h12 == T_29096 ? T_38110_18_is_jump : _GEN_19744; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19823 = 5'h12 == T_29096 ? T_38110_18_is_jal : _GEN_19745; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19824 = 5'h12 == T_29096 ? T_38110_18_is_ret : _GEN_19746; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19825 = 5'h12 == T_29096 ? T_38110_18_is_call : _GEN_19747; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19826 = 5'h12 == T_29096 ? T_38110_18_br_mask : _GEN_19748; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19827 = 5'h12 == T_29096 ? T_38110_18_br_tag : _GEN_19749; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19828 = 5'h12 == T_29096 ? T_38110_18_br_prediction_bpd_predict_val : _GEN_19750; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19829 = 5'h12 == T_29096 ? T_38110_18_br_prediction_bpd_predict_taken : _GEN_19751; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19830 = 5'h12 == T_29096 ? T_38110_18_br_prediction_btb_hit : _GEN_19752; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19831 = 5'h12 == T_29096 ? T_38110_18_br_prediction_btb_predicted : _GEN_19753; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19832 = 5'h12 == T_29096 ? T_38110_18_br_prediction_is_br_or_jalr : _GEN_19754; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19833 = 5'h12 == T_29096 ? T_38110_18_stat_brjmp_mispredicted : _GEN_19755; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19834 = 5'h12 == T_29096 ? T_38110_18_stat_btb_made_pred : _GEN_19756; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19835 = 5'h12 == T_29096 ? T_38110_18_stat_btb_mispredicted : _GEN_19757; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19836 = 5'h12 == T_29096 ? T_38110_18_stat_bpd_made_pred : _GEN_19758; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19837 = 5'h12 == T_29096 ? T_38110_18_stat_bpd_mispredicted : _GEN_19759; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19838 = 5'h12 == T_29096 ? T_38110_18_fetch_pc_lob : _GEN_19760; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19839 = 5'h12 == T_29096 ? T_38110_18_imm_packed : _GEN_19761; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19840 = 5'h12 == T_29096 ? T_38110_18_csr_addr : _GEN_19762; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19841 = 5'h12 == T_29096 ? T_38110_18_rob_idx : _GEN_19763; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19842 = 5'h12 == T_29096 ? T_38110_18_ldq_idx : _GEN_19764; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19843 = 5'h12 == T_29096 ? T_38110_18_stq_idx : _GEN_19765; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19844 = 5'h12 == T_29096 ? T_38110_18_brob_idx : _GEN_19766; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19845 = 5'h12 == T_29096 ? T_38110_18_pdst : _GEN_19767; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19846 = 5'h12 == T_29096 ? T_38110_18_pop1 : _GEN_19768; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19847 = 5'h12 == T_29096 ? T_38110_18_pop2 : _GEN_19769; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19848 = 5'h12 == T_29096 ? T_38110_18_pop3 : _GEN_19770; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19849 = 5'h12 == T_29096 ? T_38110_18_prs1_busy : _GEN_19771; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19850 = 5'h12 == T_29096 ? T_38110_18_prs2_busy : _GEN_19772; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19851 = 5'h12 == T_29096 ? T_38110_18_prs3_busy : _GEN_19773; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19852 = 5'h12 == T_29096 ? T_38110_18_stale_pdst : _GEN_19774; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19853 = 5'h12 == T_29096 ? T_38110_18_exception : _GEN_19775; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19854 = 5'h12 == T_29096 ? T_38110_18_exc_cause : _GEN_19776; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19855 = 5'h12 == T_29096 ? T_38110_18_bypassable : _GEN_19777; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19856 = 5'h12 == T_29096 ? T_38110_18_mem_cmd : _GEN_19778; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19857 = 5'h12 == T_29096 ? T_38110_18_mem_typ : _GEN_19779; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19858 = 5'h12 == T_29096 ? T_38110_18_is_fence : _GEN_19780; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19859 = 5'h12 == T_29096 ? T_38110_18_is_fencei : _GEN_19781; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19860 = 5'h12 == T_29096 ? T_38110_18_is_store : _GEN_19782; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19861 = 5'h12 == T_29096 ? T_38110_18_is_amo : _GEN_19783; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19862 = 5'h12 == T_29096 ? T_38110_18_is_load : _GEN_19784; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19863 = 5'h12 == T_29096 ? T_38110_18_is_unique : _GEN_19785; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19864 = 5'h12 == T_29096 ? T_38110_18_flush_on_commit : _GEN_19786; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19865 = 5'h12 == T_29096 ? T_38110_18_ldst : _GEN_19787; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19866 = 5'h12 == T_29096 ? T_38110_18_lrs1 : _GEN_19788; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19867 = 5'h12 == T_29096 ? T_38110_18_lrs2 : _GEN_19789; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19868 = 5'h12 == T_29096 ? T_38110_18_lrs3 : _GEN_19790; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19869 = 5'h12 == T_29096 ? T_38110_18_ldst_val : _GEN_19791; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19870 = 5'h12 == T_29096 ? T_38110_18_dst_rtype : _GEN_19792; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19871 = 5'h12 == T_29096 ? T_38110_18_lrs1_rtype : _GEN_19793; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19872 = 5'h12 == T_29096 ? T_38110_18_lrs2_rtype : _GEN_19794; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19873 = 5'h12 == T_29096 ? T_38110_18_frs3_en : _GEN_19795; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19874 = 5'h12 == T_29096 ? T_38110_18_fp_val : _GEN_19796; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19875 = 5'h12 == T_29096 ? T_38110_18_fp_single : _GEN_19797; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19876 = 5'h12 == T_29096 ? T_38110_18_xcpt_if : _GEN_19798; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19877 = 5'h12 == T_29096 ? T_38110_18_replay_if : _GEN_19799; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19879 = 5'h12 == T_29096 ? T_38110_18_debug_events_fetch_seq : _GEN_19801; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19880 = 5'h13 == T_29096 ? T_38110_19_valid : _GEN_19802; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19881 = 5'h13 == T_29096 ? T_38110_19_iw_state : _GEN_19803; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19882 = 5'h13 == T_29096 ? T_38110_19_uopc : _GEN_19804; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19883 = 5'h13 == T_29096 ? T_38110_19_inst : _GEN_19805; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19884 = 5'h13 == T_29096 ? T_38110_19_pc : _GEN_19806; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19885 = 5'h13 == T_29096 ? T_38110_19_fu_code : _GEN_19807; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19886 = 5'h13 == T_29096 ? T_38110_19_ctrl_br_type : _GEN_19808; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19887 = 5'h13 == T_29096 ? T_38110_19_ctrl_op1_sel : _GEN_19809; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19888 = 5'h13 == T_29096 ? T_38110_19_ctrl_op2_sel : _GEN_19810; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19889 = 5'h13 == T_29096 ? T_38110_19_ctrl_imm_sel : _GEN_19811; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19890 = 5'h13 == T_29096 ? T_38110_19_ctrl_op_fcn : _GEN_19812; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19891 = 5'h13 == T_29096 ? T_38110_19_ctrl_fcn_dw : _GEN_19813; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19892 = 5'h13 == T_29096 ? T_38110_19_ctrl_rf_wen : _GEN_19814; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19893 = 5'h13 == T_29096 ? T_38110_19_ctrl_csr_cmd : _GEN_19815; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19894 = 5'h13 == T_29096 ? T_38110_19_ctrl_is_load : _GEN_19816; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19895 = 5'h13 == T_29096 ? T_38110_19_ctrl_is_sta : _GEN_19817; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19896 = 5'h13 == T_29096 ? T_38110_19_ctrl_is_std : _GEN_19818; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19897 = 5'h13 == T_29096 ? T_38110_19_wakeup_delay : _GEN_19819; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19898 = 5'h13 == T_29096 ? T_38110_19_allocate_brtag : _GEN_19820; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19899 = 5'h13 == T_29096 ? T_38110_19_is_br_or_jmp : _GEN_19821; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19900 = 5'h13 == T_29096 ? T_38110_19_is_jump : _GEN_19822; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19901 = 5'h13 == T_29096 ? T_38110_19_is_jal : _GEN_19823; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19902 = 5'h13 == T_29096 ? T_38110_19_is_ret : _GEN_19824; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19903 = 5'h13 == T_29096 ? T_38110_19_is_call : _GEN_19825; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19904 = 5'h13 == T_29096 ? T_38110_19_br_mask : _GEN_19826; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19905 = 5'h13 == T_29096 ? T_38110_19_br_tag : _GEN_19827; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19906 = 5'h13 == T_29096 ? T_38110_19_br_prediction_bpd_predict_val : _GEN_19828; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19907 = 5'h13 == T_29096 ? T_38110_19_br_prediction_bpd_predict_taken : _GEN_19829; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19908 = 5'h13 == T_29096 ? T_38110_19_br_prediction_btb_hit : _GEN_19830; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19909 = 5'h13 == T_29096 ? T_38110_19_br_prediction_btb_predicted : _GEN_19831; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19910 = 5'h13 == T_29096 ? T_38110_19_br_prediction_is_br_or_jalr : _GEN_19832; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19911 = 5'h13 == T_29096 ? T_38110_19_stat_brjmp_mispredicted : _GEN_19833; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19912 = 5'h13 == T_29096 ? T_38110_19_stat_btb_made_pred : _GEN_19834; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19913 = 5'h13 == T_29096 ? T_38110_19_stat_btb_mispredicted : _GEN_19835; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19914 = 5'h13 == T_29096 ? T_38110_19_stat_bpd_made_pred : _GEN_19836; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19915 = 5'h13 == T_29096 ? T_38110_19_stat_bpd_mispredicted : _GEN_19837; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19916 = 5'h13 == T_29096 ? T_38110_19_fetch_pc_lob : _GEN_19838; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19917 = 5'h13 == T_29096 ? T_38110_19_imm_packed : _GEN_19839; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19918 = 5'h13 == T_29096 ? T_38110_19_csr_addr : _GEN_19840; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19919 = 5'h13 == T_29096 ? T_38110_19_rob_idx : _GEN_19841; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19920 = 5'h13 == T_29096 ? T_38110_19_ldq_idx : _GEN_19842; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19921 = 5'h13 == T_29096 ? T_38110_19_stq_idx : _GEN_19843; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_19922 = 5'h13 == T_29096 ? T_38110_19_brob_idx : _GEN_19844; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19923 = 5'h13 == T_29096 ? T_38110_19_pdst : _GEN_19845; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19924 = 5'h13 == T_29096 ? T_38110_19_pop1 : _GEN_19846; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19925 = 5'h13 == T_29096 ? T_38110_19_pop2 : _GEN_19847; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19926 = 5'h13 == T_29096 ? T_38110_19_pop3 : _GEN_19848; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19927 = 5'h13 == T_29096 ? T_38110_19_prs1_busy : _GEN_19849; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19928 = 5'h13 == T_29096 ? T_38110_19_prs2_busy : _GEN_19850; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19929 = 5'h13 == T_29096 ? T_38110_19_prs3_busy : _GEN_19851; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_19930 = 5'h13 == T_29096 ? T_38110_19_stale_pdst : _GEN_19852; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19931 = 5'h13 == T_29096 ? T_38110_19_exception : _GEN_19853; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_19932 = 5'h13 == T_29096 ? T_38110_19_exc_cause : _GEN_19854; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19933 = 5'h13 == T_29096 ? T_38110_19_bypassable : _GEN_19855; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19934 = 5'h13 == T_29096 ? T_38110_19_mem_cmd : _GEN_19856; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19935 = 5'h13 == T_29096 ? T_38110_19_mem_typ : _GEN_19857; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19936 = 5'h13 == T_29096 ? T_38110_19_is_fence : _GEN_19858; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19937 = 5'h13 == T_29096 ? T_38110_19_is_fencei : _GEN_19859; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19938 = 5'h13 == T_29096 ? T_38110_19_is_store : _GEN_19860; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19939 = 5'h13 == T_29096 ? T_38110_19_is_amo : _GEN_19861; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19940 = 5'h13 == T_29096 ? T_38110_19_is_load : _GEN_19862; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19941 = 5'h13 == T_29096 ? T_38110_19_is_unique : _GEN_19863; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19942 = 5'h13 == T_29096 ? T_38110_19_flush_on_commit : _GEN_19864; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19943 = 5'h13 == T_29096 ? T_38110_19_ldst : _GEN_19865; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19944 = 5'h13 == T_29096 ? T_38110_19_lrs1 : _GEN_19866; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19945 = 5'h13 == T_29096 ? T_38110_19_lrs2 : _GEN_19867; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19946 = 5'h13 == T_29096 ? T_38110_19_lrs3 : _GEN_19868; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19947 = 5'h13 == T_29096 ? T_38110_19_ldst_val : _GEN_19869; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19948 = 5'h13 == T_29096 ? T_38110_19_dst_rtype : _GEN_19870; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19949 = 5'h13 == T_29096 ? T_38110_19_lrs1_rtype : _GEN_19871; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19950 = 5'h13 == T_29096 ? T_38110_19_lrs2_rtype : _GEN_19872; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19951 = 5'h13 == T_29096 ? T_38110_19_frs3_en : _GEN_19873; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19952 = 5'h13 == T_29096 ? T_38110_19_fp_val : _GEN_19874; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19953 = 5'h13 == T_29096 ? T_38110_19_fp_single : _GEN_19875; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19954 = 5'h13 == T_29096 ? T_38110_19_xcpt_if : _GEN_19876; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19955 = 5'h13 == T_29096 ? T_38110_19_replay_if : _GEN_19877; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19957 = 5'h13 == T_29096 ? T_38110_19_debug_events_fetch_seq : _GEN_19879; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19958 = 5'h14 == T_29096 ? T_38110_20_valid : _GEN_19880; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19959 = 5'h14 == T_29096 ? T_38110_20_iw_state : _GEN_19881; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_19960 = 5'h14 == T_29096 ? T_38110_20_uopc : _GEN_19882; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_19961 = 5'h14 == T_29096 ? T_38110_20_inst : _GEN_19883; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_19962 = 5'h14 == T_29096 ? T_38110_20_pc : _GEN_19884; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19963 = 5'h14 == T_29096 ? T_38110_20_fu_code : _GEN_19885; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19964 = 5'h14 == T_29096 ? T_38110_20_ctrl_br_type : _GEN_19886; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19965 = 5'h14 == T_29096 ? T_38110_20_ctrl_op1_sel : _GEN_19887; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19966 = 5'h14 == T_29096 ? T_38110_20_ctrl_op2_sel : _GEN_19888; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19967 = 5'h14 == T_29096 ? T_38110_20_ctrl_imm_sel : _GEN_19889; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19968 = 5'h14 == T_29096 ? T_38110_20_ctrl_op_fcn : _GEN_19890; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19969 = 5'h14 == T_29096 ? T_38110_20_ctrl_fcn_dw : _GEN_19891; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19970 = 5'h14 == T_29096 ? T_38110_20_ctrl_rf_wen : _GEN_19892; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19971 = 5'h14 == T_29096 ? T_38110_20_ctrl_csr_cmd : _GEN_19893; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19972 = 5'h14 == T_29096 ? T_38110_20_ctrl_is_load : _GEN_19894; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19973 = 5'h14 == T_29096 ? T_38110_20_ctrl_is_sta : _GEN_19895; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19974 = 5'h14 == T_29096 ? T_38110_20_ctrl_is_std : _GEN_19896; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_19975 = 5'h14 == T_29096 ? T_38110_20_wakeup_delay : _GEN_19897; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19976 = 5'h14 == T_29096 ? T_38110_20_allocate_brtag : _GEN_19898; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19977 = 5'h14 == T_29096 ? T_38110_20_is_br_or_jmp : _GEN_19899; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19978 = 5'h14 == T_29096 ? T_38110_20_is_jump : _GEN_19900; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19979 = 5'h14 == T_29096 ? T_38110_20_is_jal : _GEN_19901; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19980 = 5'h14 == T_29096 ? T_38110_20_is_ret : _GEN_19902; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19981 = 5'h14 == T_29096 ? T_38110_20_is_call : _GEN_19903; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_19982 = 5'h14 == T_29096 ? T_38110_20_br_mask : _GEN_19904; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19983 = 5'h14 == T_29096 ? T_38110_20_br_tag : _GEN_19905; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19984 = 5'h14 == T_29096 ? T_38110_20_br_prediction_bpd_predict_val : _GEN_19906; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19985 = 5'h14 == T_29096 ? T_38110_20_br_prediction_bpd_predict_taken : _GEN_19907; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19986 = 5'h14 == T_29096 ? T_38110_20_br_prediction_btb_hit : _GEN_19908; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19987 = 5'h14 == T_29096 ? T_38110_20_br_prediction_btb_predicted : _GEN_19909; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19988 = 5'h14 == T_29096 ? T_38110_20_br_prediction_is_br_or_jalr : _GEN_19910; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19989 = 5'h14 == T_29096 ? T_38110_20_stat_brjmp_mispredicted : _GEN_19911; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19990 = 5'h14 == T_29096 ? T_38110_20_stat_btb_made_pred : _GEN_19912; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19991 = 5'h14 == T_29096 ? T_38110_20_stat_btb_mispredicted : _GEN_19913; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19992 = 5'h14 == T_29096 ? T_38110_20_stat_bpd_made_pred : _GEN_19914; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_19993 = 5'h14 == T_29096 ? T_38110_20_stat_bpd_mispredicted : _GEN_19915; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_19994 = 5'h14 == T_29096 ? T_38110_20_fetch_pc_lob : _GEN_19916; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_19995 = 5'h14 == T_29096 ? T_38110_20_imm_packed : _GEN_19917; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_19996 = 5'h14 == T_29096 ? T_38110_20_csr_addr : _GEN_19918; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_19997 = 5'h14 == T_29096 ? T_38110_20_rob_idx : _GEN_19919; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19998 = 5'h14 == T_29096 ? T_38110_20_ldq_idx : _GEN_19920; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_19999 = 5'h14 == T_29096 ? T_38110_20_stq_idx : _GEN_19921; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_20000 = 5'h14 == T_29096 ? T_38110_20_brob_idx : _GEN_19922; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20001 = 5'h14 == T_29096 ? T_38110_20_pdst : _GEN_19923; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20002 = 5'h14 == T_29096 ? T_38110_20_pop1 : _GEN_19924; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20003 = 5'h14 == T_29096 ? T_38110_20_pop2 : _GEN_19925; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20004 = 5'h14 == T_29096 ? T_38110_20_pop3 : _GEN_19926; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20005 = 5'h14 == T_29096 ? T_38110_20_prs1_busy : _GEN_19927; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20006 = 5'h14 == T_29096 ? T_38110_20_prs2_busy : _GEN_19928; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20007 = 5'h14 == T_29096 ? T_38110_20_prs3_busy : _GEN_19929; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20008 = 5'h14 == T_29096 ? T_38110_20_stale_pdst : _GEN_19930; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20009 = 5'h14 == T_29096 ? T_38110_20_exception : _GEN_19931; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_20010 = 5'h14 == T_29096 ? T_38110_20_exc_cause : _GEN_19932; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20011 = 5'h14 == T_29096 ? T_38110_20_bypassable : _GEN_19933; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20012 = 5'h14 == T_29096 ? T_38110_20_mem_cmd : _GEN_19934; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20013 = 5'h14 == T_29096 ? T_38110_20_mem_typ : _GEN_19935; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20014 = 5'h14 == T_29096 ? T_38110_20_is_fence : _GEN_19936; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20015 = 5'h14 == T_29096 ? T_38110_20_is_fencei : _GEN_19937; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20016 = 5'h14 == T_29096 ? T_38110_20_is_store : _GEN_19938; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20017 = 5'h14 == T_29096 ? T_38110_20_is_amo : _GEN_19939; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20018 = 5'h14 == T_29096 ? T_38110_20_is_load : _GEN_19940; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20019 = 5'h14 == T_29096 ? T_38110_20_is_unique : _GEN_19941; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20020 = 5'h14 == T_29096 ? T_38110_20_flush_on_commit : _GEN_19942; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20021 = 5'h14 == T_29096 ? T_38110_20_ldst : _GEN_19943; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20022 = 5'h14 == T_29096 ? T_38110_20_lrs1 : _GEN_19944; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20023 = 5'h14 == T_29096 ? T_38110_20_lrs2 : _GEN_19945; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20024 = 5'h14 == T_29096 ? T_38110_20_lrs3 : _GEN_19946; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20025 = 5'h14 == T_29096 ? T_38110_20_ldst_val : _GEN_19947; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20026 = 5'h14 == T_29096 ? T_38110_20_dst_rtype : _GEN_19948; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20027 = 5'h14 == T_29096 ? T_38110_20_lrs1_rtype : _GEN_19949; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20028 = 5'h14 == T_29096 ? T_38110_20_lrs2_rtype : _GEN_19950; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20029 = 5'h14 == T_29096 ? T_38110_20_frs3_en : _GEN_19951; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20030 = 5'h14 == T_29096 ? T_38110_20_fp_val : _GEN_19952; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20031 = 5'h14 == T_29096 ? T_38110_20_fp_single : _GEN_19953; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20032 = 5'h14 == T_29096 ? T_38110_20_xcpt_if : _GEN_19954; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20033 = 5'h14 == T_29096 ? T_38110_20_replay_if : _GEN_19955; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_20035 = 5'h14 == T_29096 ? T_38110_20_debug_events_fetch_seq : _GEN_19957; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20036 = 5'h15 == T_29096 ? T_38110_21_valid : _GEN_19958; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20037 = 5'h15 == T_29096 ? T_38110_21_iw_state : _GEN_19959; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_20038 = 5'h15 == T_29096 ? T_38110_21_uopc : _GEN_19960; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_20039 = 5'h15 == T_29096 ? T_38110_21_inst : _GEN_19961; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_20040 = 5'h15 == T_29096 ? T_38110_21_pc : _GEN_19962; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_20041 = 5'h15 == T_29096 ? T_38110_21_fu_code : _GEN_19963; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20042 = 5'h15 == T_29096 ? T_38110_21_ctrl_br_type : _GEN_19964; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20043 = 5'h15 == T_29096 ? T_38110_21_ctrl_op1_sel : _GEN_19965; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20044 = 5'h15 == T_29096 ? T_38110_21_ctrl_op2_sel : _GEN_19966; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20045 = 5'h15 == T_29096 ? T_38110_21_ctrl_imm_sel : _GEN_19967; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20046 = 5'h15 == T_29096 ? T_38110_21_ctrl_op_fcn : _GEN_19968; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20047 = 5'h15 == T_29096 ? T_38110_21_ctrl_fcn_dw : _GEN_19969; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20048 = 5'h15 == T_29096 ? T_38110_21_ctrl_rf_wen : _GEN_19970; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20049 = 5'h15 == T_29096 ? T_38110_21_ctrl_csr_cmd : _GEN_19971; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20050 = 5'h15 == T_29096 ? T_38110_21_ctrl_is_load : _GEN_19972; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20051 = 5'h15 == T_29096 ? T_38110_21_ctrl_is_sta : _GEN_19973; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20052 = 5'h15 == T_29096 ? T_38110_21_ctrl_is_std : _GEN_19974; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20053 = 5'h15 == T_29096 ? T_38110_21_wakeup_delay : _GEN_19975; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20054 = 5'h15 == T_29096 ? T_38110_21_allocate_brtag : _GEN_19976; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20055 = 5'h15 == T_29096 ? T_38110_21_is_br_or_jmp : _GEN_19977; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20056 = 5'h15 == T_29096 ? T_38110_21_is_jump : _GEN_19978; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20057 = 5'h15 == T_29096 ? T_38110_21_is_jal : _GEN_19979; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20058 = 5'h15 == T_29096 ? T_38110_21_is_ret : _GEN_19980; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20059 = 5'h15 == T_29096 ? T_38110_21_is_call : _GEN_19981; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_20060 = 5'h15 == T_29096 ? T_38110_21_br_mask : _GEN_19982; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20061 = 5'h15 == T_29096 ? T_38110_21_br_tag : _GEN_19983; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20062 = 5'h15 == T_29096 ? T_38110_21_br_prediction_bpd_predict_val : _GEN_19984; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20063 = 5'h15 == T_29096 ? T_38110_21_br_prediction_bpd_predict_taken : _GEN_19985; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20064 = 5'h15 == T_29096 ? T_38110_21_br_prediction_btb_hit : _GEN_19986; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20065 = 5'h15 == T_29096 ? T_38110_21_br_prediction_btb_predicted : _GEN_19987; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20066 = 5'h15 == T_29096 ? T_38110_21_br_prediction_is_br_or_jalr : _GEN_19988; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20067 = 5'h15 == T_29096 ? T_38110_21_stat_brjmp_mispredicted : _GEN_19989; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20068 = 5'h15 == T_29096 ? T_38110_21_stat_btb_made_pred : _GEN_19990; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20069 = 5'h15 == T_29096 ? T_38110_21_stat_btb_mispredicted : _GEN_19991; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20070 = 5'h15 == T_29096 ? T_38110_21_stat_bpd_made_pred : _GEN_19992; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20071 = 5'h15 == T_29096 ? T_38110_21_stat_bpd_mispredicted : _GEN_19993; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20072 = 5'h15 == T_29096 ? T_38110_21_fetch_pc_lob : _GEN_19994; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_20073 = 5'h15 == T_29096 ? T_38110_21_imm_packed : _GEN_19995; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_20074 = 5'h15 == T_29096 ? T_38110_21_csr_addr : _GEN_19996; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20075 = 5'h15 == T_29096 ? T_38110_21_rob_idx : _GEN_19997; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20076 = 5'h15 == T_29096 ? T_38110_21_ldq_idx : _GEN_19998; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20077 = 5'h15 == T_29096 ? T_38110_21_stq_idx : _GEN_19999; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_20078 = 5'h15 == T_29096 ? T_38110_21_brob_idx : _GEN_20000; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20079 = 5'h15 == T_29096 ? T_38110_21_pdst : _GEN_20001; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20080 = 5'h15 == T_29096 ? T_38110_21_pop1 : _GEN_20002; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20081 = 5'h15 == T_29096 ? T_38110_21_pop2 : _GEN_20003; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20082 = 5'h15 == T_29096 ? T_38110_21_pop3 : _GEN_20004; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20083 = 5'h15 == T_29096 ? T_38110_21_prs1_busy : _GEN_20005; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20084 = 5'h15 == T_29096 ? T_38110_21_prs2_busy : _GEN_20006; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20085 = 5'h15 == T_29096 ? T_38110_21_prs3_busy : _GEN_20007; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20086 = 5'h15 == T_29096 ? T_38110_21_stale_pdst : _GEN_20008; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20087 = 5'h15 == T_29096 ? T_38110_21_exception : _GEN_20009; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_20088 = 5'h15 == T_29096 ? T_38110_21_exc_cause : _GEN_20010; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20089 = 5'h15 == T_29096 ? T_38110_21_bypassable : _GEN_20011; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20090 = 5'h15 == T_29096 ? T_38110_21_mem_cmd : _GEN_20012; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20091 = 5'h15 == T_29096 ? T_38110_21_mem_typ : _GEN_20013; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20092 = 5'h15 == T_29096 ? T_38110_21_is_fence : _GEN_20014; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20093 = 5'h15 == T_29096 ? T_38110_21_is_fencei : _GEN_20015; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20094 = 5'h15 == T_29096 ? T_38110_21_is_store : _GEN_20016; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20095 = 5'h15 == T_29096 ? T_38110_21_is_amo : _GEN_20017; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20096 = 5'h15 == T_29096 ? T_38110_21_is_load : _GEN_20018; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20097 = 5'h15 == T_29096 ? T_38110_21_is_unique : _GEN_20019; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20098 = 5'h15 == T_29096 ? T_38110_21_flush_on_commit : _GEN_20020; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20099 = 5'h15 == T_29096 ? T_38110_21_ldst : _GEN_20021; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20100 = 5'h15 == T_29096 ? T_38110_21_lrs1 : _GEN_20022; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20101 = 5'h15 == T_29096 ? T_38110_21_lrs2 : _GEN_20023; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20102 = 5'h15 == T_29096 ? T_38110_21_lrs3 : _GEN_20024; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20103 = 5'h15 == T_29096 ? T_38110_21_ldst_val : _GEN_20025; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20104 = 5'h15 == T_29096 ? T_38110_21_dst_rtype : _GEN_20026; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20105 = 5'h15 == T_29096 ? T_38110_21_lrs1_rtype : _GEN_20027; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20106 = 5'h15 == T_29096 ? T_38110_21_lrs2_rtype : _GEN_20028; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20107 = 5'h15 == T_29096 ? T_38110_21_frs3_en : _GEN_20029; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20108 = 5'h15 == T_29096 ? T_38110_21_fp_val : _GEN_20030; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20109 = 5'h15 == T_29096 ? T_38110_21_fp_single : _GEN_20031; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20110 = 5'h15 == T_29096 ? T_38110_21_xcpt_if : _GEN_20032; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20111 = 5'h15 == T_29096 ? T_38110_21_replay_if : _GEN_20033; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_20113 = 5'h15 == T_29096 ? T_38110_21_debug_events_fetch_seq : _GEN_20035; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20114 = 5'h16 == T_29096 ? T_38110_22_valid : _GEN_20036; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20115 = 5'h16 == T_29096 ? T_38110_22_iw_state : _GEN_20037; // @[rob.scala 453:59 rob.scala 453:59]
  wire [8:0] _GEN_20116 = 5'h16 == T_29096 ? T_38110_22_uopc : _GEN_20038; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_20117 = 5'h16 == T_29096 ? T_38110_22_inst : _GEN_20039; // @[rob.scala 453:59 rob.scala 453:59]
  wire [39:0] _GEN_20118 = 5'h16 == T_29096 ? T_38110_22_pc : _GEN_20040; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_20119 = 5'h16 == T_29096 ? T_38110_22_fu_code : _GEN_20041; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20120 = 5'h16 == T_29096 ? T_38110_22_ctrl_br_type : _GEN_20042; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20121 = 5'h16 == T_29096 ? T_38110_22_ctrl_op1_sel : _GEN_20043; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20122 = 5'h16 == T_29096 ? T_38110_22_ctrl_op2_sel : _GEN_20044; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20123 = 5'h16 == T_29096 ? T_38110_22_ctrl_imm_sel : _GEN_20045; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20124 = 5'h16 == T_29096 ? T_38110_22_ctrl_op_fcn : _GEN_20046; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20125 = 5'h16 == T_29096 ? T_38110_22_ctrl_fcn_dw : _GEN_20047; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20126 = 5'h16 == T_29096 ? T_38110_22_ctrl_rf_wen : _GEN_20048; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20127 = 5'h16 == T_29096 ? T_38110_22_ctrl_csr_cmd : _GEN_20049; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20128 = 5'h16 == T_29096 ? T_38110_22_ctrl_is_load : _GEN_20050; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20129 = 5'h16 == T_29096 ? T_38110_22_ctrl_is_sta : _GEN_20051; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20130 = 5'h16 == T_29096 ? T_38110_22_ctrl_is_std : _GEN_20052; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20131 = 5'h16 == T_29096 ? T_38110_22_wakeup_delay : _GEN_20053; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20132 = 5'h16 == T_29096 ? T_38110_22_allocate_brtag : _GEN_20054; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20133 = 5'h16 == T_29096 ? T_38110_22_is_br_or_jmp : _GEN_20055; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20134 = 5'h16 == T_29096 ? T_38110_22_is_jump : _GEN_20056; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20135 = 5'h16 == T_29096 ? T_38110_22_is_jal : _GEN_20057; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20136 = 5'h16 == T_29096 ? T_38110_22_is_ret : _GEN_20058; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20137 = 5'h16 == T_29096 ? T_38110_22_is_call : _GEN_20059; // @[rob.scala 453:59 rob.scala 453:59]
  wire [7:0] _GEN_20138 = 5'h16 == T_29096 ? T_38110_22_br_mask : _GEN_20060; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20139 = 5'h16 == T_29096 ? T_38110_22_br_tag : _GEN_20061; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20140 = 5'h16 == T_29096 ? T_38110_22_br_prediction_bpd_predict_val : _GEN_20062; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20141 = 5'h16 == T_29096 ? T_38110_22_br_prediction_bpd_predict_taken : _GEN_20063; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20142 = 5'h16 == T_29096 ? T_38110_22_br_prediction_btb_hit : _GEN_20064; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20143 = 5'h16 == T_29096 ? T_38110_22_br_prediction_btb_predicted : _GEN_20065; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20144 = 5'h16 == T_29096 ? T_38110_22_br_prediction_is_br_or_jalr : _GEN_20066; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20145 = 5'h16 == T_29096 ? T_38110_22_stat_brjmp_mispredicted : _GEN_20067; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20146 = 5'h16 == T_29096 ? T_38110_22_stat_btb_made_pred : _GEN_20068; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20147 = 5'h16 == T_29096 ? T_38110_22_stat_btb_mispredicted : _GEN_20069; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20148 = 5'h16 == T_29096 ? T_38110_22_stat_bpd_made_pred : _GEN_20070; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20149 = 5'h16 == T_29096 ? T_38110_22_stat_bpd_mispredicted : _GEN_20071; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20150 = 5'h16 == T_29096 ? T_38110_22_fetch_pc_lob : _GEN_20072; // @[rob.scala 453:59 rob.scala 453:59]
  wire [19:0] _GEN_20151 = 5'h16 == T_29096 ? T_38110_22_imm_packed : _GEN_20073; // @[rob.scala 453:59 rob.scala 453:59]
  wire [11:0] _GEN_20152 = 5'h16 == T_29096 ? T_38110_22_csr_addr : _GEN_20074; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20153 = 5'h16 == T_29096 ? T_38110_22_rob_idx : _GEN_20075; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20154 = 5'h16 == T_29096 ? T_38110_22_ldq_idx : _GEN_20076; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20155 = 5'h16 == T_29096 ? T_38110_22_stq_idx : _GEN_20077; // @[rob.scala 453:59 rob.scala 453:59]
  wire [4:0] _GEN_20156 = 5'h16 == T_29096 ? T_38110_22_brob_idx : _GEN_20078; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20157 = 5'h16 == T_29096 ? T_38110_22_pdst : _GEN_20079; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20158 = 5'h16 == T_29096 ? T_38110_22_pop1 : _GEN_20080; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20159 = 5'h16 == T_29096 ? T_38110_22_pop2 : _GEN_20081; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20160 = 5'h16 == T_29096 ? T_38110_22_pop3 : _GEN_20082; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20161 = 5'h16 == T_29096 ? T_38110_22_prs1_busy : _GEN_20083; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20162 = 5'h16 == T_29096 ? T_38110_22_prs2_busy : _GEN_20084; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20163 = 5'h16 == T_29096 ? T_38110_22_prs3_busy : _GEN_20085; // @[rob.scala 453:59 rob.scala 453:59]
  wire [6:0] _GEN_20164 = 5'h16 == T_29096 ? T_38110_22_stale_pdst : _GEN_20086; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20165 = 5'h16 == T_29096 ? T_38110_22_exception : _GEN_20087; // @[rob.scala 453:59 rob.scala 453:59]
  wire [63:0] _GEN_20166 = 5'h16 == T_29096 ? T_38110_22_exc_cause : _GEN_20088; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20167 = 5'h16 == T_29096 ? T_38110_22_bypassable : _GEN_20089; // @[rob.scala 453:59 rob.scala 453:59]
  wire [3:0] _GEN_20168 = 5'h16 == T_29096 ? T_38110_22_mem_cmd : _GEN_20090; // @[rob.scala 453:59 rob.scala 453:59]
  wire [2:0] _GEN_20169 = 5'h16 == T_29096 ? T_38110_22_mem_typ : _GEN_20091; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20170 = 5'h16 == T_29096 ? T_38110_22_is_fence : _GEN_20092; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20171 = 5'h16 == T_29096 ? T_38110_22_is_fencei : _GEN_20093; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20172 = 5'h16 == T_29096 ? T_38110_22_is_store : _GEN_20094; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20173 = 5'h16 == T_29096 ? T_38110_22_is_amo : _GEN_20095; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20174 = 5'h16 == T_29096 ? T_38110_22_is_load : _GEN_20096; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20175 = 5'h16 == T_29096 ? T_38110_22_is_unique : _GEN_20097; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20176 = 5'h16 == T_29096 ? T_38110_22_flush_on_commit : _GEN_20098; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20177 = 5'h16 == T_29096 ? T_38110_22_ldst : _GEN_20099; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20178 = 5'h16 == T_29096 ? T_38110_22_lrs1 : _GEN_20100; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20179 = 5'h16 == T_29096 ? T_38110_22_lrs2 : _GEN_20101; // @[rob.scala 453:59 rob.scala 453:59]
  wire [5:0] _GEN_20180 = 5'h16 == T_29096 ? T_38110_22_lrs3 : _GEN_20102; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20181 = 5'h16 == T_29096 ? T_38110_22_ldst_val : _GEN_20103; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20182 = 5'h16 == T_29096 ? T_38110_22_dst_rtype : _GEN_20104; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20183 = 5'h16 == T_29096 ? T_38110_22_lrs1_rtype : _GEN_20105; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20184 = 5'h16 == T_29096 ? T_38110_22_lrs2_rtype : _GEN_20106; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20185 = 5'h16 == T_29096 ? T_38110_22_frs3_en : _GEN_20107; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20186 = 5'h16 == T_29096 ? T_38110_22_fp_val : _GEN_20108; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20187 = 5'h16 == T_29096 ? T_38110_22_fp_single : _GEN_20109; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20188 = 5'h16 == T_29096 ? T_38110_22_xcpt_if : _GEN_20110; // @[rob.scala 453:59 rob.scala 453:59]
  wire  _GEN_20189 = 5'h16 == T_29096 ? T_38110_22_replay_if : _GEN_20111; // @[rob.scala 453:59 rob.scala 453:59]
  wire [31:0] _GEN_20191 = 5'h16 == T_29096 ? T_38110_22_debug_events_fetch_seq : _GEN_20113; // @[rob.scala 453:59 rob.scala 453:59]
  wire [1:0] _GEN_20260 = 5'h17 == T_29096 ? T_38110_23_dst_rtype : _GEN_20182; // @[rob.scala 453:59 rob.scala 453:59]
  wire  T_41113 = _GEN_20260 == 2'h0; // @[rob.scala 453:59]
  wire  T_41199 = _GEN_20260 == 2'h1; // @[rob.scala 453:100]
  wire  T_41200 = T_41113 | T_41199; // @[rob.scala 453:70]
  wire  _GEN_20270 = 5'h0 == T_29096 ? 1'h0 : _GEN_16096; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20271 = 5'h1 == T_29096 ? 1'h0 : _GEN_16097; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20272 = 5'h2 == T_29096 ? 1'h0 : _GEN_16098; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20273 = 5'h3 == T_29096 ? 1'h0 : _GEN_16099; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20274 = 5'h4 == T_29096 ? 1'h0 : _GEN_16100; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20275 = 5'h5 == T_29096 ? 1'h0 : _GEN_16101; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20276 = 5'h6 == T_29096 ? 1'h0 : _GEN_16102; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20277 = 5'h7 == T_29096 ? 1'h0 : _GEN_16103; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20278 = 5'h8 == T_29096 ? 1'h0 : _GEN_16104; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20279 = 5'h9 == T_29096 ? 1'h0 : _GEN_16105; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20280 = 5'ha == T_29096 ? 1'h0 : _GEN_16106; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20281 = 5'hb == T_29096 ? 1'h0 : _GEN_16107; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20282 = 5'hc == T_29096 ? 1'h0 : _GEN_16108; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20283 = 5'hd == T_29096 ? 1'h0 : _GEN_16109; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20284 = 5'he == T_29096 ? 1'h0 : _GEN_16110; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20285 = 5'hf == T_29096 ? 1'h0 : _GEN_16111; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20286 = 5'h10 == T_29096 ? 1'h0 : _GEN_16112; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20287 = 5'h11 == T_29096 ? 1'h0 : _GEN_16113; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20288 = 5'h12 == T_29096 ? 1'h0 : _GEN_16114; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20289 = 5'h13 == T_29096 ? 1'h0 : _GEN_16115; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20290 = 5'h14 == T_29096 ? 1'h0 : _GEN_16116; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20291 = 5'h15 == T_29096 ? 1'h0 : _GEN_16117; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20292 = 5'h16 == T_29096 ? 1'h0 : _GEN_16118; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20293 = 5'h17 == T_29096 ? 1'h0 : _GEN_16119; // @[rob.scala 459:33 rob.scala 459:33]
  wire  _GEN_20294 = T_29097 ? _GEN_20270 : _GEN_16096; // @[rob.scala 458:7]
  wire  _GEN_20295 = T_29097 ? _GEN_20271 : _GEN_16097; // @[rob.scala 458:7]
  wire  _GEN_20296 = T_29097 ? _GEN_20272 : _GEN_16098; // @[rob.scala 458:7]
  wire  _GEN_20297 = T_29097 ? _GEN_20273 : _GEN_16099; // @[rob.scala 458:7]
  wire  _GEN_20298 = T_29097 ? _GEN_20274 : _GEN_16100; // @[rob.scala 458:7]
  wire  _GEN_20299 = T_29097 ? _GEN_20275 : _GEN_16101; // @[rob.scala 458:7]
  wire  _GEN_20300 = T_29097 ? _GEN_20276 : _GEN_16102; // @[rob.scala 458:7]
  wire  _GEN_20301 = T_29097 ? _GEN_20277 : _GEN_16103; // @[rob.scala 458:7]
  wire  _GEN_20302 = T_29097 ? _GEN_20278 : _GEN_16104; // @[rob.scala 458:7]
  wire  _GEN_20303 = T_29097 ? _GEN_20279 : _GEN_16105; // @[rob.scala 458:7]
  wire  _GEN_20304 = T_29097 ? _GEN_20280 : _GEN_16106; // @[rob.scala 458:7]
  wire  _GEN_20305 = T_29097 ? _GEN_20281 : _GEN_16107; // @[rob.scala 458:7]
  wire  _GEN_20306 = T_29097 ? _GEN_20282 : _GEN_16108; // @[rob.scala 458:7]
  wire  _GEN_20307 = T_29097 ? _GEN_20283 : _GEN_16109; // @[rob.scala 458:7]
  wire  _GEN_20308 = T_29097 ? _GEN_20284 : _GEN_16110; // @[rob.scala 458:7]
  wire  _GEN_20309 = T_29097 ? _GEN_20285 : _GEN_16111; // @[rob.scala 458:7]
  wire  _GEN_20310 = T_29097 ? _GEN_20286 : _GEN_16112; // @[rob.scala 458:7]
  wire  _GEN_20311 = T_29097 ? _GEN_20287 : _GEN_16113; // @[rob.scala 458:7]
  wire  _GEN_20312 = T_29097 ? _GEN_20288 : _GEN_16114; // @[rob.scala 458:7]
  wire  _GEN_20313 = T_29097 ? _GEN_20289 : _GEN_16115; // @[rob.scala 458:7]
  wire  _GEN_20314 = T_29097 ? _GEN_20290 : _GEN_16116; // @[rob.scala 458:7]
  wire  _GEN_20315 = T_29097 ? _GEN_20291 : _GEN_16117; // @[rob.scala 458:7]
  wire  _GEN_20316 = T_29097 ? _GEN_20292 : _GEN_16118; // @[rob.scala 458:7]
  wire  _GEN_20317 = T_29097 ? _GEN_20293 : _GEN_16119; // @[rob.scala 458:7]
  wire [7:0] T_41293 = io_brinfo_mask & T_38110_0_br_mask; // @[util.scala 45:52]
  wire  T_41295 = T_41293 != 8'h0; // @[util.scala 45:60]
  wire  T_41296 = T_35634_0 & T_41295; // @[rob.scala 481:39]
  wire  T_41298 = T_29369 & T_41296; // @[rob.scala 484:56]
  wire  _GEN_20323 = T_41298 ? 1'h0 : _GEN_20294; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20324 = T_41298 ? 32'h4033 : _GEN_18047; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_41389 = T_29460 & T_41296; // @[rob.scala 489:62]
  wire  T_41391 = ~T_41298; // @[rob.scala 485:10]
  wire  T_41392 = T_41391 & T_41389; // @[rob.scala 490:10]
  wire [7:0] T_41394 = T_38110_0_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_41395 = io_brinfo_mask & T_38110_1_br_mask; // @[util.scala 45:52]
  wire  T_41397 = T_41395 != 8'h0; // @[util.scala 45:60]
  wire  T_41398 = T_35634_1 & T_41397; // @[rob.scala 481:39]
  wire  T_41400 = T_29369 & T_41398; // @[rob.scala 484:56]
  wire  _GEN_20326 = T_41400 ? 1'h0 : _GEN_20295; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20327 = T_41400 ? 32'h4033 : _GEN_18048; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_41491 = T_29460 & T_41398; // @[rob.scala 489:62]
  wire  T_41493 = ~T_41400; // @[rob.scala 485:10]
  wire  T_41494 = T_41493 & T_41491; // @[rob.scala 490:10]
  wire [7:0] T_41496 = T_38110_1_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_41497 = io_brinfo_mask & T_38110_2_br_mask; // @[util.scala 45:52]
  wire  T_41499 = T_41497 != 8'h0; // @[util.scala 45:60]
  wire  T_41500 = T_35634_2 & T_41499; // @[rob.scala 481:39]
  wire  T_41502 = T_29369 & T_41500; // @[rob.scala 484:56]
  wire  _GEN_20329 = T_41502 ? 1'h0 : _GEN_20296; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20330 = T_41502 ? 32'h4033 : _GEN_18049; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_41593 = T_29460 & T_41500; // @[rob.scala 489:62]
  wire  T_41595 = ~T_41502; // @[rob.scala 485:10]
  wire  T_41596 = T_41595 & T_41593; // @[rob.scala 490:10]
  wire [7:0] T_41598 = T_38110_2_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_41599 = io_brinfo_mask & T_38110_3_br_mask; // @[util.scala 45:52]
  wire  T_41601 = T_41599 != 8'h0; // @[util.scala 45:60]
  wire  T_41602 = T_35634_3 & T_41601; // @[rob.scala 481:39]
  wire  T_41604 = T_29369 & T_41602; // @[rob.scala 484:56]
  wire  _GEN_20332 = T_41604 ? 1'h0 : _GEN_20297; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20333 = T_41604 ? 32'h4033 : _GEN_18050; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_41695 = T_29460 & T_41602; // @[rob.scala 489:62]
  wire  T_41697 = ~T_41604; // @[rob.scala 485:10]
  wire  T_41698 = T_41697 & T_41695; // @[rob.scala 490:10]
  wire [7:0] T_41700 = T_38110_3_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_41701 = io_brinfo_mask & T_38110_4_br_mask; // @[util.scala 45:52]
  wire  T_41703 = T_41701 != 8'h0; // @[util.scala 45:60]
  wire  T_41704 = T_35634_4 & T_41703; // @[rob.scala 481:39]
  wire  T_41706 = T_29369 & T_41704; // @[rob.scala 484:56]
  wire  _GEN_20335 = T_41706 ? 1'h0 : _GEN_20298; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20336 = T_41706 ? 32'h4033 : _GEN_18051; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_41797 = T_29460 & T_41704; // @[rob.scala 489:62]
  wire  T_41799 = ~T_41706; // @[rob.scala 485:10]
  wire  T_41800 = T_41799 & T_41797; // @[rob.scala 490:10]
  wire [7:0] T_41802 = T_38110_4_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_41803 = io_brinfo_mask & T_38110_5_br_mask; // @[util.scala 45:52]
  wire  T_41805 = T_41803 != 8'h0; // @[util.scala 45:60]
  wire  T_41806 = T_35634_5 & T_41805; // @[rob.scala 481:39]
  wire  T_41808 = T_29369 & T_41806; // @[rob.scala 484:56]
  wire  _GEN_20338 = T_41808 ? 1'h0 : _GEN_20299; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20339 = T_41808 ? 32'h4033 : _GEN_18052; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_41899 = T_29460 & T_41806; // @[rob.scala 489:62]
  wire  T_41901 = ~T_41808; // @[rob.scala 485:10]
  wire  T_41902 = T_41901 & T_41899; // @[rob.scala 490:10]
  wire [7:0] T_41904 = T_38110_5_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_41905 = io_brinfo_mask & T_38110_6_br_mask; // @[util.scala 45:52]
  wire  T_41907 = T_41905 != 8'h0; // @[util.scala 45:60]
  wire  T_41908 = T_35634_6 & T_41907; // @[rob.scala 481:39]
  wire  T_41910 = T_29369 & T_41908; // @[rob.scala 484:56]
  wire  _GEN_20341 = T_41910 ? 1'h0 : _GEN_20300; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20342 = T_41910 ? 32'h4033 : _GEN_18053; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42001 = T_29460 & T_41908; // @[rob.scala 489:62]
  wire  T_42003 = ~T_41910; // @[rob.scala 485:10]
  wire  T_42004 = T_42003 & T_42001; // @[rob.scala 490:10]
  wire [7:0] T_42006 = T_38110_6_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42007 = io_brinfo_mask & T_38110_7_br_mask; // @[util.scala 45:52]
  wire  T_42009 = T_42007 != 8'h0; // @[util.scala 45:60]
  wire  T_42010 = T_35634_7 & T_42009; // @[rob.scala 481:39]
  wire  T_42012 = T_29369 & T_42010; // @[rob.scala 484:56]
  wire  _GEN_20344 = T_42012 ? 1'h0 : _GEN_20301; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20345 = T_42012 ? 32'h4033 : _GEN_18054; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42103 = T_29460 & T_42010; // @[rob.scala 489:62]
  wire  T_42105 = ~T_42012; // @[rob.scala 485:10]
  wire  T_42106 = T_42105 & T_42103; // @[rob.scala 490:10]
  wire [7:0] T_42108 = T_38110_7_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42109 = io_brinfo_mask & T_38110_8_br_mask; // @[util.scala 45:52]
  wire  T_42111 = T_42109 != 8'h0; // @[util.scala 45:60]
  wire  T_42112 = T_35634_8 & T_42111; // @[rob.scala 481:39]
  wire  T_42114 = T_29369 & T_42112; // @[rob.scala 484:56]
  wire  _GEN_20347 = T_42114 ? 1'h0 : _GEN_20302; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20348 = T_42114 ? 32'h4033 : _GEN_18055; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42205 = T_29460 & T_42112; // @[rob.scala 489:62]
  wire  T_42207 = ~T_42114; // @[rob.scala 485:10]
  wire  T_42208 = T_42207 & T_42205; // @[rob.scala 490:10]
  wire [7:0] T_42210 = T_38110_8_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42211 = io_brinfo_mask & T_38110_9_br_mask; // @[util.scala 45:52]
  wire  T_42213 = T_42211 != 8'h0; // @[util.scala 45:60]
  wire  T_42214 = T_35634_9 & T_42213; // @[rob.scala 481:39]
  wire  T_42216 = T_29369 & T_42214; // @[rob.scala 484:56]
  wire  _GEN_20350 = T_42216 ? 1'h0 : _GEN_20303; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20351 = T_42216 ? 32'h4033 : _GEN_18056; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42307 = T_29460 & T_42214; // @[rob.scala 489:62]
  wire  T_42309 = ~T_42216; // @[rob.scala 485:10]
  wire  T_42310 = T_42309 & T_42307; // @[rob.scala 490:10]
  wire [7:0] T_42312 = T_38110_9_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42313 = io_brinfo_mask & T_38110_10_br_mask; // @[util.scala 45:52]
  wire  T_42315 = T_42313 != 8'h0; // @[util.scala 45:60]
  wire  T_42316 = T_35634_10 & T_42315; // @[rob.scala 481:39]
  wire  T_42318 = T_29369 & T_42316; // @[rob.scala 484:56]
  wire  _GEN_20353 = T_42318 ? 1'h0 : _GEN_20304; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20354 = T_42318 ? 32'h4033 : _GEN_18057; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42409 = T_29460 & T_42316; // @[rob.scala 489:62]
  wire  T_42411 = ~T_42318; // @[rob.scala 485:10]
  wire  T_42412 = T_42411 & T_42409; // @[rob.scala 490:10]
  wire [7:0] T_42414 = T_38110_10_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42415 = io_brinfo_mask & T_38110_11_br_mask; // @[util.scala 45:52]
  wire  T_42417 = T_42415 != 8'h0; // @[util.scala 45:60]
  wire  T_42418 = T_35634_11 & T_42417; // @[rob.scala 481:39]
  wire  T_42420 = T_29369 & T_42418; // @[rob.scala 484:56]
  wire  _GEN_20356 = T_42420 ? 1'h0 : _GEN_20305; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20357 = T_42420 ? 32'h4033 : _GEN_18058; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42511 = T_29460 & T_42418; // @[rob.scala 489:62]
  wire  T_42513 = ~T_42420; // @[rob.scala 485:10]
  wire  T_42514 = T_42513 & T_42511; // @[rob.scala 490:10]
  wire [7:0] T_42516 = T_38110_11_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42517 = io_brinfo_mask & T_38110_12_br_mask; // @[util.scala 45:52]
  wire  T_42519 = T_42517 != 8'h0; // @[util.scala 45:60]
  wire  T_42520 = T_35634_12 & T_42519; // @[rob.scala 481:39]
  wire  T_42522 = T_29369 & T_42520; // @[rob.scala 484:56]
  wire  _GEN_20359 = T_42522 ? 1'h0 : _GEN_20306; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20360 = T_42522 ? 32'h4033 : _GEN_18059; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42613 = T_29460 & T_42520; // @[rob.scala 489:62]
  wire  T_42615 = ~T_42522; // @[rob.scala 485:10]
  wire  T_42616 = T_42615 & T_42613; // @[rob.scala 490:10]
  wire [7:0] T_42618 = T_38110_12_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42619 = io_brinfo_mask & T_38110_13_br_mask; // @[util.scala 45:52]
  wire  T_42621 = T_42619 != 8'h0; // @[util.scala 45:60]
  wire  T_42622 = T_35634_13 & T_42621; // @[rob.scala 481:39]
  wire  T_42624 = T_29369 & T_42622; // @[rob.scala 484:56]
  wire  _GEN_20362 = T_42624 ? 1'h0 : _GEN_20307; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20363 = T_42624 ? 32'h4033 : _GEN_18060; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42715 = T_29460 & T_42622; // @[rob.scala 489:62]
  wire  T_42717 = ~T_42624; // @[rob.scala 485:10]
  wire  T_42718 = T_42717 & T_42715; // @[rob.scala 490:10]
  wire [7:0] T_42720 = T_38110_13_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42721 = io_brinfo_mask & T_38110_14_br_mask; // @[util.scala 45:52]
  wire  T_42723 = T_42721 != 8'h0; // @[util.scala 45:60]
  wire  T_42724 = T_35634_14 & T_42723; // @[rob.scala 481:39]
  wire  T_42726 = T_29369 & T_42724; // @[rob.scala 484:56]
  wire  _GEN_20365 = T_42726 ? 1'h0 : _GEN_20308; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20366 = T_42726 ? 32'h4033 : _GEN_18061; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42817 = T_29460 & T_42724; // @[rob.scala 489:62]
  wire  T_42819 = ~T_42726; // @[rob.scala 485:10]
  wire  T_42820 = T_42819 & T_42817; // @[rob.scala 490:10]
  wire [7:0] T_42822 = T_38110_14_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42823 = io_brinfo_mask & T_38110_15_br_mask; // @[util.scala 45:52]
  wire  T_42825 = T_42823 != 8'h0; // @[util.scala 45:60]
  wire  T_42826 = T_35634_15 & T_42825; // @[rob.scala 481:39]
  wire  T_42828 = T_29369 & T_42826; // @[rob.scala 484:56]
  wire  _GEN_20368 = T_42828 ? 1'h0 : _GEN_20309; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20369 = T_42828 ? 32'h4033 : _GEN_18062; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_42919 = T_29460 & T_42826; // @[rob.scala 489:62]
  wire  T_42921 = ~T_42828; // @[rob.scala 485:10]
  wire  T_42922 = T_42921 & T_42919; // @[rob.scala 490:10]
  wire [7:0] T_42924 = T_38110_15_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_42925 = io_brinfo_mask & T_38110_16_br_mask; // @[util.scala 45:52]
  wire  T_42927 = T_42925 != 8'h0; // @[util.scala 45:60]
  wire  T_42928 = T_35634_16 & T_42927; // @[rob.scala 481:39]
  wire  T_42930 = T_29369 & T_42928; // @[rob.scala 484:56]
  wire  _GEN_20371 = T_42930 ? 1'h0 : _GEN_20310; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20372 = T_42930 ? 32'h4033 : _GEN_18063; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43021 = T_29460 & T_42928; // @[rob.scala 489:62]
  wire  T_43023 = ~T_42930; // @[rob.scala 485:10]
  wire  T_43024 = T_43023 & T_43021; // @[rob.scala 490:10]
  wire [7:0] T_43026 = T_38110_16_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43027 = io_brinfo_mask & T_38110_17_br_mask; // @[util.scala 45:52]
  wire  T_43029 = T_43027 != 8'h0; // @[util.scala 45:60]
  wire  T_43030 = T_35634_17 & T_43029; // @[rob.scala 481:39]
  wire  T_43032 = T_29369 & T_43030; // @[rob.scala 484:56]
  wire  _GEN_20374 = T_43032 ? 1'h0 : _GEN_20311; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20375 = T_43032 ? 32'h4033 : _GEN_18064; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43123 = T_29460 & T_43030; // @[rob.scala 489:62]
  wire  T_43125 = ~T_43032; // @[rob.scala 485:10]
  wire  T_43126 = T_43125 & T_43123; // @[rob.scala 490:10]
  wire [7:0] T_43128 = T_38110_17_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43129 = io_brinfo_mask & T_38110_18_br_mask; // @[util.scala 45:52]
  wire  T_43131 = T_43129 != 8'h0; // @[util.scala 45:60]
  wire  T_43132 = T_35634_18 & T_43131; // @[rob.scala 481:39]
  wire  T_43134 = T_29369 & T_43132; // @[rob.scala 484:56]
  wire  _GEN_20377 = T_43134 ? 1'h0 : _GEN_20312; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20378 = T_43134 ? 32'h4033 : _GEN_18065; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43225 = T_29460 & T_43132; // @[rob.scala 489:62]
  wire  T_43227 = ~T_43134; // @[rob.scala 485:10]
  wire  T_43228 = T_43227 & T_43225; // @[rob.scala 490:10]
  wire [7:0] T_43230 = T_38110_18_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43231 = io_brinfo_mask & T_38110_19_br_mask; // @[util.scala 45:52]
  wire  T_43233 = T_43231 != 8'h0; // @[util.scala 45:60]
  wire  T_43234 = T_35634_19 & T_43233; // @[rob.scala 481:39]
  wire  T_43236 = T_29369 & T_43234; // @[rob.scala 484:56]
  wire  _GEN_20380 = T_43236 ? 1'h0 : _GEN_20313; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20381 = T_43236 ? 32'h4033 : _GEN_18066; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43327 = T_29460 & T_43234; // @[rob.scala 489:62]
  wire  T_43329 = ~T_43236; // @[rob.scala 485:10]
  wire  T_43330 = T_43329 & T_43327; // @[rob.scala 490:10]
  wire [7:0] T_43332 = T_38110_19_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43333 = io_brinfo_mask & T_38110_20_br_mask; // @[util.scala 45:52]
  wire  T_43335 = T_43333 != 8'h0; // @[util.scala 45:60]
  wire  T_43336 = T_35634_20 & T_43335; // @[rob.scala 481:39]
  wire  T_43338 = T_29369 & T_43336; // @[rob.scala 484:56]
  wire  _GEN_20383 = T_43338 ? 1'h0 : _GEN_20314; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20384 = T_43338 ? 32'h4033 : _GEN_18067; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43429 = T_29460 & T_43336; // @[rob.scala 489:62]
  wire  T_43431 = ~T_43338; // @[rob.scala 485:10]
  wire  T_43432 = T_43431 & T_43429; // @[rob.scala 490:10]
  wire [7:0] T_43434 = T_38110_20_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43435 = io_brinfo_mask & T_38110_21_br_mask; // @[util.scala 45:52]
  wire  T_43437 = T_43435 != 8'h0; // @[util.scala 45:60]
  wire  T_43438 = T_35634_21 & T_43437; // @[rob.scala 481:39]
  wire  T_43440 = T_29369 & T_43438; // @[rob.scala 484:56]
  wire  _GEN_20386 = T_43440 ? 1'h0 : _GEN_20315; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20387 = T_43440 ? 32'h4033 : _GEN_18068; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43531 = T_29460 & T_43438; // @[rob.scala 489:62]
  wire  T_43533 = ~T_43440; // @[rob.scala 485:10]
  wire  T_43534 = T_43533 & T_43531; // @[rob.scala 490:10]
  wire [7:0] T_43536 = T_38110_21_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43537 = io_brinfo_mask & T_38110_22_br_mask; // @[util.scala 45:52]
  wire  T_43539 = T_43537 != 8'h0; // @[util.scala 45:60]
  wire  T_43540 = T_35634_22 & T_43539; // @[rob.scala 481:39]
  wire  T_43542 = T_29369 & T_43540; // @[rob.scala 484:56]
  wire  _GEN_20389 = T_43542 ? 1'h0 : _GEN_20316; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20390 = T_43542 ? 32'h4033 : _GEN_18069; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43633 = T_29460 & T_43540; // @[rob.scala 489:62]
  wire  T_43635 = ~T_43542; // @[rob.scala 485:10]
  wire  T_43636 = T_43635 & T_43633; // @[rob.scala 490:10]
  wire [7:0] T_43638 = T_38110_22_br_mask & T_29465; // @[rob.scala 492:44]
  wire [7:0] T_43639 = io_brinfo_mask & T_38110_23_br_mask; // @[util.scala 45:52]
  wire  T_43641 = T_43639 != 8'h0; // @[util.scala 45:60]
  wire  T_43642 = T_35634_23 & T_43641; // @[rob.scala 481:39]
  wire  T_43644 = T_29369 & T_43642; // @[rob.scala 484:56]
  wire  _GEN_20392 = T_43644 ? 1'h0 : _GEN_20317; // @[rob.scala 485:10 rob.scala 486:24]
  wire [31:0] _GEN_20393 = T_43644 ? 32'h4033 : _GEN_18070; // @[rob.scala 485:10 rob.scala 487:35]
  wire  T_43735 = T_29460 & T_43642; // @[rob.scala 489:62]
  wire  T_43737 = ~T_43644; // @[rob.scala 485:10]
  wire  T_43738 = T_43737 & T_43735; // @[rob.scala 490:10]
  wire [7:0] T_43740 = T_38110_23_br_mask & T_29465; // @[rob.scala 492:44]
  wire  _GEN_20579 = 5'h1 == rob_head ? T_38110_1_is_store : T_38110_0_is_store; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20581 = 5'h1 == rob_head ? T_38110_1_is_load : T_38110_0_is_load; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_20597 = 5'h1 == rob_head ? T_38110_1_debug_wdata : T_38110_0_debug_wdata; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20657 = 5'h2 == rob_head ? T_38110_2_is_store : _GEN_20579; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20659 = 5'h2 == rob_head ? T_38110_2_is_load : _GEN_20581; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_20675 = 5'h2 == rob_head ? T_38110_2_debug_wdata : _GEN_20597; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20735 = 5'h3 == rob_head ? T_38110_3_is_store : _GEN_20657; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20737 = 5'h3 == rob_head ? T_38110_3_is_load : _GEN_20659; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_20753 = 5'h3 == rob_head ? T_38110_3_debug_wdata : _GEN_20675; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20813 = 5'h4 == rob_head ? T_38110_4_is_store : _GEN_20735; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20815 = 5'h4 == rob_head ? T_38110_4_is_load : _GEN_20737; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_20831 = 5'h4 == rob_head ? T_38110_4_debug_wdata : _GEN_20753; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20891 = 5'h5 == rob_head ? T_38110_5_is_store : _GEN_20813; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20893 = 5'h5 == rob_head ? T_38110_5_is_load : _GEN_20815; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_20909 = 5'h5 == rob_head ? T_38110_5_debug_wdata : _GEN_20831; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20969 = 5'h6 == rob_head ? T_38110_6_is_store : _GEN_20891; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_20971 = 5'h6 == rob_head ? T_38110_6_is_load : _GEN_20893; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_20987 = 5'h6 == rob_head ? T_38110_6_debug_wdata : _GEN_20909; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21047 = 5'h7 == rob_head ? T_38110_7_is_store : _GEN_20969; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21049 = 5'h7 == rob_head ? T_38110_7_is_load : _GEN_20971; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21065 = 5'h7 == rob_head ? T_38110_7_debug_wdata : _GEN_20987; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21125 = 5'h8 == rob_head ? T_38110_8_is_store : _GEN_21047; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21127 = 5'h8 == rob_head ? T_38110_8_is_load : _GEN_21049; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21143 = 5'h8 == rob_head ? T_38110_8_debug_wdata : _GEN_21065; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21203 = 5'h9 == rob_head ? T_38110_9_is_store : _GEN_21125; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21205 = 5'h9 == rob_head ? T_38110_9_is_load : _GEN_21127; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21221 = 5'h9 == rob_head ? T_38110_9_debug_wdata : _GEN_21143; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21281 = 5'ha == rob_head ? T_38110_10_is_store : _GEN_21203; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21283 = 5'ha == rob_head ? T_38110_10_is_load : _GEN_21205; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21299 = 5'ha == rob_head ? T_38110_10_debug_wdata : _GEN_21221; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21359 = 5'hb == rob_head ? T_38110_11_is_store : _GEN_21281; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21361 = 5'hb == rob_head ? T_38110_11_is_load : _GEN_21283; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21377 = 5'hb == rob_head ? T_38110_11_debug_wdata : _GEN_21299; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21437 = 5'hc == rob_head ? T_38110_12_is_store : _GEN_21359; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21439 = 5'hc == rob_head ? T_38110_12_is_load : _GEN_21361; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21455 = 5'hc == rob_head ? T_38110_12_debug_wdata : _GEN_21377; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21515 = 5'hd == rob_head ? T_38110_13_is_store : _GEN_21437; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21517 = 5'hd == rob_head ? T_38110_13_is_load : _GEN_21439; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21533 = 5'hd == rob_head ? T_38110_13_debug_wdata : _GEN_21455; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21593 = 5'he == rob_head ? T_38110_14_is_store : _GEN_21515; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21595 = 5'he == rob_head ? T_38110_14_is_load : _GEN_21517; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21611 = 5'he == rob_head ? T_38110_14_debug_wdata : _GEN_21533; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21671 = 5'hf == rob_head ? T_38110_15_is_store : _GEN_21593; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21673 = 5'hf == rob_head ? T_38110_15_is_load : _GEN_21595; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21689 = 5'hf == rob_head ? T_38110_15_debug_wdata : _GEN_21611; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21749 = 5'h10 == rob_head ? T_38110_16_is_store : _GEN_21671; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21751 = 5'h10 == rob_head ? T_38110_16_is_load : _GEN_21673; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21767 = 5'h10 == rob_head ? T_38110_16_debug_wdata : _GEN_21689; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21827 = 5'h11 == rob_head ? T_38110_17_is_store : _GEN_21749; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21829 = 5'h11 == rob_head ? T_38110_17_is_load : _GEN_21751; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21845 = 5'h11 == rob_head ? T_38110_17_debug_wdata : _GEN_21767; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21905 = 5'h12 == rob_head ? T_38110_18_is_store : _GEN_21827; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21907 = 5'h12 == rob_head ? T_38110_18_is_load : _GEN_21829; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_21923 = 5'h12 == rob_head ? T_38110_18_debug_wdata : _GEN_21845; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21983 = 5'h13 == rob_head ? T_38110_19_is_store : _GEN_21905; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_21985 = 5'h13 == rob_head ? T_38110_19_is_load : _GEN_21907; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_22001 = 5'h13 == rob_head ? T_38110_19_debug_wdata : _GEN_21923; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_22061 = 5'h14 == rob_head ? T_38110_20_is_store : _GEN_21983; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_22063 = 5'h14 == rob_head ? T_38110_20_is_load : _GEN_21985; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_22079 = 5'h14 == rob_head ? T_38110_20_debug_wdata : _GEN_22001; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_22139 = 5'h15 == rob_head ? T_38110_21_is_store : _GEN_22061; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_22141 = 5'h15 == rob_head ? T_38110_21_is_load : _GEN_22063; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_22157 = 5'h15 == rob_head ? T_38110_21_debug_wdata : _GEN_22079; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_22217 = 5'h16 == rob_head ? T_38110_22_is_store : _GEN_22139; // @[rob.scala 507:28 rob.scala 507:28]
  wire  _GEN_22219 = 5'h16 == rob_head ? T_38110_22_is_load : _GEN_22141; // @[rob.scala 507:28 rob.scala 507:28]
  wire [63:0] _GEN_22235 = 5'h16 == rob_head ? T_38110_22_debug_wdata : _GEN_22157; // @[rob.scala 507:28 rob.scala 507:28]
  wire  rob_head_is_store_1 = 5'h17 == rob_head ? T_38110_23_is_store : _GEN_22217; // @[rob.scala 507:28 rob.scala 507:28]
  wire  rob_head_is_load_1 = 5'h17 == rob_head ? T_38110_23_is_load : _GEN_22219; // @[rob.scala 507:28 rob.scala 507:28]
  wire [31:0] _GEN_22339 = 5'h0 == rob_head ? 32'h4033 : _GEN_20324; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22340 = 5'h1 == rob_head ? 32'h4033 : _GEN_20327; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22341 = 5'h2 == rob_head ? 32'h4033 : _GEN_20330; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22342 = 5'h3 == rob_head ? 32'h4033 : _GEN_20333; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22343 = 5'h4 == rob_head ? 32'h4033 : _GEN_20336; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22344 = 5'h5 == rob_head ? 32'h4033 : _GEN_20339; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22345 = 5'h6 == rob_head ? 32'h4033 : _GEN_20342; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22346 = 5'h7 == rob_head ? 32'h4033 : _GEN_20345; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22347 = 5'h8 == rob_head ? 32'h4033 : _GEN_20348; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22348 = 5'h9 == rob_head ? 32'h4033 : _GEN_20351; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22349 = 5'ha == rob_head ? 32'h4033 : _GEN_20354; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22350 = 5'hb == rob_head ? 32'h4033 : _GEN_20357; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22351 = 5'hc == rob_head ? 32'h4033 : _GEN_20360; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22352 = 5'hd == rob_head ? 32'h4033 : _GEN_20363; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22353 = 5'he == rob_head ? 32'h4033 : _GEN_20366; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22354 = 5'hf == rob_head ? 32'h4033 : _GEN_20369; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22355 = 5'h10 == rob_head ? 32'h4033 : _GEN_20372; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22356 = 5'h11 == rob_head ? 32'h4033 : _GEN_20375; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22357 = 5'h12 == rob_head ? 32'h4033 : _GEN_20378; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22358 = 5'h13 == rob_head ? 32'h4033 : _GEN_20381; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22359 = 5'h14 == rob_head ? 32'h4033 : _GEN_20384; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22360 = 5'h15 == rob_head ? 32'h4033 : _GEN_20387; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22361 = 5'h16 == rob_head ? 32'h4033 : _GEN_20390; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22362 = 5'h17 == rob_head ? 32'h4033 : _GEN_20393; // @[rob.scala 515:33 rob.scala 515:33]
  wire [31:0] _GEN_22363 = T_47563 ? _GEN_22339 : _GEN_20324; // @[rob.scala 514:7]
  wire [31:0] _GEN_22364 = T_47563 ? _GEN_22340 : _GEN_20327; // @[rob.scala 514:7]
  wire [31:0] _GEN_22365 = T_47563 ? _GEN_22341 : _GEN_20330; // @[rob.scala 514:7]
  wire [31:0] _GEN_22366 = T_47563 ? _GEN_22342 : _GEN_20333; // @[rob.scala 514:7]
  wire [31:0] _GEN_22367 = T_47563 ? _GEN_22343 : _GEN_20336; // @[rob.scala 514:7]
  wire [31:0] _GEN_22368 = T_47563 ? _GEN_22344 : _GEN_20339; // @[rob.scala 514:7]
  wire [31:0] _GEN_22369 = T_47563 ? _GEN_22345 : _GEN_20342; // @[rob.scala 514:7]
  wire [31:0] _GEN_22370 = T_47563 ? _GEN_22346 : _GEN_20345; // @[rob.scala 514:7]
  wire [31:0] _GEN_22371 = T_47563 ? _GEN_22347 : _GEN_20348; // @[rob.scala 514:7]
  wire [31:0] _GEN_22372 = T_47563 ? _GEN_22348 : _GEN_20351; // @[rob.scala 514:7]
  wire [31:0] _GEN_22373 = T_47563 ? _GEN_22349 : _GEN_20354; // @[rob.scala 514:7]
  wire [31:0] _GEN_22374 = T_47563 ? _GEN_22350 : _GEN_20357; // @[rob.scala 514:7]
  wire [31:0] _GEN_22375 = T_47563 ? _GEN_22351 : _GEN_20360; // @[rob.scala 514:7]
  wire [31:0] _GEN_22376 = T_47563 ? _GEN_22352 : _GEN_20363; // @[rob.scala 514:7]
  wire [31:0] _GEN_22377 = T_47563 ? _GEN_22353 : _GEN_20366; // @[rob.scala 514:7]
  wire [31:0] _GEN_22378 = T_47563 ? _GEN_22354 : _GEN_20369; // @[rob.scala 514:7]
  wire [31:0] _GEN_22379 = T_47563 ? _GEN_22355 : _GEN_20372; // @[rob.scala 514:7]
  wire [31:0] _GEN_22380 = T_47563 ? _GEN_22356 : _GEN_20375; // @[rob.scala 514:7]
  wire [31:0] _GEN_22381 = T_47563 ? _GEN_22357 : _GEN_20378; // @[rob.scala 514:7]
  wire [31:0] _GEN_22382 = T_47563 ? _GEN_22358 : _GEN_20381; // @[rob.scala 514:7]
  wire [31:0] _GEN_22383 = T_47563 ? _GEN_22359 : _GEN_20384; // @[rob.scala 514:7]
  wire [31:0] _GEN_22384 = T_47563 ? _GEN_22360 : _GEN_20387; // @[rob.scala 514:7]
  wire [31:0] _GEN_22385 = T_47563 ? _GEN_22361 : _GEN_20390; // @[rob.scala 514:7]
  wire [31:0] _GEN_22386 = T_47563 ? _GEN_22362 : _GEN_20393; // @[rob.scala 514:7]
  wire  T_44009 = ~T_47563; // @[rob.scala 514:7]
  wire  T_44010 = T_44009 & T_29097; // @[rob.scala 518:7]
  wire  T_44099 = io_debug_wb_valids_0 & T_28590; // @[rob.scala 529:38]
  wire [63:0] _GEN_22435 = 6'h0 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17949; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22436 = 6'h1 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17950; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22437 = 6'h2 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17951; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22438 = 6'h3 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17952; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22439 = 6'h4 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17953; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22440 = 6'h5 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17954; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22441 = 6'h6 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17955; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22442 = 6'h7 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17956; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22443 = 6'h8 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17957; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22444 = 6'h9 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17958; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22445 = 6'ha == T_28589 ? io_debug_wb_wdata_0 : _GEN_17959; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22446 = 6'hb == T_28589 ? io_debug_wb_wdata_0 : _GEN_17960; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22447 = 6'hc == T_28589 ? io_debug_wb_wdata_0 : _GEN_17961; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22448 = 6'hd == T_28589 ? io_debug_wb_wdata_0 : _GEN_17962; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22449 = 6'he == T_28589 ? io_debug_wb_wdata_0 : _GEN_17963; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22450 = 6'hf == T_28589 ? io_debug_wb_wdata_0 : _GEN_17964; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22451 = 6'h10 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17965; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22452 = 6'h11 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17966; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22453 = 6'h12 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17967; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22454 = 6'h13 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17968; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22455 = 6'h14 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17969; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22456 = 6'h15 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17970; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22457 = 6'h16 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17971; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22458 = 6'h17 == T_28589 ? io_debug_wb_wdata_0 : _GEN_17972; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_22459 = T_44099 ? _GEN_22435 : _GEN_17949; // @[rob.scala 530:10]
  wire [63:0] _GEN_22460 = T_44099 ? _GEN_22436 : _GEN_17950; // @[rob.scala 530:10]
  wire [63:0] _GEN_22461 = T_44099 ? _GEN_22437 : _GEN_17951; // @[rob.scala 530:10]
  wire [63:0] _GEN_22462 = T_44099 ? _GEN_22438 : _GEN_17952; // @[rob.scala 530:10]
  wire [63:0] _GEN_22463 = T_44099 ? _GEN_22439 : _GEN_17953; // @[rob.scala 530:10]
  wire [63:0] _GEN_22464 = T_44099 ? _GEN_22440 : _GEN_17954; // @[rob.scala 530:10]
  wire [63:0] _GEN_22465 = T_44099 ? _GEN_22441 : _GEN_17955; // @[rob.scala 530:10]
  wire [63:0] _GEN_22466 = T_44099 ? _GEN_22442 : _GEN_17956; // @[rob.scala 530:10]
  wire [63:0] _GEN_22467 = T_44099 ? _GEN_22443 : _GEN_17957; // @[rob.scala 530:10]
  wire [63:0] _GEN_22468 = T_44099 ? _GEN_22444 : _GEN_17958; // @[rob.scala 530:10]
  wire [63:0] _GEN_22469 = T_44099 ? _GEN_22445 : _GEN_17959; // @[rob.scala 530:10]
  wire [63:0] _GEN_22470 = T_44099 ? _GEN_22446 : _GEN_17960; // @[rob.scala 530:10]
  wire [63:0] _GEN_22471 = T_44099 ? _GEN_22447 : _GEN_17961; // @[rob.scala 530:10]
  wire [63:0] _GEN_22472 = T_44099 ? _GEN_22448 : _GEN_17962; // @[rob.scala 530:10]
  wire [63:0] _GEN_22473 = T_44099 ? _GEN_22449 : _GEN_17963; // @[rob.scala 530:10]
  wire [63:0] _GEN_22474 = T_44099 ? _GEN_22450 : _GEN_17964; // @[rob.scala 530:10]
  wire [63:0] _GEN_22475 = T_44099 ? _GEN_22451 : _GEN_17965; // @[rob.scala 530:10]
  wire [63:0] _GEN_22476 = T_44099 ? _GEN_22452 : _GEN_17966; // @[rob.scala 530:10]
  wire [63:0] _GEN_22477 = T_44099 ? _GEN_22453 : _GEN_17967; // @[rob.scala 530:10]
  wire [63:0] _GEN_22478 = T_44099 ? _GEN_22454 : _GEN_17968; // @[rob.scala 530:10]
  wire [63:0] _GEN_22479 = T_44099 ? _GEN_22455 : _GEN_17969; // @[rob.scala 530:10]
  wire [63:0] _GEN_22480 = T_44099 ? _GEN_22456 : _GEN_17970; // @[rob.scala 530:10]
  wire [63:0] _GEN_22481 = T_44099 ? _GEN_22457 : _GEN_17971; // @[rob.scala 530:10]
  wire [63:0] _GEN_22482 = T_44099 ? _GEN_22458 : _GEN_17972; // @[rob.scala 530:10]
  wire  _GEN_22484 = 6'h1 == T_28589 ? T_35634_1 : T_35634_0; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22485 = 6'h2 == T_28589 ? T_35634_2 : _GEN_22484; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22486 = 6'h3 == T_28589 ? T_35634_3 : _GEN_22485; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22487 = 6'h4 == T_28589 ? T_35634_4 : _GEN_22486; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22488 = 6'h5 == T_28589 ? T_35634_5 : _GEN_22487; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22489 = 6'h6 == T_28589 ? T_35634_6 : _GEN_22488; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22490 = 6'h7 == T_28589 ? T_35634_7 : _GEN_22489; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22491 = 6'h8 == T_28589 ? T_35634_8 : _GEN_22490; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22492 = 6'h9 == T_28589 ? T_35634_9 : _GEN_22491; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22493 = 6'ha == T_28589 ? T_35634_10 : _GEN_22492; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22494 = 6'hb == T_28589 ? T_35634_11 : _GEN_22493; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22495 = 6'hc == T_28589 ? T_35634_12 : _GEN_22494; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22496 = 6'hd == T_28589 ? T_35634_13 : _GEN_22495; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22497 = 6'he == T_28589 ? T_35634_14 : _GEN_22496; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22498 = 6'hf == T_28589 ? T_35634_15 : _GEN_22497; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22499 = 6'h10 == T_28589 ? T_35634_16 : _GEN_22498; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22500 = 6'h11 == T_28589 ? T_35634_17 : _GEN_22499; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22501 = 6'h12 == T_28589 ? T_35634_18 : _GEN_22500; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22502 = 6'h13 == T_28589 ? T_35634_19 : _GEN_22501; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22503 = 6'h14 == T_28589 ? T_35634_20 : _GEN_22502; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22504 = 6'h15 == T_28589 ? T_35634_21 : _GEN_22503; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22505 = 6'h16 == T_28589 ? T_35634_22 : _GEN_22504; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_22506 = 6'h17 == T_28589 ? T_35634_23 : _GEN_22505; // @[rob.scala 536:22 rob.scala 536:22]
  wire  T_44281 = ~_GEN_22506; // @[rob.scala 536:22]
  wire  T_44282 = T_40521 & T_44281; // @[rob.scala 535:75]
  wire  T_44284 = ~T_44282; // @[rob.scala 535:18]
  wire  T_44285 = T_44284 | reset; // @[rob.scala 535:17]
  wire  T_44287 = ~T_44285; // @[rob.scala 535:17]
  wire [6:0] _GEN_22628 = 6'h1 == T_28589 ? T_38110_1_pdst : T_38110_0_pdst; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_22652 = 6'h1 == T_28589 ? T_38110_1_ldst_val : T_38110_0_ldst_val; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_22706 = 6'h2 == T_28589 ? T_38110_2_pdst : _GEN_22628; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_22730 = 6'h2 == T_28589 ? T_38110_2_ldst_val : _GEN_22652; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_22784 = 6'h3 == T_28589 ? T_38110_3_pdst : _GEN_22706; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_22808 = 6'h3 == T_28589 ? T_38110_3_ldst_val : _GEN_22730; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_22862 = 6'h4 == T_28589 ? T_38110_4_pdst : _GEN_22784; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_22886 = 6'h4 == T_28589 ? T_38110_4_ldst_val : _GEN_22808; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_22940 = 6'h5 == T_28589 ? T_38110_5_pdst : _GEN_22862; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_22964 = 6'h5 == T_28589 ? T_38110_5_ldst_val : _GEN_22886; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23018 = 6'h6 == T_28589 ? T_38110_6_pdst : _GEN_22940; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23042 = 6'h6 == T_28589 ? T_38110_6_ldst_val : _GEN_22964; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23096 = 6'h7 == T_28589 ? T_38110_7_pdst : _GEN_23018; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23120 = 6'h7 == T_28589 ? T_38110_7_ldst_val : _GEN_23042; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23174 = 6'h8 == T_28589 ? T_38110_8_pdst : _GEN_23096; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23198 = 6'h8 == T_28589 ? T_38110_8_ldst_val : _GEN_23120; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23252 = 6'h9 == T_28589 ? T_38110_9_pdst : _GEN_23174; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23276 = 6'h9 == T_28589 ? T_38110_9_ldst_val : _GEN_23198; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23330 = 6'ha == T_28589 ? T_38110_10_pdst : _GEN_23252; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23354 = 6'ha == T_28589 ? T_38110_10_ldst_val : _GEN_23276; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23408 = 6'hb == T_28589 ? T_38110_11_pdst : _GEN_23330; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23432 = 6'hb == T_28589 ? T_38110_11_ldst_val : _GEN_23354; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23486 = 6'hc == T_28589 ? T_38110_12_pdst : _GEN_23408; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23510 = 6'hc == T_28589 ? T_38110_12_ldst_val : _GEN_23432; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23564 = 6'hd == T_28589 ? T_38110_13_pdst : _GEN_23486; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23588 = 6'hd == T_28589 ? T_38110_13_ldst_val : _GEN_23510; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23642 = 6'he == T_28589 ? T_38110_14_pdst : _GEN_23564; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23666 = 6'he == T_28589 ? T_38110_14_ldst_val : _GEN_23588; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23720 = 6'hf == T_28589 ? T_38110_15_pdst : _GEN_23642; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23744 = 6'hf == T_28589 ? T_38110_15_ldst_val : _GEN_23666; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23798 = 6'h10 == T_28589 ? T_38110_16_pdst : _GEN_23720; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23822 = 6'h10 == T_28589 ? T_38110_16_ldst_val : _GEN_23744; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23876 = 6'h11 == T_28589 ? T_38110_17_pdst : _GEN_23798; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23900 = 6'h11 == T_28589 ? T_38110_17_ldst_val : _GEN_23822; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_23954 = 6'h12 == T_28589 ? T_38110_18_pdst : _GEN_23876; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_23978 = 6'h12 == T_28589 ? T_38110_18_ldst_val : _GEN_23900; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24032 = 6'h13 == T_28589 ? T_38110_19_pdst : _GEN_23954; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24056 = 6'h13 == T_28589 ? T_38110_19_ldst_val : _GEN_23978; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24110 = 6'h14 == T_28589 ? T_38110_20_pdst : _GEN_24032; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24134 = 6'h14 == T_28589 ? T_38110_20_ldst_val : _GEN_24056; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24188 = 6'h15 == T_28589 ? T_38110_21_pdst : _GEN_24110; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24212 = 6'h15 == T_28589 ? T_38110_21_ldst_val : _GEN_24134; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24266 = 6'h16 == T_28589 ? T_38110_22_pdst : _GEN_24188; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24290 = 6'h16 == T_28589 ? T_38110_22_ldst_val : _GEN_24212; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24344 = 6'h17 == T_28589 ? T_38110_23_pdst : _GEN_24266; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24368 = 6'h17 == T_28589 ? T_38110_23_ldst_val : _GEN_24290; // @[rob.scala 538:75 rob.scala 538:75]
  wire  T_44292 = T_40521 & _GEN_24368; // @[rob.scala 538:75]
  wire  T_44293 = _GEN_24344 != io_wb_resps_0_bits_uop_pdst; // @[rob.scala 539:54]
  wire  T_44294 = T_44292 & T_44293; // @[rob.scala 539:37]
  wire  T_44296 = ~T_44294; // @[rob.scala 538:18]
  wire  T_44297 = T_44296 | reset; // @[rob.scala 538:17]
  wire  T_44299 = ~T_44297; // @[rob.scala 538:17]
  wire  T_44303 = io_debug_wb_valids_1 & T_28598; // @[rob.scala 529:38]
  wire [63:0] _GEN_24379 = 6'h0 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22459; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24380 = 6'h1 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22460; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24381 = 6'h2 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22461; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24382 = 6'h3 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22462; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24383 = 6'h4 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22463; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24384 = 6'h5 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22464; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24385 = 6'h6 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22465; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24386 = 6'h7 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22466; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24387 = 6'h8 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22467; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24388 = 6'h9 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22468; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24389 = 6'ha == T_28597 ? io_debug_wb_wdata_1 : _GEN_22469; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24390 = 6'hb == T_28597 ? io_debug_wb_wdata_1 : _GEN_22470; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24391 = 6'hc == T_28597 ? io_debug_wb_wdata_1 : _GEN_22471; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24392 = 6'hd == T_28597 ? io_debug_wb_wdata_1 : _GEN_22472; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24393 = 6'he == T_28597 ? io_debug_wb_wdata_1 : _GEN_22473; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24394 = 6'hf == T_28597 ? io_debug_wb_wdata_1 : _GEN_22474; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24395 = 6'h10 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22475; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24396 = 6'h11 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22476; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24397 = 6'h12 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22477; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24398 = 6'h13 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22478; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24399 = 6'h14 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22479; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24400 = 6'h15 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22480; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24401 = 6'h16 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22481; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24402 = 6'h17 == T_28597 ? io_debug_wb_wdata_1 : _GEN_22482; // @[rob.scala 531:53 rob.scala 531:53]
  wire [63:0] _GEN_24403 = T_44303 ? _GEN_24379 : _GEN_22459; // @[rob.scala 530:10]
  wire [63:0] _GEN_24404 = T_44303 ? _GEN_24380 : _GEN_22460; // @[rob.scala 530:10]
  wire [63:0] _GEN_24405 = T_44303 ? _GEN_24381 : _GEN_22461; // @[rob.scala 530:10]
  wire [63:0] _GEN_24406 = T_44303 ? _GEN_24382 : _GEN_22462; // @[rob.scala 530:10]
  wire [63:0] _GEN_24407 = T_44303 ? _GEN_24383 : _GEN_22463; // @[rob.scala 530:10]
  wire [63:0] _GEN_24408 = T_44303 ? _GEN_24384 : _GEN_22464; // @[rob.scala 530:10]
  wire [63:0] _GEN_24409 = T_44303 ? _GEN_24385 : _GEN_22465; // @[rob.scala 530:10]
  wire [63:0] _GEN_24410 = T_44303 ? _GEN_24386 : _GEN_22466; // @[rob.scala 530:10]
  wire [63:0] _GEN_24411 = T_44303 ? _GEN_24387 : _GEN_22467; // @[rob.scala 530:10]
  wire [63:0] _GEN_24412 = T_44303 ? _GEN_24388 : _GEN_22468; // @[rob.scala 530:10]
  wire [63:0] _GEN_24413 = T_44303 ? _GEN_24389 : _GEN_22469; // @[rob.scala 530:10]
  wire [63:0] _GEN_24414 = T_44303 ? _GEN_24390 : _GEN_22470; // @[rob.scala 530:10]
  wire [63:0] _GEN_24415 = T_44303 ? _GEN_24391 : _GEN_22471; // @[rob.scala 530:10]
  wire [63:0] _GEN_24416 = T_44303 ? _GEN_24392 : _GEN_22472; // @[rob.scala 530:10]
  wire [63:0] _GEN_24417 = T_44303 ? _GEN_24393 : _GEN_22473; // @[rob.scala 530:10]
  wire [63:0] _GEN_24418 = T_44303 ? _GEN_24394 : _GEN_22474; // @[rob.scala 530:10]
  wire [63:0] _GEN_24419 = T_44303 ? _GEN_24395 : _GEN_22475; // @[rob.scala 530:10]
  wire [63:0] _GEN_24420 = T_44303 ? _GEN_24396 : _GEN_22476; // @[rob.scala 530:10]
  wire [63:0] _GEN_24421 = T_44303 ? _GEN_24397 : _GEN_22477; // @[rob.scala 530:10]
  wire [63:0] _GEN_24422 = T_44303 ? _GEN_24398 : _GEN_22478; // @[rob.scala 530:10]
  wire [63:0] _GEN_24423 = T_44303 ? _GEN_24399 : _GEN_22479; // @[rob.scala 530:10]
  wire [63:0] _GEN_24424 = T_44303 ? _GEN_24400 : _GEN_22480; // @[rob.scala 530:10]
  wire [63:0] _GEN_24425 = T_44303 ? _GEN_24401 : _GEN_22481; // @[rob.scala 530:10]
  wire [63:0] _GEN_24426 = T_44303 ? _GEN_24402 : _GEN_22482; // @[rob.scala 530:10]
  wire  _GEN_24428 = 6'h1 == T_28597 ? T_35634_1 : T_35634_0; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24429 = 6'h2 == T_28597 ? T_35634_2 : _GEN_24428; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24430 = 6'h3 == T_28597 ? T_35634_3 : _GEN_24429; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24431 = 6'h4 == T_28597 ? T_35634_4 : _GEN_24430; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24432 = 6'h5 == T_28597 ? T_35634_5 : _GEN_24431; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24433 = 6'h6 == T_28597 ? T_35634_6 : _GEN_24432; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24434 = 6'h7 == T_28597 ? T_35634_7 : _GEN_24433; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24435 = 6'h8 == T_28597 ? T_35634_8 : _GEN_24434; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24436 = 6'h9 == T_28597 ? T_35634_9 : _GEN_24435; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24437 = 6'ha == T_28597 ? T_35634_10 : _GEN_24436; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24438 = 6'hb == T_28597 ? T_35634_11 : _GEN_24437; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24439 = 6'hc == T_28597 ? T_35634_12 : _GEN_24438; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24440 = 6'hd == T_28597 ? T_35634_13 : _GEN_24439; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24441 = 6'he == T_28597 ? T_35634_14 : _GEN_24440; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24442 = 6'hf == T_28597 ? T_35634_15 : _GEN_24441; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24443 = 6'h10 == T_28597 ? T_35634_16 : _GEN_24442; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24444 = 6'h11 == T_28597 ? T_35634_17 : _GEN_24443; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24445 = 6'h12 == T_28597 ? T_35634_18 : _GEN_24444; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24446 = 6'h13 == T_28597 ? T_35634_19 : _GEN_24445; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24447 = 6'h14 == T_28597 ? T_35634_20 : _GEN_24446; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24448 = 6'h15 == T_28597 ? T_35634_21 : _GEN_24447; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24449 = 6'h16 == T_28597 ? T_35634_22 : _GEN_24448; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_24450 = 6'h17 == T_28597 ? T_35634_23 : _GEN_24449; // @[rob.scala 536:22 rob.scala 536:22]
  wire  T_44485 = ~_GEN_24450; // @[rob.scala 536:22]
  wire  T_44486 = T_40529 & T_44485; // @[rob.scala 535:75]
  wire  T_44488 = ~T_44486; // @[rob.scala 535:18]
  wire  T_44489 = T_44488 | reset; // @[rob.scala 535:17]
  wire  T_44491 = ~T_44489; // @[rob.scala 535:17]
  wire [6:0] _GEN_24572 = 6'h1 == T_28597 ? T_38110_1_pdst : T_38110_0_pdst; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24596 = 6'h1 == T_28597 ? T_38110_1_ldst_val : T_38110_0_ldst_val; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24650 = 6'h2 == T_28597 ? T_38110_2_pdst : _GEN_24572; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24674 = 6'h2 == T_28597 ? T_38110_2_ldst_val : _GEN_24596; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24728 = 6'h3 == T_28597 ? T_38110_3_pdst : _GEN_24650; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24752 = 6'h3 == T_28597 ? T_38110_3_ldst_val : _GEN_24674; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24806 = 6'h4 == T_28597 ? T_38110_4_pdst : _GEN_24728; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24830 = 6'h4 == T_28597 ? T_38110_4_ldst_val : _GEN_24752; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24884 = 6'h5 == T_28597 ? T_38110_5_pdst : _GEN_24806; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24908 = 6'h5 == T_28597 ? T_38110_5_ldst_val : _GEN_24830; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_24962 = 6'h6 == T_28597 ? T_38110_6_pdst : _GEN_24884; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_24986 = 6'h6 == T_28597 ? T_38110_6_ldst_val : _GEN_24908; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25040 = 6'h7 == T_28597 ? T_38110_7_pdst : _GEN_24962; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25064 = 6'h7 == T_28597 ? T_38110_7_ldst_val : _GEN_24986; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25118 = 6'h8 == T_28597 ? T_38110_8_pdst : _GEN_25040; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25142 = 6'h8 == T_28597 ? T_38110_8_ldst_val : _GEN_25064; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25196 = 6'h9 == T_28597 ? T_38110_9_pdst : _GEN_25118; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25220 = 6'h9 == T_28597 ? T_38110_9_ldst_val : _GEN_25142; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25274 = 6'ha == T_28597 ? T_38110_10_pdst : _GEN_25196; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25298 = 6'ha == T_28597 ? T_38110_10_ldst_val : _GEN_25220; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25352 = 6'hb == T_28597 ? T_38110_11_pdst : _GEN_25274; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25376 = 6'hb == T_28597 ? T_38110_11_ldst_val : _GEN_25298; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25430 = 6'hc == T_28597 ? T_38110_12_pdst : _GEN_25352; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25454 = 6'hc == T_28597 ? T_38110_12_ldst_val : _GEN_25376; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25508 = 6'hd == T_28597 ? T_38110_13_pdst : _GEN_25430; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25532 = 6'hd == T_28597 ? T_38110_13_ldst_val : _GEN_25454; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25586 = 6'he == T_28597 ? T_38110_14_pdst : _GEN_25508; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25610 = 6'he == T_28597 ? T_38110_14_ldst_val : _GEN_25532; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25664 = 6'hf == T_28597 ? T_38110_15_pdst : _GEN_25586; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25688 = 6'hf == T_28597 ? T_38110_15_ldst_val : _GEN_25610; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25742 = 6'h10 == T_28597 ? T_38110_16_pdst : _GEN_25664; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25766 = 6'h10 == T_28597 ? T_38110_16_ldst_val : _GEN_25688; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25820 = 6'h11 == T_28597 ? T_38110_17_pdst : _GEN_25742; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25844 = 6'h11 == T_28597 ? T_38110_17_ldst_val : _GEN_25766; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25898 = 6'h12 == T_28597 ? T_38110_18_pdst : _GEN_25820; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_25922 = 6'h12 == T_28597 ? T_38110_18_ldst_val : _GEN_25844; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_25976 = 6'h13 == T_28597 ? T_38110_19_pdst : _GEN_25898; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26000 = 6'h13 == T_28597 ? T_38110_19_ldst_val : _GEN_25922; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26054 = 6'h14 == T_28597 ? T_38110_20_pdst : _GEN_25976; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26078 = 6'h14 == T_28597 ? T_38110_20_ldst_val : _GEN_26000; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26132 = 6'h15 == T_28597 ? T_38110_21_pdst : _GEN_26054; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26156 = 6'h15 == T_28597 ? T_38110_21_ldst_val : _GEN_26078; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26210 = 6'h16 == T_28597 ? T_38110_22_pdst : _GEN_26132; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26234 = 6'h16 == T_28597 ? T_38110_22_ldst_val : _GEN_26156; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26288 = 6'h17 == T_28597 ? T_38110_23_pdst : _GEN_26210; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26312 = 6'h17 == T_28597 ? T_38110_23_ldst_val : _GEN_26234; // @[rob.scala 538:75 rob.scala 538:75]
  wire  T_44496 = T_40529 & _GEN_26312; // @[rob.scala 538:75]
  wire  T_44497 = _GEN_26288 != io_wb_resps_1_bits_uop_pdst; // @[rob.scala 539:54]
  wire  T_44498 = T_44496 & T_44497; // @[rob.scala 539:37]
  wire  T_44500 = ~T_44498; // @[rob.scala 538:18]
  wire  T_44501 = T_44500 | reset; // @[rob.scala 538:17]
  wire  T_44503 = ~T_44501; // @[rob.scala 538:17]
  wire  T_44507 = io_debug_wb_valids_2 & T_28606; // @[rob.scala 529:38]
  wire  _GEN_26372 = 6'h1 == T_28605 ? T_35634_1 : T_35634_0; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26373 = 6'h2 == T_28605 ? T_35634_2 : _GEN_26372; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26374 = 6'h3 == T_28605 ? T_35634_3 : _GEN_26373; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26375 = 6'h4 == T_28605 ? T_35634_4 : _GEN_26374; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26376 = 6'h5 == T_28605 ? T_35634_5 : _GEN_26375; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26377 = 6'h6 == T_28605 ? T_35634_6 : _GEN_26376; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26378 = 6'h7 == T_28605 ? T_35634_7 : _GEN_26377; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26379 = 6'h8 == T_28605 ? T_35634_8 : _GEN_26378; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26380 = 6'h9 == T_28605 ? T_35634_9 : _GEN_26379; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26381 = 6'ha == T_28605 ? T_35634_10 : _GEN_26380; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26382 = 6'hb == T_28605 ? T_35634_11 : _GEN_26381; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26383 = 6'hc == T_28605 ? T_35634_12 : _GEN_26382; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26384 = 6'hd == T_28605 ? T_35634_13 : _GEN_26383; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26385 = 6'he == T_28605 ? T_35634_14 : _GEN_26384; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26386 = 6'hf == T_28605 ? T_35634_15 : _GEN_26385; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26387 = 6'h10 == T_28605 ? T_35634_16 : _GEN_26386; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26388 = 6'h11 == T_28605 ? T_35634_17 : _GEN_26387; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26389 = 6'h12 == T_28605 ? T_35634_18 : _GEN_26388; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26390 = 6'h13 == T_28605 ? T_35634_19 : _GEN_26389; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26391 = 6'h14 == T_28605 ? T_35634_20 : _GEN_26390; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26392 = 6'h15 == T_28605 ? T_35634_21 : _GEN_26391; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26393 = 6'h16 == T_28605 ? T_35634_22 : _GEN_26392; // @[rob.scala 536:22 rob.scala 536:22]
  wire  _GEN_26394 = 6'h17 == T_28605 ? T_35634_23 : _GEN_26393; // @[rob.scala 536:22 rob.scala 536:22]
  wire  T_44689 = ~_GEN_26394; // @[rob.scala 536:22]
  wire  T_44690 = T_40537 & T_44689; // @[rob.scala 535:75]
  wire  T_44692 = ~T_44690; // @[rob.scala 535:18]
  wire  T_44693 = T_44692 | reset; // @[rob.scala 535:17]
  wire  T_44695 = ~T_44693; // @[rob.scala 535:17]
  wire [6:0] _GEN_26516 = 6'h1 == T_28605 ? T_38110_1_pdst : T_38110_0_pdst; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26540 = 6'h1 == T_28605 ? T_38110_1_ldst_val : T_38110_0_ldst_val; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26594 = 6'h2 == T_28605 ? T_38110_2_pdst : _GEN_26516; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26618 = 6'h2 == T_28605 ? T_38110_2_ldst_val : _GEN_26540; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26672 = 6'h3 == T_28605 ? T_38110_3_pdst : _GEN_26594; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26696 = 6'h3 == T_28605 ? T_38110_3_ldst_val : _GEN_26618; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26750 = 6'h4 == T_28605 ? T_38110_4_pdst : _GEN_26672; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26774 = 6'h4 == T_28605 ? T_38110_4_ldst_val : _GEN_26696; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26828 = 6'h5 == T_28605 ? T_38110_5_pdst : _GEN_26750; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26852 = 6'h5 == T_28605 ? T_38110_5_ldst_val : _GEN_26774; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26906 = 6'h6 == T_28605 ? T_38110_6_pdst : _GEN_26828; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_26930 = 6'h6 == T_28605 ? T_38110_6_ldst_val : _GEN_26852; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_26984 = 6'h7 == T_28605 ? T_38110_7_pdst : _GEN_26906; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27008 = 6'h7 == T_28605 ? T_38110_7_ldst_val : _GEN_26930; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27062 = 6'h8 == T_28605 ? T_38110_8_pdst : _GEN_26984; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27086 = 6'h8 == T_28605 ? T_38110_8_ldst_val : _GEN_27008; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27140 = 6'h9 == T_28605 ? T_38110_9_pdst : _GEN_27062; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27164 = 6'h9 == T_28605 ? T_38110_9_ldst_val : _GEN_27086; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27218 = 6'ha == T_28605 ? T_38110_10_pdst : _GEN_27140; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27242 = 6'ha == T_28605 ? T_38110_10_ldst_val : _GEN_27164; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27296 = 6'hb == T_28605 ? T_38110_11_pdst : _GEN_27218; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27320 = 6'hb == T_28605 ? T_38110_11_ldst_val : _GEN_27242; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27374 = 6'hc == T_28605 ? T_38110_12_pdst : _GEN_27296; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27398 = 6'hc == T_28605 ? T_38110_12_ldst_val : _GEN_27320; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27452 = 6'hd == T_28605 ? T_38110_13_pdst : _GEN_27374; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27476 = 6'hd == T_28605 ? T_38110_13_ldst_val : _GEN_27398; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27530 = 6'he == T_28605 ? T_38110_14_pdst : _GEN_27452; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27554 = 6'he == T_28605 ? T_38110_14_ldst_val : _GEN_27476; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27608 = 6'hf == T_28605 ? T_38110_15_pdst : _GEN_27530; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27632 = 6'hf == T_28605 ? T_38110_15_ldst_val : _GEN_27554; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27686 = 6'h10 == T_28605 ? T_38110_16_pdst : _GEN_27608; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27710 = 6'h10 == T_28605 ? T_38110_16_ldst_val : _GEN_27632; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27764 = 6'h11 == T_28605 ? T_38110_17_pdst : _GEN_27686; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27788 = 6'h11 == T_28605 ? T_38110_17_ldst_val : _GEN_27710; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27842 = 6'h12 == T_28605 ? T_38110_18_pdst : _GEN_27764; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27866 = 6'h12 == T_28605 ? T_38110_18_ldst_val : _GEN_27788; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27920 = 6'h13 == T_28605 ? T_38110_19_pdst : _GEN_27842; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_27944 = 6'h13 == T_28605 ? T_38110_19_ldst_val : _GEN_27866; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_27998 = 6'h14 == T_28605 ? T_38110_20_pdst : _GEN_27920; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_28022 = 6'h14 == T_28605 ? T_38110_20_ldst_val : _GEN_27944; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_28076 = 6'h15 == T_28605 ? T_38110_21_pdst : _GEN_27998; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_28100 = 6'h15 == T_28605 ? T_38110_21_ldst_val : _GEN_28022; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_28154 = 6'h16 == T_28605 ? T_38110_22_pdst : _GEN_28076; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_28178 = 6'h16 == T_28605 ? T_38110_22_ldst_val : _GEN_28100; // @[rob.scala 538:75 rob.scala 538:75]
  wire [6:0] _GEN_28232 = 6'h17 == T_28605 ? T_38110_23_pdst : _GEN_28154; // @[rob.scala 538:75 rob.scala 538:75]
  wire  _GEN_28256 = 6'h17 == T_28605 ? T_38110_23_ldst_val : _GEN_28178; // @[rob.scala 538:75 rob.scala 538:75]
  wire  T_44700 = T_40537 & _GEN_28256; // @[rob.scala 538:75]
  wire  T_44701 = _GEN_28232 != io_wb_resps_2_bits_uop_pdst; // @[rob.scala 539:54]
  wire  T_44702 = T_44700 & T_44701; // @[rob.scala 539:37]
  wire  T_44704 = ~T_44702; // @[rob.scala 538:18]
  wire  T_44705 = T_44704 | reset; // @[rob.scala 538:17]
  wire  T_44707 = ~T_44705; // @[rob.scala 538:17]
  wire [39:0] T_44888 = {T_23555_T_44886_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_44883 = {{24'd0}, T_44888}; // @[rob.scala 899:26]
  wire [39:0] T_44895 = T_44883[39:0]; // @[rob.scala 906:20]
  wire  T_44896 = T_44895[39]; // @[util.scala 114:43]
  wire [23:0] T_44900 = T_44896 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_44901 = {T_44900,T_44895}; // @[Cat.scala 20:58]
  wire [63:0] T_44904 = T_44901 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45008 = {T_23558_T_45006_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_44997 = {{24'd0}, T_45008}; // @[rob.scala 899:26]
  wire [39:0] T_45009 = T_44997[39:0]; // @[rob.scala 906:20]
  wire  T_45010 = T_45009[39]; // @[util.scala 114:43]
  wire [23:0] T_45014 = T_45010 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45015 = {T_45014,T_45009}; // @[Cat.scala 20:58]
  wire [63:0] T_45018 = T_45015 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45116 = {T_23555_T_45114_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_45111 = {{24'd0}, T_45116}; // @[rob.scala 899:26]
  wire [39:0] T_45123 = T_45111[39:0]; // @[rob.scala 906:20]
  wire  T_45124 = T_45123[39]; // @[util.scala 114:43]
  wire [23:0] T_45128 = T_45124 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45129 = {T_45128,T_45123}; // @[Cat.scala 20:58]
  wire [63:0] T_45132 = T_45129 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45236 = {T_23558_T_45234_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_45225 = {{24'd0}, T_45236}; // @[rob.scala 899:26]
  wire [39:0] T_45237 = T_45225[39:0]; // @[rob.scala 906:20]
  wire  T_45238 = T_45237[39]; // @[util.scala 114:43]
  wire [23:0] T_45242 = T_45238 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45243 = {T_45242,T_45237}; // @[Cat.scala 20:58]
  wire [63:0] T_45246 = T_45243 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45344 = {T_23555_T_45342_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_45339 = {{24'd0}, T_45344}; // @[rob.scala 899:26]
  wire [39:0] T_45351 = T_45339[39:0]; // @[rob.scala 906:20]
  wire  T_45352 = T_45351[39]; // @[util.scala 114:43]
  wire [23:0] T_45356 = T_45352 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45357 = {T_45356,T_45351}; // @[Cat.scala 20:58]
  wire [63:0] T_45360 = T_45357 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45464 = {T_23558_T_45462_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_45453 = {{24'd0}, T_45464}; // @[rob.scala 899:26]
  wire [39:0] T_45465 = T_45453[39:0]; // @[rob.scala 906:20]
  wire  T_45466 = T_45465[39]; // @[util.scala 114:43]
  wire [23:0] T_45470 = T_45466 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45471 = {T_45470,T_45465}; // @[Cat.scala 20:58]
  wire [63:0] T_45474 = T_45471 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45572 = {T_23555_T_45570_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_45567 = {{24'd0}, T_45572}; // @[rob.scala 899:26]
  wire [39:0] T_45579 = T_45567[39:0]; // @[rob.scala 906:20]
  wire  T_45580 = T_45579[39]; // @[util.scala 114:43]
  wire [23:0] T_45584 = T_45580 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45585 = {T_45584,T_45579}; // @[Cat.scala 20:58]
  wire [63:0] T_45588 = T_45585 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45692 = {T_23558_T_45690_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_45681 = {{24'd0}, T_45692}; // @[rob.scala 899:26]
  wire [39:0] T_45693 = T_45681[39:0]; // @[rob.scala 906:20]
  wire  T_45694 = T_45693[39]; // @[util.scala 114:43]
  wire [23:0] T_45698 = T_45694 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45699 = {T_45698,T_45693}; // @[Cat.scala 20:58]
  wire [63:0] T_45702 = T_45699 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45800 = {T_23555_T_45798_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_45795 = {{24'd0}, T_45800}; // @[rob.scala 899:26]
  wire [39:0] T_45807 = T_45795[39:0]; // @[rob.scala 906:20]
  wire  T_45808 = T_45807[39]; // @[util.scala 114:43]
  wire [23:0] T_45812 = T_45808 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45813 = {T_45812,T_45807}; // @[Cat.scala 20:58]
  wire [63:0] T_45816 = T_45813 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_45920 = {T_23558_T_45918_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_45909 = {{24'd0}, T_45920}; // @[rob.scala 899:26]
  wire [39:0] T_45921 = T_45909[39:0]; // @[rob.scala 906:20]
  wire  T_45922 = T_45921[39]; // @[util.scala 114:43]
  wire [23:0] T_45926 = T_45922 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_45927 = {T_45926,T_45921}; // @[Cat.scala 20:58]
  wire [63:0] T_45930 = T_45927 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46028 = {T_23555_T_46026_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_46023 = {{24'd0}, T_46028}; // @[rob.scala 899:26]
  wire [39:0] T_46035 = T_46023[39:0]; // @[rob.scala 906:20]
  wire  T_46036 = T_46035[39]; // @[util.scala 114:43]
  wire [23:0] T_46040 = T_46036 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46041 = {T_46040,T_46035}; // @[Cat.scala 20:58]
  wire [63:0] T_46044 = T_46041 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46148 = {T_23558_T_46146_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_46137 = {{24'd0}, T_46148}; // @[rob.scala 899:26]
  wire [39:0] T_46149 = T_46137[39:0]; // @[rob.scala 906:20]
  wire  T_46150 = T_46149[39]; // @[util.scala 114:43]
  wire [23:0] T_46154 = T_46150 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46155 = {T_46154,T_46149}; // @[Cat.scala 20:58]
  wire [63:0] T_46158 = T_46155 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46256 = {T_23555_T_46254_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_46251 = {{24'd0}, T_46256}; // @[rob.scala 899:26]
  wire [39:0] T_46263 = T_46251[39:0]; // @[rob.scala 906:20]
  wire  T_46264 = T_46263[39]; // @[util.scala 114:43]
  wire [23:0] T_46268 = T_46264 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46269 = {T_46268,T_46263}; // @[Cat.scala 20:58]
  wire [63:0] T_46272 = T_46269 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46376 = {T_23558_T_46374_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_46365 = {{24'd0}, T_46376}; // @[rob.scala 899:26]
  wire [39:0] T_46377 = T_46365[39:0]; // @[rob.scala 906:20]
  wire  T_46378 = T_46377[39]; // @[util.scala 114:43]
  wire [23:0] T_46382 = T_46378 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46383 = {T_46382,T_46377}; // @[Cat.scala 20:58]
  wire [63:0] T_46386 = T_46383 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46484 = {T_23555_T_46482_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_46479 = {{24'd0}, T_46484}; // @[rob.scala 899:26]
  wire [39:0] T_46491 = T_46479[39:0]; // @[rob.scala 906:20]
  wire  T_46492 = T_46491[39]; // @[util.scala 114:43]
  wire [23:0] T_46496 = T_46492 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46497 = {T_46496,T_46491}; // @[Cat.scala 20:58]
  wire [63:0] T_46500 = T_46497 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46604 = {T_23558_T_46602_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_46593 = {{24'd0}, T_46604}; // @[rob.scala 899:26]
  wire [39:0] T_46605 = T_46593[39:0]; // @[rob.scala 906:20]
  wire  T_46606 = T_46605[39]; // @[util.scala 114:43]
  wire [23:0] T_46610 = T_46606 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46611 = {T_46610,T_46605}; // @[Cat.scala 20:58]
  wire [63:0] T_46614 = T_46611 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46712 = {T_23555_T_46710_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_46707 = {{24'd0}, T_46712}; // @[rob.scala 899:26]
  wire [39:0] T_46719 = T_46707[39:0]; // @[rob.scala 906:20]
  wire  T_46720 = T_46719[39]; // @[util.scala 114:43]
  wire [23:0] T_46724 = T_46720 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46725 = {T_46724,T_46719}; // @[Cat.scala 20:58]
  wire [63:0] T_46728 = T_46725 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46832 = {T_23558_T_46830_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_46821 = {{24'd0}, T_46832}; // @[rob.scala 899:26]
  wire [39:0] T_46833 = T_46821[39:0]; // @[rob.scala 906:20]
  wire  T_46834 = T_46833[39]; // @[util.scala 114:43]
  wire [23:0] T_46838 = T_46834 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46839 = {T_46838,T_46833}; // @[Cat.scala 20:58]
  wire [63:0] T_46842 = T_46839 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_46940 = {T_23555_T_46938_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_46935 = {{24'd0}, T_46940}; // @[rob.scala 899:26]
  wire [39:0] T_46947 = T_46935[39:0]; // @[rob.scala 906:20]
  wire  T_46948 = T_46947[39]; // @[util.scala 114:43]
  wire [23:0] T_46952 = T_46948 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_46953 = {T_46952,T_46947}; // @[Cat.scala 20:58]
  wire [63:0] T_46956 = T_46953 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_47060 = {T_23558_T_47058_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_47049 = {{24'd0}, T_47060}; // @[rob.scala 899:26]
  wire [39:0] T_47061 = T_47049[39:0]; // @[rob.scala 906:20]
  wire  T_47062 = T_47061[39]; // @[util.scala 114:43]
  wire [23:0] T_47066 = T_47062 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_47067 = {T_47066,T_47061}; // @[Cat.scala 20:58]
  wire [63:0] T_47070 = T_47067 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_47168 = {T_23555_T_47166_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_47163 = {{24'd0}, T_47168}; // @[rob.scala 899:26]
  wire [39:0] T_47175 = T_47163[39:0]; // @[rob.scala 906:20]
  wire  T_47176 = T_47175[39]; // @[util.scala 114:43]
  wire [23:0] T_47180 = T_47176 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_47181 = {T_47180,T_47175}; // @[Cat.scala 20:58]
  wire [63:0] T_47184 = T_47181 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_47288 = {T_23558_T_47286_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_47277 = {{24'd0}, T_47288}; // @[rob.scala 899:26]
  wire [39:0] T_47289 = T_47277[39:0]; // @[rob.scala 906:20]
  wire  T_47290 = T_47289[39]; // @[util.scala 114:43]
  wire [23:0] T_47294 = T_47290 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_47295 = {T_47294,T_47289}; // @[Cat.scala 20:58]
  wire [63:0] T_47298 = T_47295 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_47396 = {T_23555_T_47394_data, 3'h0}; // @[rob.scala 900:45]
  wire [63:0] T_47391 = {{24'd0}, T_47396}; // @[rob.scala 899:26]
  wire [39:0] T_47403 = T_47391[39:0]; // @[rob.scala 906:20]
  wire  T_47404 = T_47403[39]; // @[util.scala 114:43]
  wire [23:0] T_47408 = T_47404 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_47409 = {T_47408,T_47403}; // @[Cat.scala 20:58]
  wire [63:0] T_47412 = T_47409 + 64'h4; // @[rob.scala 554:94]
  wire [39:0] T_47516 = {T_23558_T_47514_data, 3'h0}; // @[rob.scala 904:48]
  wire [63:0] T_47505 = {{24'd0}, T_47516}; // @[rob.scala 899:26]
  wire [39:0] T_47517 = T_47505[39:0]; // @[rob.scala 906:20]
  wire  T_47518 = T_47517[39]; // @[util.scala 114:43]
  wire [23:0] T_47522 = T_47518 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_47523 = {T_47522,T_47517}; // @[Cat.scala 20:58]
  wire [63:0] T_47526 = T_47523 + 64'h4; // @[rob.scala 554:94]
  wire  T_47536 = T_29090 & T_47545; // @[rob.scala 583:54]
  wire  T_47554 = T_41018 & T_47562; // @[rob.scala 583:54]
  wire  T_47557 = T_47554 & T_32081; // @[rob.scala 583:71]
  wire  will_throw_exception = T_47557 | T_47536; // @[rob.scala 583:87]
  wire  T_47568 = will_throw_exception | io_cxcpt_valid; // @[rob.scala 593:48]
  wire  T_47569 = io_com_exc_cause == 64'hd; // @[rob.scala 594:45]
  wire  T_47570 = io_com_exc_cause == 64'he; // @[rob.scala 595:45]
  wire  is_mini_exception = T_47569 | T_47570; // @[rob.scala 594:77]
  wire  T_47572 = ~is_mini_exception; // @[rob.scala 596:47]
  reg  T_47576;
  wire  T_47577 = r_xcpt_badvaddr[39]; // @[util.scala 114:43]
  wire [23:0] T_47581 = T_47577 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [4:0] T_47586 = {{1'd0}, rob_head[4:1]}; // @[rob.scala 900:33]
  wire [39:0] T_47589 = {T_23555_T_47587_data, 3'h0}; // @[rob.scala 900:45]
  wire  T_47590 = rob_head[0]; // @[rob.scala 902:23]
  wire [39:0] T_47595 = {T_23558_T_47593_data, 3'h0}; // @[rob.scala 904:48]
  wire [39:0] _GEN_28318 = T_47590 ? T_47595 : T_47589; // @[rob.scala 903:10 rob.scala 904:19 rob.scala 900:16]
  wire [63:0] T_47584 = {{24'd0}, _GEN_28318}; // @[rob.scala 899:26]
  wire [39:0] T_47596 = T_47584[39:0]; // @[rob.scala 906:20]
  wire  T_47597 = T_47596[39]; // @[util.scala 114:43]
  wire [23:0] T_47601 = T_47597 ? 24'hffffff : 24'h0; // @[Bitwise.scala 33:12]
  wire [63:0] T_47602 = {T_47601,T_47596}; // @[Cat.scala 20:58]
  wire [2:0] T_47605 = rob_head_vals_0 ? 3'h0 : 3'h4; // @[Mux.scala 31:69]
  wire [63:0] _GEN_28920 = {{61'd0}, T_47605}; // @[rob.scala 605:46]
  wire [63:0] T_47607 = T_47602 + _GEN_28920; // @[rob.scala 605:46]
  wire [2:0] T_47610 = T_47568 ? 3'h0 : 3'h4; // @[rob.scala 607:23]
  wire [63:0] _GEN_28921 = {{61'd0}, T_47610}; // @[rob.scala 606:86]
  wire [63:0] T_47612 = T_47607 + _GEN_28921; // @[rob.scala 606:86]
  wire  T_47613 = io_com_valids_0 & io_com_uops_0_flush_on_commit; // @[rob.scala 609:64]
  wire  T_47614 = io_com_valids_1 & io_com_uops_1_flush_on_commit; // @[rob.scala 609:64]
  wire  T_47615 = T_47613 | T_47614; // @[rob.scala 609:108]
  reg  T_47616;
  wire  T_47631 = io_com_valids_0 & io_com_uops_0_fp_val; // @[rob.scala 624:41]
  wire  T_47632 = io_com_uops_0_is_load | io_com_uops_0_is_store; // @[rob.scala 626:48]
  wire  T_47634 = ~T_47632; // @[rob.scala 626:23]
  wire  T_47635 = T_47631 & T_47634; // @[rob.scala 625:46]
  wire [4:0] rob_head_fflags_0 = T_28314_T_31814_data; // @[rob.scala 201:34 rob.scala 506:28]
  wire [4:0] T_47637 = T_47635 ? rob_head_fflags_0 : 5'h0; // @[rob.scala 628:23]
  wire  T_47639 = ~io_com_uops_0_fp_val; // @[rob.scala 631:16]
  wire  T_47640 = io_com_valids_0 & T_47639; // @[rob.scala 630:34]
  wire  T_47642 = rob_head_fflags_0 != 5'h0; // @[rob.scala 632:35]
  wire  T_47643 = T_47640 & T_47642; // @[rob.scala 631:39]
  wire  T_47645 = ~T_47643; // @[rob.scala 630:15]
  wire  T_47646 = T_47645 | reset; // @[rob.scala 630:14]
  wire  T_47648 = ~T_47646; // @[rob.scala 630:14]
  wire  T_47651 = T_47631 & T_47632; // @[rob.scala 635:38]
  wire  T_47654 = T_47651 & T_47642; // @[rob.scala 636:68]
  wire  T_47656 = ~T_47654; // @[rob.scala 634:15]
  wire  T_47657 = T_47656 | reset; // @[rob.scala 634:14]
  wire  T_47659 = ~T_47657; // @[rob.scala 634:14]
  wire  T_47660 = io_com_valids_1 & io_com_uops_1_fp_val; // @[rob.scala 624:41]
  wire  T_47661 = io_com_uops_1_is_load | io_com_uops_1_is_store; // @[rob.scala 626:48]
  wire  T_47663 = ~T_47661; // @[rob.scala 626:23]
  wire  T_47664 = T_47660 & T_47663; // @[rob.scala 625:46]
  wire [4:0] rob_head_fflags_1 = T_40242_T_43742_data; // @[rob.scala 201:34 rob.scala 506:28]
  wire [4:0] T_47666 = T_47664 ? rob_head_fflags_1 : 5'h0; // @[rob.scala 628:23]
  wire  T_47668 = ~io_com_uops_1_fp_val; // @[rob.scala 631:16]
  wire  T_47669 = io_com_valids_1 & T_47668; // @[rob.scala 630:34]
  wire  T_47671 = rob_head_fflags_1 != 5'h0; // @[rob.scala 632:35]
  wire  T_47672 = T_47669 & T_47671; // @[rob.scala 631:39]
  wire  T_47674 = ~T_47672; // @[rob.scala 630:15]
  wire  T_47675 = T_47674 | reset; // @[rob.scala 630:14]
  wire  T_47677 = ~T_47675; // @[rob.scala 630:14]
  wire  T_47680 = T_47660 & T_47661; // @[rob.scala 635:38]
  wire  T_47683 = T_47680 & T_47671; // @[rob.scala 636:68]
  wire  T_47685 = ~T_47683; // @[rob.scala 634:15]
  wire  T_47686 = T_47685 | reset; // @[rob.scala 634:14]
  wire  T_47688 = ~T_47686; // @[rob.scala 634:14]
  wire  T_47869 = io_dis_valids_0 & io_dis_uops_0_exception; // @[rob.scala 656:40]
  wire  T_47870 = io_dis_valids_1 & io_dis_uops_1_exception; // @[rob.scala 656:40]
  wire  T_47871 = io_flush_pipeline | T_47568; // @[rob.scala 659:30]
  wire  T_47873 = ~T_47871; // @[rob.scala 659:10]
  wire  T_47874 = rob_state != 2'h2; // @[rob.scala 659:64]
  wire  T_47875 = T_47873 & T_47874; // @[rob.scala 659:51]
  wire  T_47876 = io_lxcpt_valid | io_bxcpt_valid; // @[rob.scala 661:28]
  wire  T_47878 = ~io_bxcpt_valid; // @[rob.scala 663:49]
  wire  T_47879 = io_lxcpt_valid & T_47878; // @[rob.scala 663:46]
  wire  T_47880 = io_lxcpt_valid & io_bxcpt_valid; // @[rob.scala 664:46]
  wire  T_47881 = io_lxcpt_bits_uop_rob_idx <= rob_tail_idx; // @[rob.scala 650:58]
  wire [6:0] T_47882 = {T_47881,io_lxcpt_bits_uop_rob_idx}; // @[Cat.scala 20:58]
  wire  T_47883 = io_bxcpt_bits_uop_rob_idx <= rob_tail_idx; // @[rob.scala 650:80]
  wire [6:0] T_47884 = {T_47883,io_bxcpt_bits_uop_rob_idx}; // @[Cat.scala 20:58]
  wire  T_47885 = T_47882 < T_47884; // @[rob.scala 650:71]
  wire  T_47886 = T_47880 & T_47885; // @[rob.scala 664:64]
  wire  T_47887 = T_47879 | T_47886; // @[rob.scala 663:66]
  wire  T_47888_valid = T_47887 ? io_lxcpt_bits_uop_valid : io_bxcpt_bits_uop_valid; // @[rob.scala 666:32]
  wire [1:0] T_47888_iw_state = T_47887 ? io_lxcpt_bits_uop_iw_state : io_bxcpt_bits_uop_iw_state; // @[rob.scala 666:32]
  wire [8:0] T_47888_uopc = T_47887 ? io_lxcpt_bits_uop_uopc : io_bxcpt_bits_uop_uopc; // @[rob.scala 666:32]
  wire [31:0] T_47888_inst = T_47887 ? io_lxcpt_bits_uop_inst : io_bxcpt_bits_uop_inst; // @[rob.scala 666:32]
  wire [39:0] T_47888_pc = T_47887 ? io_lxcpt_bits_uop_pc : io_bxcpt_bits_uop_pc; // @[rob.scala 666:32]
  wire [7:0] T_47888_fu_code = T_47887 ? io_lxcpt_bits_uop_fu_code : io_bxcpt_bits_uop_fu_code; // @[rob.scala 666:32]
  wire [3:0] T_47888_ctrl_br_type = T_47887 ? io_lxcpt_bits_uop_ctrl_br_type : io_bxcpt_bits_uop_ctrl_br_type; // @[rob.scala 666:32]
  wire [1:0] T_47888_ctrl_op1_sel = T_47887 ? io_lxcpt_bits_uop_ctrl_op1_sel : io_bxcpt_bits_uop_ctrl_op1_sel; // @[rob.scala 666:32]
  wire [2:0] T_47888_ctrl_op2_sel = T_47887 ? io_lxcpt_bits_uop_ctrl_op2_sel : io_bxcpt_bits_uop_ctrl_op2_sel; // @[rob.scala 666:32]
  wire [2:0] T_47888_ctrl_imm_sel = T_47887 ? io_lxcpt_bits_uop_ctrl_imm_sel : io_bxcpt_bits_uop_ctrl_imm_sel; // @[rob.scala 666:32]
  wire [3:0] T_47888_ctrl_op_fcn = T_47887 ? io_lxcpt_bits_uop_ctrl_op_fcn : io_bxcpt_bits_uop_ctrl_op_fcn; // @[rob.scala 666:32]
  wire  T_47888_ctrl_fcn_dw = T_47887 ? io_lxcpt_bits_uop_ctrl_fcn_dw : io_bxcpt_bits_uop_ctrl_fcn_dw; // @[rob.scala 666:32]
  wire  T_47888_ctrl_rf_wen = T_47887 ? io_lxcpt_bits_uop_ctrl_rf_wen : io_bxcpt_bits_uop_ctrl_rf_wen; // @[rob.scala 666:32]
  wire [2:0] T_47888_ctrl_csr_cmd = T_47887 ? io_lxcpt_bits_uop_ctrl_csr_cmd : io_bxcpt_bits_uop_ctrl_csr_cmd; // @[rob.scala 666:32]
  wire  T_47888_ctrl_is_load = T_47887 ? io_lxcpt_bits_uop_ctrl_is_load : io_bxcpt_bits_uop_ctrl_is_load; // @[rob.scala 666:32]
  wire  T_47888_ctrl_is_sta = T_47887 ? io_lxcpt_bits_uop_ctrl_is_sta : io_bxcpt_bits_uop_ctrl_is_sta; // @[rob.scala 666:32]
  wire  T_47888_ctrl_is_std = T_47887 ? io_lxcpt_bits_uop_ctrl_is_std : io_bxcpt_bits_uop_ctrl_is_std; // @[rob.scala 666:32]
  wire [1:0] T_47888_wakeup_delay = T_47887 ? io_lxcpt_bits_uop_wakeup_delay : io_bxcpt_bits_uop_wakeup_delay; // @[rob.scala 666:32]
  wire  T_47888_allocate_brtag = T_47887 ? io_lxcpt_bits_uop_allocate_brtag : io_bxcpt_bits_uop_allocate_brtag; // @[rob.scala 666:32]
  wire  T_47888_is_br_or_jmp = T_47887 ? io_lxcpt_bits_uop_is_br_or_jmp : io_bxcpt_bits_uop_is_br_or_jmp; // @[rob.scala 666:32]
  wire  T_47888_is_jump = T_47887 ? io_lxcpt_bits_uop_is_jump : io_bxcpt_bits_uop_is_jump; // @[rob.scala 666:32]
  wire  T_47888_is_jal = T_47887 ? io_lxcpt_bits_uop_is_jal : io_bxcpt_bits_uop_is_jal; // @[rob.scala 666:32]
  wire  T_47888_is_ret = T_47887 ? io_lxcpt_bits_uop_is_ret : io_bxcpt_bits_uop_is_ret; // @[rob.scala 666:32]
  wire  T_47888_is_call = T_47887 ? io_lxcpt_bits_uop_is_call : io_bxcpt_bits_uop_is_call; // @[rob.scala 666:32]
  wire [7:0] T_47888_br_mask = T_47887 ? io_lxcpt_bits_uop_br_mask : io_bxcpt_bits_uop_br_mask; // @[rob.scala 666:32]
  wire [2:0] T_47888_br_tag = T_47887 ? io_lxcpt_bits_uop_br_tag : io_bxcpt_bits_uop_br_tag; // @[rob.scala 666:32]
  wire  T_47888_br_prediction_bpd_predict_val = T_47887 ? io_lxcpt_bits_uop_br_prediction_bpd_predict_val :
    io_bxcpt_bits_uop_br_prediction_bpd_predict_val; // @[rob.scala 666:32]
  wire  T_47888_br_prediction_bpd_predict_taken = T_47887 ? io_lxcpt_bits_uop_br_prediction_bpd_predict_taken :
    io_bxcpt_bits_uop_br_prediction_bpd_predict_taken; // @[rob.scala 666:32]
  wire  T_47888_br_prediction_btb_hit = T_47887 ? io_lxcpt_bits_uop_br_prediction_btb_hit :
    io_bxcpt_bits_uop_br_prediction_btb_hit; // @[rob.scala 666:32]
  wire  T_47888_br_prediction_btb_predicted = T_47887 ? io_lxcpt_bits_uop_br_prediction_btb_predicted :
    io_bxcpt_bits_uop_br_prediction_btb_predicted; // @[rob.scala 666:32]
  wire  T_47888_br_prediction_is_br_or_jalr = T_47887 ? io_lxcpt_bits_uop_br_prediction_is_br_or_jalr :
    io_bxcpt_bits_uop_br_prediction_is_br_or_jalr; // @[rob.scala 666:32]
  wire  T_47888_stat_brjmp_mispredicted = T_47887 ? io_lxcpt_bits_uop_stat_brjmp_mispredicted :
    io_bxcpt_bits_uop_stat_brjmp_mispredicted; // @[rob.scala 666:32]
  wire  T_47888_stat_btb_made_pred = T_47887 ? io_lxcpt_bits_uop_stat_btb_made_pred :
    io_bxcpt_bits_uop_stat_btb_made_pred; // @[rob.scala 666:32]
  wire  T_47888_stat_btb_mispredicted = T_47887 ? io_lxcpt_bits_uop_stat_btb_mispredicted :
    io_bxcpt_bits_uop_stat_btb_mispredicted; // @[rob.scala 666:32]
  wire  T_47888_stat_bpd_made_pred = T_47887 ? io_lxcpt_bits_uop_stat_bpd_made_pred :
    io_bxcpt_bits_uop_stat_bpd_made_pred; // @[rob.scala 666:32]
  wire  T_47888_stat_bpd_mispredicted = T_47887 ? io_lxcpt_bits_uop_stat_bpd_mispredicted :
    io_bxcpt_bits_uop_stat_bpd_mispredicted; // @[rob.scala 666:32]
  wire [2:0] T_47888_fetch_pc_lob = T_47887 ? io_lxcpt_bits_uop_fetch_pc_lob : io_bxcpt_bits_uop_fetch_pc_lob; // @[rob.scala 666:32]
  wire [19:0] T_47888_imm_packed = T_47887 ? io_lxcpt_bits_uop_imm_packed : io_bxcpt_bits_uop_imm_packed; // @[rob.scala 666:32]
  wire [11:0] T_47888_csr_addr = T_47887 ? io_lxcpt_bits_uop_csr_addr : io_bxcpt_bits_uop_csr_addr; // @[rob.scala 666:32]
  wire [5:0] T_47888_rob_idx = T_47887 ? io_lxcpt_bits_uop_rob_idx : io_bxcpt_bits_uop_rob_idx; // @[rob.scala 666:32]
  wire [3:0] T_47888_ldq_idx = T_47887 ? io_lxcpt_bits_uop_ldq_idx : io_bxcpt_bits_uop_ldq_idx; // @[rob.scala 666:32]
  wire [3:0] T_47888_stq_idx = T_47887 ? io_lxcpt_bits_uop_stq_idx : io_bxcpt_bits_uop_stq_idx; // @[rob.scala 666:32]
  wire [4:0] T_47888_brob_idx = T_47887 ? io_lxcpt_bits_uop_brob_idx : io_bxcpt_bits_uop_brob_idx; // @[rob.scala 666:32]
  wire [6:0] T_47888_pdst = T_47887 ? io_lxcpt_bits_uop_pdst : io_bxcpt_bits_uop_pdst; // @[rob.scala 666:32]
  wire [6:0] T_47888_pop1 = T_47887 ? io_lxcpt_bits_uop_pop1 : io_bxcpt_bits_uop_pop1; // @[rob.scala 666:32]
  wire [6:0] T_47888_pop2 = T_47887 ? io_lxcpt_bits_uop_pop2 : io_bxcpt_bits_uop_pop2; // @[rob.scala 666:32]
  wire [6:0] T_47888_pop3 = T_47887 ? io_lxcpt_bits_uop_pop3 : io_bxcpt_bits_uop_pop3; // @[rob.scala 666:32]
  wire  T_47888_prs1_busy = T_47887 ? io_lxcpt_bits_uop_prs1_busy : io_bxcpt_bits_uop_prs1_busy; // @[rob.scala 666:32]
  wire  T_47888_prs2_busy = T_47887 ? io_lxcpt_bits_uop_prs2_busy : io_bxcpt_bits_uop_prs2_busy; // @[rob.scala 666:32]
  wire  T_47888_prs3_busy = T_47887 ? io_lxcpt_bits_uop_prs3_busy : io_bxcpt_bits_uop_prs3_busy; // @[rob.scala 666:32]
  wire [6:0] T_47888_stale_pdst = T_47887 ? io_lxcpt_bits_uop_stale_pdst : io_bxcpt_bits_uop_stale_pdst; // @[rob.scala 666:32]
  wire  T_47888_exception = T_47887 ? io_lxcpt_bits_uop_exception : io_bxcpt_bits_uop_exception; // @[rob.scala 666:32]
  wire  T_47888_bypassable = T_47887 ? io_lxcpt_bits_uop_bypassable : io_bxcpt_bits_uop_bypassable; // @[rob.scala 666:32]
  wire [3:0] T_47888_mem_cmd = T_47887 ? io_lxcpt_bits_uop_mem_cmd : io_bxcpt_bits_uop_mem_cmd; // @[rob.scala 666:32]
  wire [2:0] T_47888_mem_typ = T_47887 ? io_lxcpt_bits_uop_mem_typ : io_bxcpt_bits_uop_mem_typ; // @[rob.scala 666:32]
  wire  T_47888_is_fence = T_47887 ? io_lxcpt_bits_uop_is_fence : io_bxcpt_bits_uop_is_fence; // @[rob.scala 666:32]
  wire  T_47888_is_fencei = T_47887 ? io_lxcpt_bits_uop_is_fencei : io_bxcpt_bits_uop_is_fencei; // @[rob.scala 666:32]
  wire  T_47888_is_store = T_47887 ? io_lxcpt_bits_uop_is_store : io_bxcpt_bits_uop_is_store; // @[rob.scala 666:32]
  wire  T_47888_is_amo = T_47887 ? io_lxcpt_bits_uop_is_amo : io_bxcpt_bits_uop_is_amo; // @[rob.scala 666:32]
  wire  T_47888_is_load = T_47887 ? io_lxcpt_bits_uop_is_load : io_bxcpt_bits_uop_is_load; // @[rob.scala 666:32]
  wire  T_47888_is_unique = T_47887 ? io_lxcpt_bits_uop_is_unique : io_bxcpt_bits_uop_is_unique; // @[rob.scala 666:32]
  wire  T_47888_flush_on_commit = T_47887 ? io_lxcpt_bits_uop_flush_on_commit : io_bxcpt_bits_uop_flush_on_commit; // @[rob.scala 666:32]
  wire [5:0] T_47888_ldst = T_47887 ? io_lxcpt_bits_uop_ldst : io_bxcpt_bits_uop_ldst; // @[rob.scala 666:32]
  wire [5:0] T_47888_lrs1 = T_47887 ? io_lxcpt_bits_uop_lrs1 : io_bxcpt_bits_uop_lrs1; // @[rob.scala 666:32]
  wire [5:0] T_47888_lrs2 = T_47887 ? io_lxcpt_bits_uop_lrs2 : io_bxcpt_bits_uop_lrs2; // @[rob.scala 666:32]
  wire [5:0] T_47888_lrs3 = T_47887 ? io_lxcpt_bits_uop_lrs3 : io_bxcpt_bits_uop_lrs3; // @[rob.scala 666:32]
  wire  T_47888_ldst_val = T_47887 ? io_lxcpt_bits_uop_ldst_val : io_bxcpt_bits_uop_ldst_val; // @[rob.scala 666:32]
  wire [1:0] T_47888_dst_rtype = T_47887 ? io_lxcpt_bits_uop_dst_rtype : io_bxcpt_bits_uop_dst_rtype; // @[rob.scala 666:32]
  wire [1:0] T_47888_lrs1_rtype = T_47887 ? io_lxcpt_bits_uop_lrs1_rtype : io_bxcpt_bits_uop_lrs1_rtype; // @[rob.scala 666:32]
  wire [1:0] T_47888_lrs2_rtype = T_47887 ? io_lxcpt_bits_uop_lrs2_rtype : io_bxcpt_bits_uop_lrs2_rtype; // @[rob.scala 666:32]
  wire  T_47888_frs3_en = T_47887 ? io_lxcpt_bits_uop_frs3_en : io_bxcpt_bits_uop_frs3_en; // @[rob.scala 666:32]
  wire  T_47888_fp_val = T_47887 ? io_lxcpt_bits_uop_fp_val : io_bxcpt_bits_uop_fp_val; // @[rob.scala 666:32]
  wire  T_47888_fp_single = T_47887 ? io_lxcpt_bits_uop_fp_single : io_bxcpt_bits_uop_fp_single; // @[rob.scala 666:32]
  wire  T_47888_xcpt_if = T_47887 ? io_lxcpt_bits_uop_xcpt_if : io_bxcpt_bits_uop_xcpt_if; // @[rob.scala 666:32]
  wire  T_47888_replay_if = T_47887 ? io_lxcpt_bits_uop_replay_if : io_bxcpt_bits_uop_replay_if; // @[rob.scala 666:32]
  wire [63:0] T_47888_debug_wdata = T_47887 ? io_lxcpt_bits_uop_debug_wdata : io_bxcpt_bits_uop_debug_wdata; // @[rob.scala 666:32]
  wire [31:0] T_47888_debug_events_fetch_seq = T_47887 ? io_lxcpt_bits_uop_debug_events_fetch_seq :
    io_bxcpt_bits_uop_debug_events_fetch_seq; // @[rob.scala 666:32]
  wire  T_47975 = ~r_xcpt_val; // @[rob.scala 667:16]
  wire  T_47976 = T_47888_rob_idx <= rob_tail_idx; // @[rob.scala 650:58]
  wire [6:0] T_47977 = {T_47976,T_47888_rob_idx}; // @[Cat.scala 20:58]
  wire  T_47978 = r_xcpt_uop_rob_idx <= rob_tail_idx; // @[rob.scala 650:80]
  wire [6:0] T_47979 = {T_47978,r_xcpt_uop_rob_idx}; // @[Cat.scala 20:58]
  wire  T_47980 = T_47977 < T_47979; // @[rob.scala 650:71]
  wire  T_47981 = T_47975 | T_47980; // @[rob.scala 667:28]
  wire [3:0] T_47983 = io_lxcpt_valid ? io_lxcpt_bits_cause : io_bxcpt_bits_cause; // @[rob.scala 671:43]
  wire [39:0] T_47984 = io_lxcpt_valid ? io_lxcpt_bits_badvaddr : io_bxcpt_bits_badvaddr; // @[rob.scala 672:43]
  wire  _GEN_28319 = T_47981 | r_xcpt_val; // @[rob.scala 668:10 rob.scala 669:37]
  wire  _GEN_28320 = T_47981 ? T_47888_valid : r_xcpt_uop_valid; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [1:0] _GEN_28321 = T_47981 ? T_47888_iw_state : r_xcpt_uop_iw_state; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [8:0] _GEN_28322 = T_47981 ? T_47888_uopc : r_xcpt_uop_uopc; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [31:0] _GEN_28323 = T_47981 ? T_47888_inst : r_xcpt_uop_inst; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [39:0] _GEN_28324 = T_47981 ? T_47888_pc : r_xcpt_uop_pc; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [7:0] _GEN_28325 = T_47981 ? T_47888_fu_code : r_xcpt_uop_fu_code; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [3:0] _GEN_28326 = T_47981 ? T_47888_ctrl_br_type : r_xcpt_uop_ctrl_br_type; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [1:0] _GEN_28327 = T_47981 ? T_47888_ctrl_op1_sel : r_xcpt_uop_ctrl_op1_sel; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [2:0] _GEN_28328 = T_47981 ? T_47888_ctrl_op2_sel : r_xcpt_uop_ctrl_op2_sel; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [2:0] _GEN_28329 = T_47981 ? T_47888_ctrl_imm_sel : r_xcpt_uop_ctrl_imm_sel; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [3:0] _GEN_28330 = T_47981 ? T_47888_ctrl_op_fcn : r_xcpt_uop_ctrl_op_fcn; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28331 = T_47981 ? T_47888_ctrl_fcn_dw : r_xcpt_uop_ctrl_fcn_dw; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28332 = T_47981 ? T_47888_ctrl_rf_wen : r_xcpt_uop_ctrl_rf_wen; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [2:0] _GEN_28333 = T_47981 ? T_47888_ctrl_csr_cmd : r_xcpt_uop_ctrl_csr_cmd; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28334 = T_47981 ? T_47888_ctrl_is_load : r_xcpt_uop_ctrl_is_load; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28335 = T_47981 ? T_47888_ctrl_is_sta : r_xcpt_uop_ctrl_is_sta; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28336 = T_47981 ? T_47888_ctrl_is_std : r_xcpt_uop_ctrl_is_std; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [1:0] _GEN_28337 = T_47981 ? T_47888_wakeup_delay : r_xcpt_uop_wakeup_delay; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28338 = T_47981 ? T_47888_allocate_brtag : r_xcpt_uop_allocate_brtag; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28339 = T_47981 ? T_47888_is_br_or_jmp : r_xcpt_uop_is_br_or_jmp; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28340 = T_47981 ? T_47888_is_jump : r_xcpt_uop_is_jump; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28341 = T_47981 ? T_47888_is_jal : r_xcpt_uop_is_jal; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28342 = T_47981 ? T_47888_is_ret : r_xcpt_uop_is_ret; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28343 = T_47981 ? T_47888_is_call : r_xcpt_uop_is_call; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [7:0] _GEN_28344 = T_47981 ? T_47888_br_mask : r_xcpt_uop_br_mask; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [2:0] _GEN_28345 = T_47981 ? T_47888_br_tag : r_xcpt_uop_br_tag; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28346 = T_47981 ? T_47888_br_prediction_bpd_predict_val : r_xcpt_uop_br_prediction_bpd_predict_val; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28347 = T_47981 ? T_47888_br_prediction_bpd_predict_taken : r_xcpt_uop_br_prediction_bpd_predict_taken; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28348 = T_47981 ? T_47888_br_prediction_btb_hit : r_xcpt_uop_br_prediction_btb_hit; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28349 = T_47981 ? T_47888_br_prediction_btb_predicted : r_xcpt_uop_br_prediction_btb_predicted; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28350 = T_47981 ? T_47888_br_prediction_is_br_or_jalr : r_xcpt_uop_br_prediction_is_br_or_jalr; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28351 = T_47981 ? T_47888_stat_brjmp_mispredicted : r_xcpt_uop_stat_brjmp_mispredicted; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28352 = T_47981 ? T_47888_stat_btb_made_pred : r_xcpt_uop_stat_btb_made_pred; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28353 = T_47981 ? T_47888_stat_btb_mispredicted : r_xcpt_uop_stat_btb_mispredicted; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28354 = T_47981 ? T_47888_stat_bpd_made_pred : r_xcpt_uop_stat_bpd_made_pred; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28355 = T_47981 ? T_47888_stat_bpd_mispredicted : r_xcpt_uop_stat_bpd_mispredicted; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [2:0] _GEN_28356 = T_47981 ? T_47888_fetch_pc_lob : r_xcpt_uop_fetch_pc_lob; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [19:0] _GEN_28357 = T_47981 ? T_47888_imm_packed : r_xcpt_uop_imm_packed; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [11:0] _GEN_28358 = T_47981 ? T_47888_csr_addr : r_xcpt_uop_csr_addr; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [5:0] _GEN_28359 = T_47981 ? T_47888_rob_idx : r_xcpt_uop_rob_idx; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [3:0] _GEN_28360 = T_47981 ? T_47888_ldq_idx : r_xcpt_uop_ldq_idx; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [3:0] _GEN_28361 = T_47981 ? T_47888_stq_idx : r_xcpt_uop_stq_idx; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [4:0] _GEN_28362 = T_47981 ? T_47888_brob_idx : r_xcpt_uop_brob_idx; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [6:0] _GEN_28363 = T_47981 ? T_47888_pdst : r_xcpt_uop_pdst; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [6:0] _GEN_28364 = T_47981 ? T_47888_pop1 : r_xcpt_uop_pop1; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [6:0] _GEN_28365 = T_47981 ? T_47888_pop2 : r_xcpt_uop_pop2; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [6:0] _GEN_28366 = T_47981 ? T_47888_pop3 : r_xcpt_uop_pop3; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28367 = T_47981 ? T_47888_prs1_busy : r_xcpt_uop_prs1_busy; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28368 = T_47981 ? T_47888_prs2_busy : r_xcpt_uop_prs2_busy; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28369 = T_47981 ? T_47888_prs3_busy : r_xcpt_uop_prs3_busy; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [6:0] _GEN_28370 = T_47981 ? T_47888_stale_pdst : r_xcpt_uop_stale_pdst; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28371 = T_47981 ? T_47888_exception : r_xcpt_uop_exception; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [63:0] _GEN_28372 = T_47981 ? {{60'd0}, T_47983} : r_xcpt_uop_exc_cause; // @[rob.scala 668:10 rob.scala 671:37 rob.scala 652:18]
  wire  _GEN_28373 = T_47981 ? T_47888_bypassable : r_xcpt_uop_bypassable; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [3:0] _GEN_28374 = T_47981 ? T_47888_mem_cmd : r_xcpt_uop_mem_cmd; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [2:0] _GEN_28375 = T_47981 ? T_47888_mem_typ : r_xcpt_uop_mem_typ; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28376 = T_47981 ? T_47888_is_fence : r_xcpt_uop_is_fence; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28377 = T_47981 ? T_47888_is_fencei : r_xcpt_uop_is_fencei; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28378 = T_47981 ? T_47888_is_store : r_xcpt_uop_is_store; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28379 = T_47981 ? T_47888_is_amo : r_xcpt_uop_is_amo; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28380 = T_47981 ? T_47888_is_load : r_xcpt_uop_is_load; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28381 = T_47981 ? T_47888_is_unique : r_xcpt_uop_is_unique; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28382 = T_47981 ? T_47888_flush_on_commit : r_xcpt_uop_flush_on_commit; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [5:0] _GEN_28383 = T_47981 ? T_47888_ldst : r_xcpt_uop_ldst; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [5:0] _GEN_28384 = T_47981 ? T_47888_lrs1 : r_xcpt_uop_lrs1; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [5:0] _GEN_28385 = T_47981 ? T_47888_lrs2 : r_xcpt_uop_lrs2; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [5:0] _GEN_28386 = T_47981 ? T_47888_lrs3 : r_xcpt_uop_lrs3; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28387 = T_47981 ? T_47888_ldst_val : r_xcpt_uop_ldst_val; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [1:0] _GEN_28388 = T_47981 ? T_47888_dst_rtype : r_xcpt_uop_dst_rtype; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [1:0] _GEN_28389 = T_47981 ? T_47888_lrs1_rtype : r_xcpt_uop_lrs1_rtype; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [1:0] _GEN_28390 = T_47981 ? T_47888_lrs2_rtype : r_xcpt_uop_lrs2_rtype; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28391 = T_47981 ? T_47888_frs3_en : r_xcpt_uop_frs3_en; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28392 = T_47981 ? T_47888_fp_val : r_xcpt_uop_fp_val; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28393 = T_47981 ? T_47888_fp_single : r_xcpt_uop_fp_single; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28394 = T_47981 ? T_47888_xcpt_if : r_xcpt_uop_xcpt_if; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28395 = T_47981 ? T_47888_replay_if : r_xcpt_uop_replay_if; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [63:0] _GEN_28396 = T_47981 ? T_47888_debug_wdata : r_xcpt_uop_debug_wdata; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire [31:0] _GEN_28397 = T_47981 ? T_47888_debug_events_fetch_seq : r_xcpt_uop_debug_events_fetch_seq; // @[rob.scala 668:10 rob.scala 670:37 rob.scala 652:18]
  wire  _GEN_28399 = T_47876 ? _GEN_28319 : r_xcpt_val; // @[rob.scala 662:7]
  wire  _GEN_28400 = T_47876 ? _GEN_28320 : r_xcpt_uop_valid; // @[rob.scala 662:7 rob.scala 652:18]
  wire [1:0] _GEN_28401 = T_47876 ? _GEN_28321 : r_xcpt_uop_iw_state; // @[rob.scala 662:7 rob.scala 652:18]
  wire [8:0] _GEN_28402 = T_47876 ? _GEN_28322 : r_xcpt_uop_uopc; // @[rob.scala 662:7 rob.scala 652:18]
  wire [31:0] _GEN_28403 = T_47876 ? _GEN_28323 : r_xcpt_uop_inst; // @[rob.scala 662:7 rob.scala 652:18]
  wire [39:0] _GEN_28404 = T_47876 ? _GEN_28324 : r_xcpt_uop_pc; // @[rob.scala 662:7 rob.scala 652:18]
  wire [7:0] _GEN_28405 = T_47876 ? _GEN_28325 : r_xcpt_uop_fu_code; // @[rob.scala 662:7 rob.scala 652:18]
  wire [3:0] _GEN_28406 = T_47876 ? _GEN_28326 : r_xcpt_uop_ctrl_br_type; // @[rob.scala 662:7 rob.scala 652:18]
  wire [1:0] _GEN_28407 = T_47876 ? _GEN_28327 : r_xcpt_uop_ctrl_op1_sel; // @[rob.scala 662:7 rob.scala 652:18]
  wire [2:0] _GEN_28408 = T_47876 ? _GEN_28328 : r_xcpt_uop_ctrl_op2_sel; // @[rob.scala 662:7 rob.scala 652:18]
  wire [2:0] _GEN_28409 = T_47876 ? _GEN_28329 : r_xcpt_uop_ctrl_imm_sel; // @[rob.scala 662:7 rob.scala 652:18]
  wire [3:0] _GEN_28410 = T_47876 ? _GEN_28330 : r_xcpt_uop_ctrl_op_fcn; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28411 = T_47876 ? _GEN_28331 : r_xcpt_uop_ctrl_fcn_dw; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28412 = T_47876 ? _GEN_28332 : r_xcpt_uop_ctrl_rf_wen; // @[rob.scala 662:7 rob.scala 652:18]
  wire [2:0] _GEN_28413 = T_47876 ? _GEN_28333 : r_xcpt_uop_ctrl_csr_cmd; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28414 = T_47876 ? _GEN_28334 : r_xcpt_uop_ctrl_is_load; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28415 = T_47876 ? _GEN_28335 : r_xcpt_uop_ctrl_is_sta; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28416 = T_47876 ? _GEN_28336 : r_xcpt_uop_ctrl_is_std; // @[rob.scala 662:7 rob.scala 652:18]
  wire [1:0] _GEN_28417 = T_47876 ? _GEN_28337 : r_xcpt_uop_wakeup_delay; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28418 = T_47876 ? _GEN_28338 : r_xcpt_uop_allocate_brtag; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28419 = T_47876 ? _GEN_28339 : r_xcpt_uop_is_br_or_jmp; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28420 = T_47876 ? _GEN_28340 : r_xcpt_uop_is_jump; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28421 = T_47876 ? _GEN_28341 : r_xcpt_uop_is_jal; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28422 = T_47876 ? _GEN_28342 : r_xcpt_uop_is_ret; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28423 = T_47876 ? _GEN_28343 : r_xcpt_uop_is_call; // @[rob.scala 662:7 rob.scala 652:18]
  wire [7:0] _GEN_28424 = T_47876 ? _GEN_28344 : r_xcpt_uop_br_mask; // @[rob.scala 662:7 rob.scala 652:18]
  wire [2:0] _GEN_28425 = T_47876 ? _GEN_28345 : r_xcpt_uop_br_tag; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28426 = T_47876 ? _GEN_28346 : r_xcpt_uop_br_prediction_bpd_predict_val; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28427 = T_47876 ? _GEN_28347 : r_xcpt_uop_br_prediction_bpd_predict_taken; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28428 = T_47876 ? _GEN_28348 : r_xcpt_uop_br_prediction_btb_hit; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28429 = T_47876 ? _GEN_28349 : r_xcpt_uop_br_prediction_btb_predicted; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28430 = T_47876 ? _GEN_28350 : r_xcpt_uop_br_prediction_is_br_or_jalr; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28431 = T_47876 ? _GEN_28351 : r_xcpt_uop_stat_brjmp_mispredicted; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28432 = T_47876 ? _GEN_28352 : r_xcpt_uop_stat_btb_made_pred; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28433 = T_47876 ? _GEN_28353 : r_xcpt_uop_stat_btb_mispredicted; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28434 = T_47876 ? _GEN_28354 : r_xcpt_uop_stat_bpd_made_pred; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28435 = T_47876 ? _GEN_28355 : r_xcpt_uop_stat_bpd_mispredicted; // @[rob.scala 662:7 rob.scala 652:18]
  wire [2:0] _GEN_28436 = T_47876 ? _GEN_28356 : r_xcpt_uop_fetch_pc_lob; // @[rob.scala 662:7 rob.scala 652:18]
  wire [19:0] _GEN_28437 = T_47876 ? _GEN_28357 : r_xcpt_uop_imm_packed; // @[rob.scala 662:7 rob.scala 652:18]
  wire [11:0] _GEN_28438 = T_47876 ? _GEN_28358 : r_xcpt_uop_csr_addr; // @[rob.scala 662:7 rob.scala 652:18]
  wire [5:0] _GEN_28439 = T_47876 ? _GEN_28359 : r_xcpt_uop_rob_idx; // @[rob.scala 662:7 rob.scala 652:18]
  wire [3:0] _GEN_28440 = T_47876 ? _GEN_28360 : r_xcpt_uop_ldq_idx; // @[rob.scala 662:7 rob.scala 652:18]
  wire [3:0] _GEN_28441 = T_47876 ? _GEN_28361 : r_xcpt_uop_stq_idx; // @[rob.scala 662:7 rob.scala 652:18]
  wire [4:0] _GEN_28442 = T_47876 ? _GEN_28362 : r_xcpt_uop_brob_idx; // @[rob.scala 662:7 rob.scala 652:18]
  wire [6:0] _GEN_28443 = T_47876 ? _GEN_28363 : r_xcpt_uop_pdst; // @[rob.scala 662:7 rob.scala 652:18]
  wire [6:0] _GEN_28444 = T_47876 ? _GEN_28364 : r_xcpt_uop_pop1; // @[rob.scala 662:7 rob.scala 652:18]
  wire [6:0] _GEN_28445 = T_47876 ? _GEN_28365 : r_xcpt_uop_pop2; // @[rob.scala 662:7 rob.scala 652:18]
  wire [6:0] _GEN_28446 = T_47876 ? _GEN_28366 : r_xcpt_uop_pop3; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28447 = T_47876 ? _GEN_28367 : r_xcpt_uop_prs1_busy; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28448 = T_47876 ? _GEN_28368 : r_xcpt_uop_prs2_busy; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28449 = T_47876 ? _GEN_28369 : r_xcpt_uop_prs3_busy; // @[rob.scala 662:7 rob.scala 652:18]
  wire [6:0] _GEN_28450 = T_47876 ? _GEN_28370 : r_xcpt_uop_stale_pdst; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28451 = T_47876 ? _GEN_28371 : r_xcpt_uop_exception; // @[rob.scala 662:7 rob.scala 652:18]
  wire [63:0] _GEN_28452 = T_47876 ? _GEN_28372 : r_xcpt_uop_exc_cause; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28453 = T_47876 ? _GEN_28373 : r_xcpt_uop_bypassable; // @[rob.scala 662:7 rob.scala 652:18]
  wire [3:0] _GEN_28454 = T_47876 ? _GEN_28374 : r_xcpt_uop_mem_cmd; // @[rob.scala 662:7 rob.scala 652:18]
  wire [2:0] _GEN_28455 = T_47876 ? _GEN_28375 : r_xcpt_uop_mem_typ; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28456 = T_47876 ? _GEN_28376 : r_xcpt_uop_is_fence; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28457 = T_47876 ? _GEN_28377 : r_xcpt_uop_is_fencei; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28458 = T_47876 ? _GEN_28378 : r_xcpt_uop_is_store; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28459 = T_47876 ? _GEN_28379 : r_xcpt_uop_is_amo; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28460 = T_47876 ? _GEN_28380 : r_xcpt_uop_is_load; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28461 = T_47876 ? _GEN_28381 : r_xcpt_uop_is_unique; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28462 = T_47876 ? _GEN_28382 : r_xcpt_uop_flush_on_commit; // @[rob.scala 662:7 rob.scala 652:18]
  wire [5:0] _GEN_28463 = T_47876 ? _GEN_28383 : r_xcpt_uop_ldst; // @[rob.scala 662:7 rob.scala 652:18]
  wire [5:0] _GEN_28464 = T_47876 ? _GEN_28384 : r_xcpt_uop_lrs1; // @[rob.scala 662:7 rob.scala 652:18]
  wire [5:0] _GEN_28465 = T_47876 ? _GEN_28385 : r_xcpt_uop_lrs2; // @[rob.scala 662:7 rob.scala 652:18]
  wire [5:0] _GEN_28466 = T_47876 ? _GEN_28386 : r_xcpt_uop_lrs3; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28467 = T_47876 ? _GEN_28387 : r_xcpt_uop_ldst_val; // @[rob.scala 662:7 rob.scala 652:18]
  wire [1:0] _GEN_28468 = T_47876 ? _GEN_28388 : r_xcpt_uop_dst_rtype; // @[rob.scala 662:7 rob.scala 652:18]
  wire [1:0] _GEN_28469 = T_47876 ? _GEN_28389 : r_xcpt_uop_lrs1_rtype; // @[rob.scala 662:7 rob.scala 652:18]
  wire [1:0] _GEN_28470 = T_47876 ? _GEN_28390 : r_xcpt_uop_lrs2_rtype; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28471 = T_47876 ? _GEN_28391 : r_xcpt_uop_frs3_en; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28472 = T_47876 ? _GEN_28392 : r_xcpt_uop_fp_val; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28473 = T_47876 ? _GEN_28393 : r_xcpt_uop_fp_single; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28474 = T_47876 ? _GEN_28394 : r_xcpt_uop_xcpt_if; // @[rob.scala 662:7 rob.scala 652:18]
  wire  _GEN_28475 = T_47876 ? _GEN_28395 : r_xcpt_uop_replay_if; // @[rob.scala 662:7 rob.scala 652:18]
  wire [63:0] _GEN_28476 = T_47876 ? _GEN_28396 : r_xcpt_uop_debug_wdata; // @[rob.scala 662:7 rob.scala 652:18]
  wire [31:0] _GEN_28477 = T_47876 ? _GEN_28397 : r_xcpt_uop_debug_events_fetch_seq; // @[rob.scala 662:7 rob.scala 652:18]
  wire  T_47987 = T_47869 | T_47870; // @[rob.scala 675:51]
  wire  T_47988 = T_47975 & T_47987; // @[rob.scala 675:30]
  wire  T_47990 = ~T_47876; // @[rob.scala 662:7]
  wire  T_47991 = T_47990 & T_47988; // @[rob.scala 676:7]
  wire  T_47994 = T_47869 ? 1'h0 : 1'h1; // @[rob.scala 677:40]
  wire  _GEN_28557 = T_47994 ? io_dis_uops_1_valid : io_dis_uops_0_valid; // @[rob.scala 681:26 rob.scala 681:26]
  wire [1:0] _GEN_28558 = T_47994 ? io_dis_uops_1_iw_state : io_dis_uops_0_iw_state; // @[rob.scala 681:26 rob.scala 681:26]
  wire [8:0] _GEN_28559 = T_47994 ? io_dis_uops_1_uopc : io_dis_uops_0_uopc; // @[rob.scala 681:26 rob.scala 681:26]
  wire [31:0] _GEN_28560 = T_47994 ? io_dis_uops_1_inst : io_dis_uops_0_inst; // @[rob.scala 681:26 rob.scala 681:26]
  wire [39:0] _GEN_28561 = T_47994 ? io_dis_uops_1_pc : io_dis_uops_0_pc; // @[rob.scala 681:26 rob.scala 681:26]
  wire [7:0] _GEN_28562 = T_47994 ? io_dis_uops_1_fu_code : io_dis_uops_0_fu_code; // @[rob.scala 681:26 rob.scala 681:26]
  wire [3:0] _GEN_28563 = T_47994 ? io_dis_uops_1_ctrl_br_type : io_dis_uops_0_ctrl_br_type; // @[rob.scala 681:26 rob.scala 681:26]
  wire [1:0] _GEN_28564 = T_47994 ? io_dis_uops_1_ctrl_op1_sel : io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28565 = T_47994 ? io_dis_uops_1_ctrl_op2_sel : io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28566 = T_47994 ? io_dis_uops_1_ctrl_imm_sel : io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 681:26 rob.scala 681:26]
  wire [3:0] _GEN_28567 = T_47994 ? io_dis_uops_1_ctrl_op_fcn : io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28568 = T_47994 ? io_dis_uops_1_ctrl_fcn_dw : io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28569 = T_47994 ? io_dis_uops_1_ctrl_rf_wen : io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28570 = T_47994 ? io_dis_uops_1_ctrl_csr_cmd : io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28571 = T_47994 ? io_dis_uops_1_ctrl_is_load : io_dis_uops_0_ctrl_is_load; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28572 = T_47994 ? io_dis_uops_1_ctrl_is_sta : io_dis_uops_0_ctrl_is_sta; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28573 = T_47994 ? io_dis_uops_1_ctrl_is_std : io_dis_uops_0_ctrl_is_std; // @[rob.scala 681:26 rob.scala 681:26]
  wire [1:0] _GEN_28574 = T_47994 ? io_dis_uops_1_wakeup_delay : io_dis_uops_0_wakeup_delay; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28575 = T_47994 ? io_dis_uops_1_allocate_brtag : io_dis_uops_0_allocate_brtag; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28576 = T_47994 ? io_dis_uops_1_is_br_or_jmp : io_dis_uops_0_is_br_or_jmp; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28577 = T_47994 ? io_dis_uops_1_is_jump : io_dis_uops_0_is_jump; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28578 = T_47994 ? io_dis_uops_1_is_jal : io_dis_uops_0_is_jal; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28579 = T_47994 ? io_dis_uops_1_is_ret : io_dis_uops_0_is_ret; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28580 = T_47994 ? io_dis_uops_1_is_call : io_dis_uops_0_is_call; // @[rob.scala 681:26 rob.scala 681:26]
  wire [7:0] _GEN_28581 = T_47994 ? io_dis_uops_1_br_mask : io_dis_uops_0_br_mask; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28582 = T_47994 ? io_dis_uops_1_br_tag : io_dis_uops_0_br_tag; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28583 = T_47994 ? io_dis_uops_1_br_prediction_bpd_predict_val : io_dis_uops_0_br_prediction_bpd_predict_val
    ; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28584 = T_47994 ? io_dis_uops_1_br_prediction_bpd_predict_taken :
    io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28585 = T_47994 ? io_dis_uops_1_br_prediction_btb_hit : io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28586 = T_47994 ? io_dis_uops_1_br_prediction_btb_predicted : io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28587 = T_47994 ? io_dis_uops_1_br_prediction_is_br_or_jalr : io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28588 = T_47994 ? io_dis_uops_1_stat_brjmp_mispredicted : io_dis_uops_0_stat_brjmp_mispredicted; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28589 = T_47994 ? io_dis_uops_1_stat_btb_made_pred : io_dis_uops_0_stat_btb_made_pred; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28590 = T_47994 ? io_dis_uops_1_stat_btb_mispredicted : io_dis_uops_0_stat_btb_mispredicted; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28591 = T_47994 ? io_dis_uops_1_stat_bpd_made_pred : io_dis_uops_0_stat_bpd_made_pred; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28592 = T_47994 ? io_dis_uops_1_stat_bpd_mispredicted : io_dis_uops_0_stat_bpd_mispredicted; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28593 = T_47994 ? io_dis_uops_1_fetch_pc_lob : io_dis_uops_0_fetch_pc_lob; // @[rob.scala 681:26 rob.scala 681:26]
  wire [19:0] _GEN_28594 = T_47994 ? io_dis_uops_1_imm_packed : io_dis_uops_0_imm_packed; // @[rob.scala 681:26 rob.scala 681:26]
  wire [11:0] _GEN_28595 = T_47994 ? io_dis_uops_1_csr_addr : io_dis_uops_0_csr_addr; // @[rob.scala 681:26 rob.scala 681:26]
  wire [5:0] _GEN_28596 = T_47994 ? io_dis_uops_1_rob_idx : io_dis_uops_0_rob_idx; // @[rob.scala 681:26 rob.scala 681:26]
  wire [3:0] _GEN_28597 = T_47994 ? io_dis_uops_1_ldq_idx : io_dis_uops_0_ldq_idx; // @[rob.scala 681:26 rob.scala 681:26]
  wire [3:0] _GEN_28598 = T_47994 ? io_dis_uops_1_stq_idx : io_dis_uops_0_stq_idx; // @[rob.scala 681:26 rob.scala 681:26]
  wire [4:0] _GEN_28599 = T_47994 ? io_dis_uops_1_brob_idx : io_dis_uops_0_brob_idx; // @[rob.scala 681:26 rob.scala 681:26]
  wire [6:0] _GEN_28600 = T_47994 ? io_dis_uops_1_pdst : io_dis_uops_0_pdst; // @[rob.scala 681:26 rob.scala 681:26]
  wire [6:0] _GEN_28601 = T_47994 ? io_dis_uops_1_pop1 : io_dis_uops_0_pop1; // @[rob.scala 681:26 rob.scala 681:26]
  wire [6:0] _GEN_28602 = T_47994 ? io_dis_uops_1_pop2 : io_dis_uops_0_pop2; // @[rob.scala 681:26 rob.scala 681:26]
  wire [6:0] _GEN_28603 = T_47994 ? io_dis_uops_1_pop3 : io_dis_uops_0_pop3; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28604 = T_47994 ? io_dis_uops_1_prs1_busy : io_dis_uops_0_prs1_busy; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28605 = T_47994 ? io_dis_uops_1_prs2_busy : io_dis_uops_0_prs2_busy; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28606 = T_47994 ? io_dis_uops_1_prs3_busy : io_dis_uops_0_prs3_busy; // @[rob.scala 681:26 rob.scala 681:26]
  wire [6:0] _GEN_28607 = T_47994 ? io_dis_uops_1_stale_pdst : io_dis_uops_0_stale_pdst; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28608 = T_47994 ? io_dis_uops_1_exception : io_dis_uops_0_exception; // @[rob.scala 681:26 rob.scala 681:26]
  wire [63:0] _GEN_28609 = T_47994 ? io_dis_uops_1_exc_cause : io_dis_uops_0_exc_cause; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28610 = T_47994 ? io_dis_uops_1_bypassable : io_dis_uops_0_bypassable; // @[rob.scala 681:26 rob.scala 681:26]
  wire [3:0] _GEN_28611 = T_47994 ? io_dis_uops_1_mem_cmd : io_dis_uops_0_mem_cmd; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28612 = T_47994 ? io_dis_uops_1_mem_typ : io_dis_uops_0_mem_typ; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28613 = T_47994 ? io_dis_uops_1_is_fence : io_dis_uops_0_is_fence; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28614 = T_47994 ? io_dis_uops_1_is_fencei : io_dis_uops_0_is_fencei; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28615 = T_47994 ? io_dis_uops_1_is_store : io_dis_uops_0_is_store; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28616 = T_47994 ? io_dis_uops_1_is_amo : io_dis_uops_0_is_amo; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28617 = T_47994 ? io_dis_uops_1_is_load : io_dis_uops_0_is_load; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28618 = T_47994 ? io_dis_uops_1_is_unique : io_dis_uops_0_is_unique; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28619 = T_47994 ? io_dis_uops_1_flush_on_commit : io_dis_uops_0_flush_on_commit; // @[rob.scala 681:26 rob.scala 681:26]
  wire [5:0] _GEN_28620 = T_47994 ? io_dis_uops_1_ldst : io_dis_uops_0_ldst; // @[rob.scala 681:26 rob.scala 681:26]
  wire [5:0] _GEN_28621 = T_47994 ? io_dis_uops_1_lrs1 : io_dis_uops_0_lrs1; // @[rob.scala 681:26 rob.scala 681:26]
  wire [5:0] _GEN_28622 = T_47994 ? io_dis_uops_1_lrs2 : io_dis_uops_0_lrs2; // @[rob.scala 681:26 rob.scala 681:26]
  wire [5:0] _GEN_28623 = T_47994 ? io_dis_uops_1_lrs3 : io_dis_uops_0_lrs3; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28624 = T_47994 ? io_dis_uops_1_ldst_val : io_dis_uops_0_ldst_val; // @[rob.scala 681:26 rob.scala 681:26]
  wire [1:0] _GEN_28625 = T_47994 ? io_dis_uops_1_dst_rtype : io_dis_uops_0_dst_rtype; // @[rob.scala 681:26 rob.scala 681:26]
  wire [1:0] _GEN_28626 = T_47994 ? io_dis_uops_1_lrs1_rtype : io_dis_uops_0_lrs1_rtype; // @[rob.scala 681:26 rob.scala 681:26]
  wire [1:0] _GEN_28627 = T_47994 ? io_dis_uops_1_lrs2_rtype : io_dis_uops_0_lrs2_rtype; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28628 = T_47994 ? io_dis_uops_1_frs3_en : io_dis_uops_0_frs3_en; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28629 = T_47994 ? io_dis_uops_1_fp_val : io_dis_uops_0_fp_val; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28630 = T_47994 ? io_dis_uops_1_fp_single : io_dis_uops_0_fp_single; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28631 = T_47994 ? io_dis_uops_1_xcpt_if : io_dis_uops_0_xcpt_if; // @[rob.scala 681:26 rob.scala 681:26]
  wire  _GEN_28632 = T_47994 ? io_dis_uops_1_replay_if : io_dis_uops_0_replay_if; // @[rob.scala 681:26 rob.scala 681:26]
  wire [63:0] _GEN_28633 = T_47994 ? io_dis_uops_1_debug_wdata : io_dis_uops_0_debug_wdata; // @[rob.scala 681:26 rob.scala 681:26]
  wire [31:0] _GEN_28634 = T_47994 ? io_dis_uops_1_debug_events_fetch_seq : io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 681:26 rob.scala 681:26]
  wire [2:0] _GEN_28922 = {T_47994, 2'h0}; // @[rob.scala 682:54]
  wire [3:0] T_48082 = {{1'd0}, _GEN_28922}; // @[rob.scala 682:54]
  wire [39:0] _GEN_28923 = {{36'd0}, T_48082}; // @[rob.scala 682:47]
  wire [39:0] T_48084 = io_dis_uops_0_pc + _GEN_28923; // @[rob.scala 682:47]
  wire  _GEN_28635 = T_47991 | _GEN_28399; // @[rob.scala 676:7 rob.scala 680:26]
  wire  _GEN_28636 = T_47991 ? _GEN_28557 : _GEN_28400; // @[rob.scala 676:7 rob.scala 681:26]
  wire [1:0] _GEN_28637 = T_47991 ? _GEN_28558 : _GEN_28401; // @[rob.scala 676:7 rob.scala 681:26]
  wire [8:0] _GEN_28638 = T_47991 ? _GEN_28559 : _GEN_28402; // @[rob.scala 676:7 rob.scala 681:26]
  wire [31:0] _GEN_28639 = T_47991 ? _GEN_28560 : _GEN_28403; // @[rob.scala 676:7 rob.scala 681:26]
  wire [39:0] _GEN_28640 = T_47991 ? _GEN_28561 : _GEN_28404; // @[rob.scala 676:7 rob.scala 681:26]
  wire [7:0] _GEN_28641 = T_47991 ? _GEN_28562 : _GEN_28405; // @[rob.scala 676:7 rob.scala 681:26]
  wire [3:0] _GEN_28642 = T_47991 ? _GEN_28563 : _GEN_28406; // @[rob.scala 676:7 rob.scala 681:26]
  wire [1:0] _GEN_28643 = T_47991 ? _GEN_28564 : _GEN_28407; // @[rob.scala 676:7 rob.scala 681:26]
  wire [2:0] _GEN_28644 = T_47991 ? _GEN_28565 : _GEN_28408; // @[rob.scala 676:7 rob.scala 681:26]
  wire [2:0] _GEN_28645 = T_47991 ? _GEN_28566 : _GEN_28409; // @[rob.scala 676:7 rob.scala 681:26]
  wire [3:0] _GEN_28646 = T_47991 ? _GEN_28567 : _GEN_28410; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28647 = T_47991 ? _GEN_28568 : _GEN_28411; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28648 = T_47991 ? _GEN_28569 : _GEN_28412; // @[rob.scala 676:7 rob.scala 681:26]
  wire [2:0] _GEN_28649 = T_47991 ? _GEN_28570 : _GEN_28413; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28650 = T_47991 ? _GEN_28571 : _GEN_28414; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28651 = T_47991 ? _GEN_28572 : _GEN_28415; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28652 = T_47991 ? _GEN_28573 : _GEN_28416; // @[rob.scala 676:7 rob.scala 681:26]
  wire [1:0] _GEN_28653 = T_47991 ? _GEN_28574 : _GEN_28417; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28654 = T_47991 ? _GEN_28575 : _GEN_28418; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28655 = T_47991 ? _GEN_28576 : _GEN_28419; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28656 = T_47991 ? _GEN_28577 : _GEN_28420; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28657 = T_47991 ? _GEN_28578 : _GEN_28421; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28658 = T_47991 ? _GEN_28579 : _GEN_28422; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28659 = T_47991 ? _GEN_28580 : _GEN_28423; // @[rob.scala 676:7 rob.scala 681:26]
  wire [7:0] _GEN_28660 = T_47991 ? _GEN_28581 : _GEN_28424; // @[rob.scala 676:7 rob.scala 681:26]
  wire [2:0] _GEN_28661 = T_47991 ? _GEN_28582 : _GEN_28425; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28662 = T_47991 ? _GEN_28583 : _GEN_28426; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28663 = T_47991 ? _GEN_28584 : _GEN_28427; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28664 = T_47991 ? _GEN_28585 : _GEN_28428; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28665 = T_47991 ? _GEN_28586 : _GEN_28429; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28666 = T_47991 ? _GEN_28587 : _GEN_28430; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28667 = T_47991 ? _GEN_28588 : _GEN_28431; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28668 = T_47991 ? _GEN_28589 : _GEN_28432; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28669 = T_47991 ? _GEN_28590 : _GEN_28433; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28670 = T_47991 ? _GEN_28591 : _GEN_28434; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28671 = T_47991 ? _GEN_28592 : _GEN_28435; // @[rob.scala 676:7 rob.scala 681:26]
  wire [2:0] _GEN_28672 = T_47991 ? _GEN_28593 : _GEN_28436; // @[rob.scala 676:7 rob.scala 681:26]
  wire [19:0] _GEN_28673 = T_47991 ? _GEN_28594 : _GEN_28437; // @[rob.scala 676:7 rob.scala 681:26]
  wire [11:0] _GEN_28674 = T_47991 ? _GEN_28595 : _GEN_28438; // @[rob.scala 676:7 rob.scala 681:26]
  wire [5:0] _GEN_28675 = T_47991 ? _GEN_28596 : _GEN_28439; // @[rob.scala 676:7 rob.scala 681:26]
  wire [3:0] _GEN_28676 = T_47991 ? _GEN_28597 : _GEN_28440; // @[rob.scala 676:7 rob.scala 681:26]
  wire [3:0] _GEN_28677 = T_47991 ? _GEN_28598 : _GEN_28441; // @[rob.scala 676:7 rob.scala 681:26]
  wire [4:0] _GEN_28678 = T_47991 ? _GEN_28599 : _GEN_28442; // @[rob.scala 676:7 rob.scala 681:26]
  wire [6:0] _GEN_28679 = T_47991 ? _GEN_28600 : _GEN_28443; // @[rob.scala 676:7 rob.scala 681:26]
  wire [6:0] _GEN_28680 = T_47991 ? _GEN_28601 : _GEN_28444; // @[rob.scala 676:7 rob.scala 681:26]
  wire [6:0] _GEN_28681 = T_47991 ? _GEN_28602 : _GEN_28445; // @[rob.scala 676:7 rob.scala 681:26]
  wire [6:0] _GEN_28682 = T_47991 ? _GEN_28603 : _GEN_28446; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28683 = T_47991 ? _GEN_28604 : _GEN_28447; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28684 = T_47991 ? _GEN_28605 : _GEN_28448; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28685 = T_47991 ? _GEN_28606 : _GEN_28449; // @[rob.scala 676:7 rob.scala 681:26]
  wire [6:0] _GEN_28686 = T_47991 ? _GEN_28607 : _GEN_28450; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28687 = T_47991 ? _GEN_28608 : _GEN_28451; // @[rob.scala 676:7 rob.scala 681:26]
  wire [63:0] _GEN_28688 = T_47991 ? _GEN_28609 : _GEN_28452; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28689 = T_47991 ? _GEN_28610 : _GEN_28453; // @[rob.scala 676:7 rob.scala 681:26]
  wire [3:0] _GEN_28690 = T_47991 ? _GEN_28611 : _GEN_28454; // @[rob.scala 676:7 rob.scala 681:26]
  wire [2:0] _GEN_28691 = T_47991 ? _GEN_28612 : _GEN_28455; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28692 = T_47991 ? _GEN_28613 : _GEN_28456; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28693 = T_47991 ? _GEN_28614 : _GEN_28457; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28694 = T_47991 ? _GEN_28615 : _GEN_28458; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28695 = T_47991 ? _GEN_28616 : _GEN_28459; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28696 = T_47991 ? _GEN_28617 : _GEN_28460; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28697 = T_47991 ? _GEN_28618 : _GEN_28461; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28698 = T_47991 ? _GEN_28619 : _GEN_28462; // @[rob.scala 676:7 rob.scala 681:26]
  wire [5:0] _GEN_28699 = T_47991 ? _GEN_28620 : _GEN_28463; // @[rob.scala 676:7 rob.scala 681:26]
  wire [5:0] _GEN_28700 = T_47991 ? _GEN_28621 : _GEN_28464; // @[rob.scala 676:7 rob.scala 681:26]
  wire [5:0] _GEN_28701 = T_47991 ? _GEN_28622 : _GEN_28465; // @[rob.scala 676:7 rob.scala 681:26]
  wire [5:0] _GEN_28702 = T_47991 ? _GEN_28623 : _GEN_28466; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28703 = T_47991 ? _GEN_28624 : _GEN_28467; // @[rob.scala 676:7 rob.scala 681:26]
  wire [1:0] _GEN_28704 = T_47991 ? _GEN_28625 : _GEN_28468; // @[rob.scala 676:7 rob.scala 681:26]
  wire [1:0] _GEN_28705 = T_47991 ? _GEN_28626 : _GEN_28469; // @[rob.scala 676:7 rob.scala 681:26]
  wire [1:0] _GEN_28706 = T_47991 ? _GEN_28627 : _GEN_28470; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28707 = T_47991 ? _GEN_28628 : _GEN_28471; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28708 = T_47991 ? _GEN_28629 : _GEN_28472; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28709 = T_47991 ? _GEN_28630 : _GEN_28473; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28710 = T_47991 ? _GEN_28631 : _GEN_28474; // @[rob.scala 676:7 rob.scala 681:26]
  wire  _GEN_28711 = T_47991 ? _GEN_28632 : _GEN_28475; // @[rob.scala 676:7 rob.scala 681:26]
  wire [63:0] _GEN_28712 = T_47991 ? _GEN_28633 : _GEN_28476; // @[rob.scala 676:7 rob.scala 681:26]
  wire [31:0] _GEN_28713 = T_47991 ? _GEN_28634 : _GEN_28477; // @[rob.scala 676:7 rob.scala 681:26]
  wire  next_xcpt_uop_valid = T_47875 ? _GEN_28636 : r_xcpt_uop_valid; // @[rob.scala 660:4 rob.scala 652:18]
  wire [1:0] next_xcpt_uop_iw_state = T_47875 ? _GEN_28637 : r_xcpt_uop_iw_state; // @[rob.scala 660:4 rob.scala 652:18]
  wire [8:0] next_xcpt_uop_uopc = T_47875 ? _GEN_28638 : r_xcpt_uop_uopc; // @[rob.scala 660:4 rob.scala 652:18]
  wire [31:0] next_xcpt_uop_inst = T_47875 ? _GEN_28639 : r_xcpt_uop_inst; // @[rob.scala 660:4 rob.scala 652:18]
  wire [39:0] next_xcpt_uop_pc = T_47875 ? _GEN_28640 : r_xcpt_uop_pc; // @[rob.scala 660:4 rob.scala 652:18]
  wire [7:0] next_xcpt_uop_fu_code = T_47875 ? _GEN_28641 : r_xcpt_uop_fu_code; // @[rob.scala 660:4 rob.scala 652:18]
  wire [3:0] next_xcpt_uop_ctrl_br_type = T_47875 ? _GEN_28642 : r_xcpt_uop_ctrl_br_type; // @[rob.scala 660:4 rob.scala 652:18]
  wire [1:0] next_xcpt_uop_ctrl_op1_sel = T_47875 ? _GEN_28643 : r_xcpt_uop_ctrl_op1_sel; // @[rob.scala 660:4 rob.scala 652:18]
  wire [2:0] next_xcpt_uop_ctrl_op2_sel = T_47875 ? _GEN_28644 : r_xcpt_uop_ctrl_op2_sel; // @[rob.scala 660:4 rob.scala 652:18]
  wire [2:0] next_xcpt_uop_ctrl_imm_sel = T_47875 ? _GEN_28645 : r_xcpt_uop_ctrl_imm_sel; // @[rob.scala 660:4 rob.scala 652:18]
  wire [3:0] next_xcpt_uop_ctrl_op_fcn = T_47875 ? _GEN_28646 : r_xcpt_uop_ctrl_op_fcn; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_ctrl_fcn_dw = T_47875 ? _GEN_28647 : r_xcpt_uop_ctrl_fcn_dw; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_ctrl_rf_wen = T_47875 ? _GEN_28648 : r_xcpt_uop_ctrl_rf_wen; // @[rob.scala 660:4 rob.scala 652:18]
  wire [2:0] next_xcpt_uop_ctrl_csr_cmd = T_47875 ? _GEN_28649 : r_xcpt_uop_ctrl_csr_cmd; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_ctrl_is_load = T_47875 ? _GEN_28650 : r_xcpt_uop_ctrl_is_load; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_ctrl_is_sta = T_47875 ? _GEN_28651 : r_xcpt_uop_ctrl_is_sta; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_ctrl_is_std = T_47875 ? _GEN_28652 : r_xcpt_uop_ctrl_is_std; // @[rob.scala 660:4 rob.scala 652:18]
  wire [1:0] next_xcpt_uop_wakeup_delay = T_47875 ? _GEN_28653 : r_xcpt_uop_wakeup_delay; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_allocate_brtag = T_47875 ? _GEN_28654 : r_xcpt_uop_allocate_brtag; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_br_or_jmp = T_47875 ? _GEN_28655 : r_xcpt_uop_is_br_or_jmp; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_jump = T_47875 ? _GEN_28656 : r_xcpt_uop_is_jump; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_jal = T_47875 ? _GEN_28657 : r_xcpt_uop_is_jal; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_ret = T_47875 ? _GEN_28658 : r_xcpt_uop_is_ret; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_call = T_47875 ? _GEN_28659 : r_xcpt_uop_is_call; // @[rob.scala 660:4 rob.scala 652:18]
  wire [7:0] next_xcpt_uop_br_mask = T_47875 ? _GEN_28660 : r_xcpt_uop_br_mask; // @[rob.scala 660:4 rob.scala 652:18]
  wire [2:0] next_xcpt_uop_br_tag = T_47875 ? _GEN_28661 : r_xcpt_uop_br_tag; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_br_prediction_bpd_predict_val = T_47875 ? _GEN_28662 : r_xcpt_uop_br_prediction_bpd_predict_val; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_br_prediction_bpd_predict_taken = T_47875 ? _GEN_28663 :
    r_xcpt_uop_br_prediction_bpd_predict_taken; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_br_prediction_btb_hit = T_47875 ? _GEN_28664 : r_xcpt_uop_br_prediction_btb_hit; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_br_prediction_btb_predicted = T_47875 ? _GEN_28665 : r_xcpt_uop_br_prediction_btb_predicted; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_br_prediction_is_br_or_jalr = T_47875 ? _GEN_28666 : r_xcpt_uop_br_prediction_is_br_or_jalr; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_stat_brjmp_mispredicted = T_47875 ? _GEN_28667 : r_xcpt_uop_stat_brjmp_mispredicted; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_stat_btb_made_pred = T_47875 ? _GEN_28668 : r_xcpt_uop_stat_btb_made_pred; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_stat_btb_mispredicted = T_47875 ? _GEN_28669 : r_xcpt_uop_stat_btb_mispredicted; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_stat_bpd_made_pred = T_47875 ? _GEN_28670 : r_xcpt_uop_stat_bpd_made_pred; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_stat_bpd_mispredicted = T_47875 ? _GEN_28671 : r_xcpt_uop_stat_bpd_mispredicted; // @[rob.scala 660:4 rob.scala 652:18]
  wire [2:0] next_xcpt_uop_fetch_pc_lob = T_47875 ? _GEN_28672 : r_xcpt_uop_fetch_pc_lob; // @[rob.scala 660:4 rob.scala 652:18]
  wire [19:0] next_xcpt_uop_imm_packed = T_47875 ? _GEN_28673 : r_xcpt_uop_imm_packed; // @[rob.scala 660:4 rob.scala 652:18]
  wire [11:0] next_xcpt_uop_csr_addr = T_47875 ? _GEN_28674 : r_xcpt_uop_csr_addr; // @[rob.scala 660:4 rob.scala 652:18]
  wire [5:0] next_xcpt_uop_rob_idx = T_47875 ? _GEN_28675 : r_xcpt_uop_rob_idx; // @[rob.scala 660:4 rob.scala 652:18]
  wire [3:0] next_xcpt_uop_ldq_idx = T_47875 ? _GEN_28676 : r_xcpt_uop_ldq_idx; // @[rob.scala 660:4 rob.scala 652:18]
  wire [3:0] next_xcpt_uop_stq_idx = T_47875 ? _GEN_28677 : r_xcpt_uop_stq_idx; // @[rob.scala 660:4 rob.scala 652:18]
  wire [4:0] next_xcpt_uop_brob_idx = T_47875 ? _GEN_28678 : r_xcpt_uop_brob_idx; // @[rob.scala 660:4 rob.scala 652:18]
  wire [6:0] next_xcpt_uop_pdst = T_47875 ? _GEN_28679 : r_xcpt_uop_pdst; // @[rob.scala 660:4 rob.scala 652:18]
  wire [6:0] next_xcpt_uop_pop1 = T_47875 ? _GEN_28680 : r_xcpt_uop_pop1; // @[rob.scala 660:4 rob.scala 652:18]
  wire [6:0] next_xcpt_uop_pop2 = T_47875 ? _GEN_28681 : r_xcpt_uop_pop2; // @[rob.scala 660:4 rob.scala 652:18]
  wire [6:0] next_xcpt_uop_pop3 = T_47875 ? _GEN_28682 : r_xcpt_uop_pop3; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_prs1_busy = T_47875 ? _GEN_28683 : r_xcpt_uop_prs1_busy; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_prs2_busy = T_47875 ? _GEN_28684 : r_xcpt_uop_prs2_busy; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_prs3_busy = T_47875 ? _GEN_28685 : r_xcpt_uop_prs3_busy; // @[rob.scala 660:4 rob.scala 652:18]
  wire [6:0] next_xcpt_uop_stale_pdst = T_47875 ? _GEN_28686 : r_xcpt_uop_stale_pdst; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_exception = T_47875 ? _GEN_28687 : r_xcpt_uop_exception; // @[rob.scala 660:4 rob.scala 652:18]
  wire [63:0] next_xcpt_uop_exc_cause = T_47875 ? _GEN_28688 : r_xcpt_uop_exc_cause; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_bypassable = T_47875 ? _GEN_28689 : r_xcpt_uop_bypassable; // @[rob.scala 660:4 rob.scala 652:18]
  wire [3:0] next_xcpt_uop_mem_cmd = T_47875 ? _GEN_28690 : r_xcpt_uop_mem_cmd; // @[rob.scala 660:4 rob.scala 652:18]
  wire [2:0] next_xcpt_uop_mem_typ = T_47875 ? _GEN_28691 : r_xcpt_uop_mem_typ; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_fence = T_47875 ? _GEN_28692 : r_xcpt_uop_is_fence; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_fencei = T_47875 ? _GEN_28693 : r_xcpt_uop_is_fencei; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_store = T_47875 ? _GEN_28694 : r_xcpt_uop_is_store; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_amo = T_47875 ? _GEN_28695 : r_xcpt_uop_is_amo; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_load = T_47875 ? _GEN_28696 : r_xcpt_uop_is_load; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_is_unique = T_47875 ? _GEN_28697 : r_xcpt_uop_is_unique; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_flush_on_commit = T_47875 ? _GEN_28698 : r_xcpt_uop_flush_on_commit; // @[rob.scala 660:4 rob.scala 652:18]
  wire [5:0] next_xcpt_uop_ldst = T_47875 ? _GEN_28699 : r_xcpt_uop_ldst; // @[rob.scala 660:4 rob.scala 652:18]
  wire [5:0] next_xcpt_uop_lrs1 = T_47875 ? _GEN_28700 : r_xcpt_uop_lrs1; // @[rob.scala 660:4 rob.scala 652:18]
  wire [5:0] next_xcpt_uop_lrs2 = T_47875 ? _GEN_28701 : r_xcpt_uop_lrs2; // @[rob.scala 660:4 rob.scala 652:18]
  wire [5:0] next_xcpt_uop_lrs3 = T_47875 ? _GEN_28702 : r_xcpt_uop_lrs3; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_ldst_val = T_47875 ? _GEN_28703 : r_xcpt_uop_ldst_val; // @[rob.scala 660:4 rob.scala 652:18]
  wire [1:0] next_xcpt_uop_dst_rtype = T_47875 ? _GEN_28704 : r_xcpt_uop_dst_rtype; // @[rob.scala 660:4 rob.scala 652:18]
  wire [1:0] next_xcpt_uop_lrs1_rtype = T_47875 ? _GEN_28705 : r_xcpt_uop_lrs1_rtype; // @[rob.scala 660:4 rob.scala 652:18]
  wire [1:0] next_xcpt_uop_lrs2_rtype = T_47875 ? _GEN_28706 : r_xcpt_uop_lrs2_rtype; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_frs3_en = T_47875 ? _GEN_28707 : r_xcpt_uop_frs3_en; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_fp_val = T_47875 ? _GEN_28708 : r_xcpt_uop_fp_val; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_fp_single = T_47875 ? _GEN_28709 : r_xcpt_uop_fp_single; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_xcpt_if = T_47875 ? _GEN_28710 : r_xcpt_uop_xcpt_if; // @[rob.scala 660:4 rob.scala 652:18]
  wire  next_xcpt_uop_replay_if = T_47875 ? _GEN_28711 : r_xcpt_uop_replay_if; // @[rob.scala 660:4 rob.scala 652:18]
  wire [63:0] next_xcpt_uop_debug_wdata = T_47875 ? _GEN_28712 : r_xcpt_uop_debug_wdata; // @[rob.scala 660:4 rob.scala 652:18]
  wire [31:0] next_xcpt_uop_debug_events_fetch_seq = T_47875 ? _GEN_28713 : r_xcpt_uop_debug_events_fetch_seq; // @[rob.scala 660:4 rob.scala 652:18]
  wire [7:0] T_48086 = next_xcpt_uop_br_mask & T_29465; // @[util.scala 32:45]
  wire [7:0] T_48087 = io_brinfo_valid ? T_48086 : next_xcpt_uop_br_mask; // @[util.scala 32:17]
  wire [7:0] T_48089 = io_brinfo_mask & next_xcpt_uop_br_mask; // @[util.scala 45:52]
  wire  T_48091 = T_48089 != 8'h0; // @[util.scala 45:60]
  wire  T_48092 = T_29369 & T_48091; // @[util.scala 23:33]
  wire  T_48093 = io_flush_pipeline | T_48092; // @[rob.scala 688:28]
  wire  T_48096 = ~io_cxcpt_valid; // @[rob.scala 693:34]
  wire  T_48097 = T_47568 & T_48096; // @[rob.scala 693:31]
  wire  T_48100 = T_48097 & T_47975; // @[rob.scala 693:50]
  wire  T_48102 = ~T_48100; // @[rob.scala 693:12]
  wire  T_48103 = T_48102 | reset; // @[rob.scala 693:11]
  wire  T_48105 = ~T_48103; // @[rob.scala 693:11]
  wire  T_48106 = io_empty & r_xcpt_val; // @[rob.scala 696:23]
  wire  T_48108 = ~T_48106; // @[rob.scala 696:12]
  wire  T_48109 = T_48108 | reset; // @[rob.scala 696:11]
  wire  T_48111 = ~T_48109; // @[rob.scala 696:11]
  wire [5:0] T_48113 = {{1'd0}, r_xcpt_uop_rob_idx[5:1]}; // @[rob.scala 222:27]
  wire [5:0] _GEN_28925 = {{1'd0}, rob_head}; // @[rob.scala 699:69]
  wire  T_48114 = T_48113 != _GEN_28925; // @[rob.scala 699:69]
  wire  T_48115 = will_throw_exception & T_48114; // @[rob.scala 699:35]
  wire  T_48117 = ~T_48115; // @[rob.scala 699:12]
  wire  T_48118 = T_48117 | reset; // @[rob.scala 699:11]
  wire  T_48120 = ~T_48118; // @[rob.scala 699:11]
  wire  T_48136 = rob_head == 5'h17; // @[util.scala 75:28]
  wire [4:0] T_48140 = rob_head + 5'h1; // @[util.scala 76:35]
  wire  T_48143 = rob_tail != rob_head; // @[rob.scala 726:47]
  wire  T_48144 = T_29097 & T_48143; // @[rob.scala 726:35]
  wire  T_48146 = rob_tail == 5'h0; // @[util.scala 91:28]
  wire [4:0] T_48150 = rob_tail - 5'h1; // @[util.scala 92:39]
  wire [4:0] T_48151 = T_48146 ? 5'h17 : T_48150; // @[util.scala 92:13]
  wire [4:0] _GEN_28797 = T_48144 ? T_48151 : rob_tail; // @[rob.scala 727:4 rob.scala 728:16]
  wire  T_48154 = ~T_48144; // @[rob.scala 727:4]
  wire  T_48155 = T_48154 & T_29369; // @[rob.scala 731:4]
  wire  T_48159 = T_28625 == 6'h17; // @[util.scala 75:28]
  wire [5:0] T_48163 = T_28625 + 6'h1; // @[util.scala 76:35]
  wire [5:0] T_48164 = T_48159 ? 6'h0 : T_48163; // @[util.scala 76:13]
  wire [5:0] _GEN_28798 = T_48155 ? T_48164 : {{1'd0}, _GEN_28797}; // @[rob.scala 731:4 rob.scala 732:16]
  wire  T_48167 = T_23625 != 2'h0; // @[rob.scala 734:36]
  wire  T_48169 = ~io_dis_partial_stall; // @[rob.scala 734:51]
  wire  T_48170 = T_48167 & T_48169; // @[rob.scala 734:48]
  wire  T_48175 = ~(T_48144 | T_29369);
  wire  T_48176 = T_48175 & T_48170; // @[rob.scala 735:4]
  wire  T_48178 = rob_tail == 5'h17; // @[util.scala 75:28]
  wire [4:0] T_48182 = rob_tail + 5'h1; // @[util.scala 76:35]
  wire [4:0] T_48183 = T_48178 ? 5'h0 : T_48182; // @[util.scala 76:13]
  wire [5:0] _GEN_28799 = T_48176 ? {{1'd0}, T_48183} : _GEN_28798; // @[rob.scala 735:4 rob.scala 736:16]
  wire  full = T_48183 == rob_head; // @[rob.scala 757:47]
  wire  T_48194 = T_48125 == 2'h0; // @[rob.scala 759:65]
  wire  T_48196 = rob_state == 2'h1; // @[rob.scala 764:27]
  wire  T_48198 = ~full; // @[rob.scala 764:44]
  wire  T_48200 = 2'h0 == rob_state; // @[Conditional.scala 24:42]
  wire [1:0] _GEN_28800 = T_48200 ? 2'h1 : rob_state; // @[Conditional.scala 24:73 rob.scala 777:23]
  wire  T_48201 = 2'h1 == rob_state; // @[Conditional.scala 24:42]
  wire [1:0] _GEN_28801 = T_47568 ? 2'h2 : _GEN_28800; // @[rob.scala 782:13 rob.scala 783:26]
  wire  T_48203 = ~T_47568; // @[rob.scala 782:13]
  wire [1:0] _GEN_28802 = T_23670 ? 2'h3 : _GEN_28801; // @[rob.scala 790:19 rob.scala 791:32]
  wire [1:0] _GEN_28803 = T_23671 ? 2'h3 : _GEN_28802; // @[rob.scala 790:19 rob.scala 791:32]
  wire [1:0] _GEN_28804 = T_48203 ? _GEN_28803 : _GEN_28801; // @[rob.scala 786:13]
  wire [1:0] _GEN_28805 = T_48201 ? _GEN_28804 : _GEN_28800; // @[Conditional.scala 24:73]
  wire  T_48206 = 2'h2 == rob_state; // @[Conditional.scala 24:42]
  wire [1:0] _GEN_28806 = io_empty ? 2'h1 : _GEN_28805; // @[rob.scala 799:13 rob.scala 800:26]
  wire [1:0] _GEN_28807 = T_48206 ? _GEN_28806 : _GEN_28805; // @[Conditional.scala 24:73]
  wire  T_48207 = 2'h3 == rob_state; // @[Conditional.scala 24:42]
  wire  T_48210 = T_48203 & io_empty; // @[rob.scala 810:13]
  wire  T_48216 = T_48125[0]; // @[OneHot.scala 35:40]
  wire  T_48220 = T_48216 ? 1'h0 : 1'h1; // @[Mux.scala 31:69]
  wire [7:0] T_48223 = r_xcpt_val ? 8'h45 : 8'h2d; // @[rob.scala 946:18]
  wire  T_48225 = ~reset; // @[rob.scala 945:13]
  wire  T_48228 = rob_head == 5'h0; // @[rob.scala 970:26]
  wire  T_48231 = T_48228 & T_48146; // @[rob.scala 970:40]
  wire [7:0] T_48240 = T_48146 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48241 = T_48228 ? 8'h48 : T_48240; // @[rob.scala 971:18]
  wire [7:0] T_48242 = T_48231 ? 8'h42 : T_48241; // @[rob.scala 970:18]
  wire [7:0] T_48252 = T_23706_0 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48255 = T_35634_0 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_0_busy = T_23710_T_32866_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48258 = debug_entry_0_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_1_busy = T_35638_T_44794_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48261 = debug_entry_1_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_0_uop_pc = T_32976[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48262 = debug_entry_0_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_1_uop_pc = T_44904[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48263 = debug_entry_1_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_0_exception = T_28311_T_32978_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48274 = debug_entry_0_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_1_exception = T_40239_T_44906_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48277 = debug_entry_1_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48280 = T_26182_0_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48282 = T_26182_0_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48284 = T_26182_0_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48286 = T_26182_0_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48289 = T_48286 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48290 = T_48284 ? 8'h66 : T_48289; // @[rob.scala 1050:21]
  wire [7:0] T_48291 = T_48282 ? 8'h43 : T_48290; // @[rob.scala 1049:21]
  wire [7:0] T_48292 = T_48280 ? 8'h58 : T_48291; // @[rob.scala 1048:21]
  wire  T_48295 = T_38110_0_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48297 = T_38110_0_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48299 = T_38110_0_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48301 = T_38110_0_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48304 = T_48301 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48305 = T_48299 ? 8'h66 : T_48304; // @[rob.scala 1050:21]
  wire [7:0] T_48306 = T_48297 ? 8'h43 : T_48305; // @[rob.scala 1049:21]
  wire [7:0] T_48307 = T_48295 ? 8'h58 : T_48306; // @[rob.scala 1048:21]
  wire  T_48314 = rob_head == 5'h1; // @[rob.scala 970:26]
  wire  T_48316 = rob_tail == 5'h1; // @[rob.scala 970:50]
  wire  T_48317 = T_48314 & T_48316; // @[rob.scala 970:40]
  wire [7:0] T_48326 = T_48316 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48327 = T_48314 ? 8'h48 : T_48326; // @[rob.scala 971:18]
  wire [7:0] T_48328 = T_48317 ? 8'h42 : T_48327; // @[rob.scala 970:18]
  wire [7:0] T_48338 = T_23706_1 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48341 = T_35634_1 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_2_busy = T_23710_T_32980_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48344 = debug_entry_2_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_3_busy = T_35638_T_44908_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48347 = debug_entry_3_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_2_uop_pc = T_33090[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48348 = debug_entry_2_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_3_uop_pc = T_45018[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48349 = debug_entry_3_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_2_exception = T_28311_T_33092_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48360 = debug_entry_2_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_3_exception = T_40239_T_45020_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48363 = debug_entry_3_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48366 = T_26182_1_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48368 = T_26182_1_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48370 = T_26182_1_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48372 = T_26182_1_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48375 = T_48372 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48376 = T_48370 ? 8'h66 : T_48375; // @[rob.scala 1050:21]
  wire [7:0] T_48377 = T_48368 ? 8'h43 : T_48376; // @[rob.scala 1049:21]
  wire [7:0] T_48378 = T_48366 ? 8'h58 : T_48377; // @[rob.scala 1048:21]
  wire  T_48381 = T_38110_1_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48383 = T_38110_1_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48385 = T_38110_1_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48387 = T_38110_1_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48390 = T_48387 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48391 = T_48385 ? 8'h66 : T_48390; // @[rob.scala 1050:21]
  wire [7:0] T_48392 = T_48383 ? 8'h43 : T_48391; // @[rob.scala 1049:21]
  wire [7:0] T_48393 = T_48381 ? 8'h58 : T_48392; // @[rob.scala 1048:21]
  wire  T_48400 = rob_head == 5'h2; // @[rob.scala 970:26]
  wire  T_48402 = rob_tail == 5'h2; // @[rob.scala 970:50]
  wire  T_48403 = T_48400 & T_48402; // @[rob.scala 970:40]
  wire [7:0] T_48412 = T_48402 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48413 = T_48400 ? 8'h48 : T_48412; // @[rob.scala 971:18]
  wire [7:0] T_48414 = T_48403 ? 8'h42 : T_48413; // @[rob.scala 970:18]
  wire [7:0] T_48424 = T_23706_2 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48427 = T_35634_2 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_4_busy = T_23710_T_33094_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48430 = debug_entry_4_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_5_busy = T_35638_T_45022_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48433 = debug_entry_5_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_4_uop_pc = T_33204[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48434 = debug_entry_4_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_5_uop_pc = T_45132[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48435 = debug_entry_5_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_4_exception = T_28311_T_33206_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48446 = debug_entry_4_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_5_exception = T_40239_T_45134_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48449 = debug_entry_5_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48452 = T_26182_2_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48454 = T_26182_2_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48456 = T_26182_2_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48458 = T_26182_2_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48461 = T_48458 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48462 = T_48456 ? 8'h66 : T_48461; // @[rob.scala 1050:21]
  wire [7:0] T_48463 = T_48454 ? 8'h43 : T_48462; // @[rob.scala 1049:21]
  wire [7:0] T_48464 = T_48452 ? 8'h58 : T_48463; // @[rob.scala 1048:21]
  wire  T_48467 = T_38110_2_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48469 = T_38110_2_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48471 = T_38110_2_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48473 = T_38110_2_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48476 = T_48473 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48477 = T_48471 ? 8'h66 : T_48476; // @[rob.scala 1050:21]
  wire [7:0] T_48478 = T_48469 ? 8'h43 : T_48477; // @[rob.scala 1049:21]
  wire [7:0] T_48479 = T_48467 ? 8'h58 : T_48478; // @[rob.scala 1048:21]
  wire  T_48486 = rob_head == 5'h3; // @[rob.scala 970:26]
  wire  T_48488 = rob_tail == 5'h3; // @[rob.scala 970:50]
  wire  T_48489 = T_48486 & T_48488; // @[rob.scala 970:40]
  wire [7:0] T_48498 = T_48488 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48499 = T_48486 ? 8'h48 : T_48498; // @[rob.scala 971:18]
  wire [7:0] T_48500 = T_48489 ? 8'h42 : T_48499; // @[rob.scala 970:18]
  wire [7:0] T_48510 = T_23706_3 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48513 = T_35634_3 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_6_busy = T_23710_T_33208_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48516 = debug_entry_6_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_7_busy = T_35638_T_45136_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48519 = debug_entry_7_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_6_uop_pc = T_33318[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48520 = debug_entry_6_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_7_uop_pc = T_45246[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48521 = debug_entry_7_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_6_exception = T_28311_T_33320_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48532 = debug_entry_6_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_7_exception = T_40239_T_45248_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48535 = debug_entry_7_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48538 = T_26182_3_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48540 = T_26182_3_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48542 = T_26182_3_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48544 = T_26182_3_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48547 = T_48544 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48548 = T_48542 ? 8'h66 : T_48547; // @[rob.scala 1050:21]
  wire [7:0] T_48549 = T_48540 ? 8'h43 : T_48548; // @[rob.scala 1049:21]
  wire [7:0] T_48550 = T_48538 ? 8'h58 : T_48549; // @[rob.scala 1048:21]
  wire  T_48553 = T_38110_3_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48555 = T_38110_3_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48557 = T_38110_3_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48559 = T_38110_3_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48562 = T_48559 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48563 = T_48557 ? 8'h66 : T_48562; // @[rob.scala 1050:21]
  wire [7:0] T_48564 = T_48555 ? 8'h43 : T_48563; // @[rob.scala 1049:21]
  wire [7:0] T_48565 = T_48553 ? 8'h58 : T_48564; // @[rob.scala 1048:21]
  wire  T_48572 = rob_head == 5'h4; // @[rob.scala 970:26]
  wire  T_48574 = rob_tail == 5'h4; // @[rob.scala 970:50]
  wire  T_48575 = T_48572 & T_48574; // @[rob.scala 970:40]
  wire [7:0] T_48584 = T_48574 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48585 = T_48572 ? 8'h48 : T_48584; // @[rob.scala 971:18]
  wire [7:0] T_48586 = T_48575 ? 8'h42 : T_48585; // @[rob.scala 970:18]
  wire [7:0] T_48596 = T_23706_4 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48599 = T_35634_4 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_8_busy = T_23710_T_33322_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48602 = debug_entry_8_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_9_busy = T_35638_T_45250_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48605 = debug_entry_9_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_8_uop_pc = T_33432[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48606 = debug_entry_8_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_9_uop_pc = T_45360[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48607 = debug_entry_9_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_8_exception = T_28311_T_33434_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48618 = debug_entry_8_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_9_exception = T_40239_T_45362_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48621 = debug_entry_9_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48624 = T_26182_4_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48626 = T_26182_4_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48628 = T_26182_4_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48630 = T_26182_4_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48633 = T_48630 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48634 = T_48628 ? 8'h66 : T_48633; // @[rob.scala 1050:21]
  wire [7:0] T_48635 = T_48626 ? 8'h43 : T_48634; // @[rob.scala 1049:21]
  wire [7:0] T_48636 = T_48624 ? 8'h58 : T_48635; // @[rob.scala 1048:21]
  wire  T_48639 = T_38110_4_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48641 = T_38110_4_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48643 = T_38110_4_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48645 = T_38110_4_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48648 = T_48645 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48649 = T_48643 ? 8'h66 : T_48648; // @[rob.scala 1050:21]
  wire [7:0] T_48650 = T_48641 ? 8'h43 : T_48649; // @[rob.scala 1049:21]
  wire [7:0] T_48651 = T_48639 ? 8'h58 : T_48650; // @[rob.scala 1048:21]
  wire  T_48658 = rob_head == 5'h5; // @[rob.scala 970:26]
  wire  T_48660 = rob_tail == 5'h5; // @[rob.scala 970:50]
  wire  T_48661 = T_48658 & T_48660; // @[rob.scala 970:40]
  wire [7:0] T_48670 = T_48660 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48671 = T_48658 ? 8'h48 : T_48670; // @[rob.scala 971:18]
  wire [7:0] T_48672 = T_48661 ? 8'h42 : T_48671; // @[rob.scala 970:18]
  wire [7:0] T_48682 = T_23706_5 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48685 = T_35634_5 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_10_busy = T_23710_T_33436_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48688 = debug_entry_10_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_11_busy = T_35638_T_45364_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48691 = debug_entry_11_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_10_uop_pc = T_33546[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48692 = debug_entry_10_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_11_uop_pc = T_45474[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48693 = debug_entry_11_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_10_exception = T_28311_T_33548_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48704 = debug_entry_10_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_11_exception = T_40239_T_45476_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48707 = debug_entry_11_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48710 = T_26182_5_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48712 = T_26182_5_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48714 = T_26182_5_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48716 = T_26182_5_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48719 = T_48716 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48720 = T_48714 ? 8'h66 : T_48719; // @[rob.scala 1050:21]
  wire [7:0] T_48721 = T_48712 ? 8'h43 : T_48720; // @[rob.scala 1049:21]
  wire [7:0] T_48722 = T_48710 ? 8'h58 : T_48721; // @[rob.scala 1048:21]
  wire  T_48725 = T_38110_5_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48727 = T_38110_5_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48729 = T_38110_5_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48731 = T_38110_5_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48734 = T_48731 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48735 = T_48729 ? 8'h66 : T_48734; // @[rob.scala 1050:21]
  wire [7:0] T_48736 = T_48727 ? 8'h43 : T_48735; // @[rob.scala 1049:21]
  wire [7:0] T_48737 = T_48725 ? 8'h58 : T_48736; // @[rob.scala 1048:21]
  wire  T_48744 = rob_head == 5'h6; // @[rob.scala 970:26]
  wire  T_48746 = rob_tail == 5'h6; // @[rob.scala 970:50]
  wire  T_48747 = T_48744 & T_48746; // @[rob.scala 970:40]
  wire [7:0] T_48756 = T_48746 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48757 = T_48744 ? 8'h48 : T_48756; // @[rob.scala 971:18]
  wire [7:0] T_48758 = T_48747 ? 8'h42 : T_48757; // @[rob.scala 970:18]
  wire [7:0] T_48768 = T_23706_6 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48771 = T_35634_6 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_12_busy = T_23710_T_33550_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48774 = debug_entry_12_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_13_busy = T_35638_T_45478_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48777 = debug_entry_13_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_12_uop_pc = T_33660[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48778 = debug_entry_12_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_13_uop_pc = T_45588[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48779 = debug_entry_13_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_12_exception = T_28311_T_33662_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48790 = debug_entry_12_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_13_exception = T_40239_T_45590_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48793 = debug_entry_13_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48796 = T_26182_6_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48798 = T_26182_6_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48800 = T_26182_6_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48802 = T_26182_6_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48805 = T_48802 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48806 = T_48800 ? 8'h66 : T_48805; // @[rob.scala 1050:21]
  wire [7:0] T_48807 = T_48798 ? 8'h43 : T_48806; // @[rob.scala 1049:21]
  wire [7:0] T_48808 = T_48796 ? 8'h58 : T_48807; // @[rob.scala 1048:21]
  wire  T_48811 = T_38110_6_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48813 = T_38110_6_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48815 = T_38110_6_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48817 = T_38110_6_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48820 = T_48817 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48821 = T_48815 ? 8'h66 : T_48820; // @[rob.scala 1050:21]
  wire [7:0] T_48822 = T_48813 ? 8'h43 : T_48821; // @[rob.scala 1049:21]
  wire [7:0] T_48823 = T_48811 ? 8'h58 : T_48822; // @[rob.scala 1048:21]
  wire  T_48830 = rob_head == 5'h7; // @[rob.scala 970:26]
  wire  T_48832 = rob_tail == 5'h7; // @[rob.scala 970:50]
  wire  T_48833 = T_48830 & T_48832; // @[rob.scala 970:40]
  wire [7:0] T_48842 = T_48832 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48843 = T_48830 ? 8'h48 : T_48842; // @[rob.scala 971:18]
  wire [7:0] T_48844 = T_48833 ? 8'h42 : T_48843; // @[rob.scala 970:18]
  wire [7:0] T_48854 = T_23706_7 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48857 = T_35634_7 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_14_busy = T_23710_T_33664_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48860 = debug_entry_14_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_15_busy = T_35638_T_45592_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48863 = debug_entry_15_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_14_uop_pc = T_33774[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48864 = debug_entry_14_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_15_uop_pc = T_45702[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48865 = debug_entry_15_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_14_exception = T_28311_T_33776_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48876 = debug_entry_14_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_15_exception = T_40239_T_45704_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48879 = debug_entry_15_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48882 = T_26182_7_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48884 = T_26182_7_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48886 = T_26182_7_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48888 = T_26182_7_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48891 = T_48888 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48892 = T_48886 ? 8'h66 : T_48891; // @[rob.scala 1050:21]
  wire [7:0] T_48893 = T_48884 ? 8'h43 : T_48892; // @[rob.scala 1049:21]
  wire [7:0] T_48894 = T_48882 ? 8'h58 : T_48893; // @[rob.scala 1048:21]
  wire  T_48897 = T_38110_7_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48899 = T_38110_7_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48901 = T_38110_7_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48903 = T_38110_7_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48906 = T_48903 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48907 = T_48901 ? 8'h66 : T_48906; // @[rob.scala 1050:21]
  wire [7:0] T_48908 = T_48899 ? 8'h43 : T_48907; // @[rob.scala 1049:21]
  wire [7:0] T_48909 = T_48897 ? 8'h58 : T_48908; // @[rob.scala 1048:21]
  wire  T_48916 = rob_head == 5'h8; // @[rob.scala 970:26]
  wire  T_48918 = rob_tail == 5'h8; // @[rob.scala 970:50]
  wire  T_48919 = T_48916 & T_48918; // @[rob.scala 970:40]
  wire [7:0] T_48928 = T_48918 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_48929 = T_48916 ? 8'h48 : T_48928; // @[rob.scala 971:18]
  wire [7:0] T_48930 = T_48919 ? 8'h42 : T_48929; // @[rob.scala 970:18]
  wire [7:0] T_48940 = T_23706_8 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_48943 = T_35634_8 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_16_busy = T_23710_T_33778_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48946 = debug_entry_16_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_17_busy = T_35638_T_45706_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_48949 = debug_entry_17_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_16_uop_pc = T_33888[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_48950 = debug_entry_16_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_17_uop_pc = T_45816[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_48951 = debug_entry_17_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_16_exception = T_28311_T_33890_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48962 = debug_entry_16_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_17_exception = T_40239_T_45818_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_48965 = debug_entry_17_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_48968 = T_26182_8_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48970 = T_26182_8_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48972 = T_26182_8_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48974 = T_26182_8_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48977 = T_48974 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48978 = T_48972 ? 8'h66 : T_48977; // @[rob.scala 1050:21]
  wire [7:0] T_48979 = T_48970 ? 8'h43 : T_48978; // @[rob.scala 1049:21]
  wire [7:0] T_48980 = T_48968 ? 8'h58 : T_48979; // @[rob.scala 1048:21]
  wire  T_48983 = T_38110_8_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_48985 = T_38110_8_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_48987 = T_38110_8_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_48989 = T_38110_8_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_48992 = T_48989 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_48993 = T_48987 ? 8'h66 : T_48992; // @[rob.scala 1050:21]
  wire [7:0] T_48994 = T_48985 ? 8'h43 : T_48993; // @[rob.scala 1049:21]
  wire [7:0] T_48995 = T_48983 ? 8'h58 : T_48994; // @[rob.scala 1048:21]
  wire  T_49002 = rob_head == 5'h9; // @[rob.scala 970:26]
  wire  T_49004 = rob_tail == 5'h9; // @[rob.scala 970:50]
  wire  T_49005 = T_49002 & T_49004; // @[rob.scala 970:40]
  wire [7:0] T_49014 = T_49004 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49015 = T_49002 ? 8'h48 : T_49014; // @[rob.scala 971:18]
  wire [7:0] T_49016 = T_49005 ? 8'h42 : T_49015; // @[rob.scala 970:18]
  wire [7:0] T_49026 = T_23706_9 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49029 = T_35634_9 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_18_busy = T_23710_T_33892_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49032 = debug_entry_18_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_19_busy = T_35638_T_45820_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49035 = debug_entry_19_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_18_uop_pc = T_34002[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49036 = debug_entry_18_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_19_uop_pc = T_45930[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49037 = debug_entry_19_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_18_exception = T_28311_T_34004_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49048 = debug_entry_18_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_19_exception = T_40239_T_45932_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49051 = debug_entry_19_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49054 = T_26182_9_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49056 = T_26182_9_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49058 = T_26182_9_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49060 = T_26182_9_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49063 = T_49060 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49064 = T_49058 ? 8'h66 : T_49063; // @[rob.scala 1050:21]
  wire [7:0] T_49065 = T_49056 ? 8'h43 : T_49064; // @[rob.scala 1049:21]
  wire [7:0] T_49066 = T_49054 ? 8'h58 : T_49065; // @[rob.scala 1048:21]
  wire  T_49069 = T_38110_9_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49071 = T_38110_9_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49073 = T_38110_9_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49075 = T_38110_9_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49078 = T_49075 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49079 = T_49073 ? 8'h66 : T_49078; // @[rob.scala 1050:21]
  wire [7:0] T_49080 = T_49071 ? 8'h43 : T_49079; // @[rob.scala 1049:21]
  wire [7:0] T_49081 = T_49069 ? 8'h58 : T_49080; // @[rob.scala 1048:21]
  wire  T_49088 = rob_head == 5'ha; // @[rob.scala 970:26]
  wire  T_49090 = rob_tail == 5'ha; // @[rob.scala 970:50]
  wire  T_49091 = T_49088 & T_49090; // @[rob.scala 970:40]
  wire [7:0] T_49100 = T_49090 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49101 = T_49088 ? 8'h48 : T_49100; // @[rob.scala 971:18]
  wire [7:0] T_49102 = T_49091 ? 8'h42 : T_49101; // @[rob.scala 970:18]
  wire [7:0] T_49112 = T_23706_10 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49115 = T_35634_10 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_20_busy = T_23710_T_34006_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49118 = debug_entry_20_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_21_busy = T_35638_T_45934_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49121 = debug_entry_21_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_20_uop_pc = T_34116[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49122 = debug_entry_20_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_21_uop_pc = T_46044[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49123 = debug_entry_21_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_20_exception = T_28311_T_34118_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49134 = debug_entry_20_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_21_exception = T_40239_T_46046_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49137 = debug_entry_21_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49140 = T_26182_10_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49142 = T_26182_10_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49144 = T_26182_10_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49146 = T_26182_10_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49149 = T_49146 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49150 = T_49144 ? 8'h66 : T_49149; // @[rob.scala 1050:21]
  wire [7:0] T_49151 = T_49142 ? 8'h43 : T_49150; // @[rob.scala 1049:21]
  wire [7:0] T_49152 = T_49140 ? 8'h58 : T_49151; // @[rob.scala 1048:21]
  wire  T_49155 = T_38110_10_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49157 = T_38110_10_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49159 = T_38110_10_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49161 = T_38110_10_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49164 = T_49161 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49165 = T_49159 ? 8'h66 : T_49164; // @[rob.scala 1050:21]
  wire [7:0] T_49166 = T_49157 ? 8'h43 : T_49165; // @[rob.scala 1049:21]
  wire [7:0] T_49167 = T_49155 ? 8'h58 : T_49166; // @[rob.scala 1048:21]
  wire  T_49174 = rob_head == 5'hb; // @[rob.scala 970:26]
  wire  T_49176 = rob_tail == 5'hb; // @[rob.scala 970:50]
  wire  T_49177 = T_49174 & T_49176; // @[rob.scala 970:40]
  wire [7:0] T_49186 = T_49176 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49187 = T_49174 ? 8'h48 : T_49186; // @[rob.scala 971:18]
  wire [7:0] T_49188 = T_49177 ? 8'h42 : T_49187; // @[rob.scala 970:18]
  wire [7:0] T_49198 = T_23706_11 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49201 = T_35634_11 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_22_busy = T_23710_T_34120_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49204 = debug_entry_22_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_23_busy = T_35638_T_46048_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49207 = debug_entry_23_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_22_uop_pc = T_34230[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49208 = debug_entry_22_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_23_uop_pc = T_46158[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49209 = debug_entry_23_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_22_exception = T_28311_T_34232_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49220 = debug_entry_22_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_23_exception = T_40239_T_46160_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49223 = debug_entry_23_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49226 = T_26182_11_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49228 = T_26182_11_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49230 = T_26182_11_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49232 = T_26182_11_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49235 = T_49232 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49236 = T_49230 ? 8'h66 : T_49235; // @[rob.scala 1050:21]
  wire [7:0] T_49237 = T_49228 ? 8'h43 : T_49236; // @[rob.scala 1049:21]
  wire [7:0] T_49238 = T_49226 ? 8'h58 : T_49237; // @[rob.scala 1048:21]
  wire  T_49241 = T_38110_11_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49243 = T_38110_11_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49245 = T_38110_11_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49247 = T_38110_11_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49250 = T_49247 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49251 = T_49245 ? 8'h66 : T_49250; // @[rob.scala 1050:21]
  wire [7:0] T_49252 = T_49243 ? 8'h43 : T_49251; // @[rob.scala 1049:21]
  wire [7:0] T_49253 = T_49241 ? 8'h58 : T_49252; // @[rob.scala 1048:21]
  wire  T_49260 = rob_head == 5'hc; // @[rob.scala 970:26]
  wire  T_49262 = rob_tail == 5'hc; // @[rob.scala 970:50]
  wire  T_49263 = T_49260 & T_49262; // @[rob.scala 970:40]
  wire [7:0] T_49272 = T_49262 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49273 = T_49260 ? 8'h48 : T_49272; // @[rob.scala 971:18]
  wire [7:0] T_49274 = T_49263 ? 8'h42 : T_49273; // @[rob.scala 970:18]
  wire [7:0] T_49284 = T_23706_12 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49287 = T_35634_12 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_24_busy = T_23710_T_34234_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49290 = debug_entry_24_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_25_busy = T_35638_T_46162_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49293 = debug_entry_25_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_24_uop_pc = T_34344[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49294 = debug_entry_24_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_25_uop_pc = T_46272[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49295 = debug_entry_25_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_24_exception = T_28311_T_34346_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49306 = debug_entry_24_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_25_exception = T_40239_T_46274_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49309 = debug_entry_25_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49312 = T_26182_12_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49314 = T_26182_12_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49316 = T_26182_12_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49318 = T_26182_12_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49321 = T_49318 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49322 = T_49316 ? 8'h66 : T_49321; // @[rob.scala 1050:21]
  wire [7:0] T_49323 = T_49314 ? 8'h43 : T_49322; // @[rob.scala 1049:21]
  wire [7:0] T_49324 = T_49312 ? 8'h58 : T_49323; // @[rob.scala 1048:21]
  wire  T_49327 = T_38110_12_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49329 = T_38110_12_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49331 = T_38110_12_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49333 = T_38110_12_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49336 = T_49333 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49337 = T_49331 ? 8'h66 : T_49336; // @[rob.scala 1050:21]
  wire [7:0] T_49338 = T_49329 ? 8'h43 : T_49337; // @[rob.scala 1049:21]
  wire [7:0] T_49339 = T_49327 ? 8'h58 : T_49338; // @[rob.scala 1048:21]
  wire  T_49346 = rob_head == 5'hd; // @[rob.scala 970:26]
  wire  T_49348 = rob_tail == 5'hd; // @[rob.scala 970:50]
  wire  T_49349 = T_49346 & T_49348; // @[rob.scala 970:40]
  wire [7:0] T_49358 = T_49348 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49359 = T_49346 ? 8'h48 : T_49358; // @[rob.scala 971:18]
  wire [7:0] T_49360 = T_49349 ? 8'h42 : T_49359; // @[rob.scala 970:18]
  wire [7:0] T_49370 = T_23706_13 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49373 = T_35634_13 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_26_busy = T_23710_T_34348_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49376 = debug_entry_26_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_27_busy = T_35638_T_46276_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49379 = debug_entry_27_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_26_uop_pc = T_34458[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49380 = debug_entry_26_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_27_uop_pc = T_46386[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49381 = debug_entry_27_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_26_exception = T_28311_T_34460_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49392 = debug_entry_26_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_27_exception = T_40239_T_46388_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49395 = debug_entry_27_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49398 = T_26182_13_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49400 = T_26182_13_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49402 = T_26182_13_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49404 = T_26182_13_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49407 = T_49404 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49408 = T_49402 ? 8'h66 : T_49407; // @[rob.scala 1050:21]
  wire [7:0] T_49409 = T_49400 ? 8'h43 : T_49408; // @[rob.scala 1049:21]
  wire [7:0] T_49410 = T_49398 ? 8'h58 : T_49409; // @[rob.scala 1048:21]
  wire  T_49413 = T_38110_13_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49415 = T_38110_13_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49417 = T_38110_13_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49419 = T_38110_13_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49422 = T_49419 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49423 = T_49417 ? 8'h66 : T_49422; // @[rob.scala 1050:21]
  wire [7:0] T_49424 = T_49415 ? 8'h43 : T_49423; // @[rob.scala 1049:21]
  wire [7:0] T_49425 = T_49413 ? 8'h58 : T_49424; // @[rob.scala 1048:21]
  wire  T_49432 = rob_head == 5'he; // @[rob.scala 970:26]
  wire  T_49434 = rob_tail == 5'he; // @[rob.scala 970:50]
  wire  T_49435 = T_49432 & T_49434; // @[rob.scala 970:40]
  wire [7:0] T_49444 = T_49434 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49445 = T_49432 ? 8'h48 : T_49444; // @[rob.scala 971:18]
  wire [7:0] T_49446 = T_49435 ? 8'h42 : T_49445; // @[rob.scala 970:18]
  wire [7:0] T_49456 = T_23706_14 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49459 = T_35634_14 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_28_busy = T_23710_T_34462_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49462 = debug_entry_28_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_29_busy = T_35638_T_46390_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49465 = debug_entry_29_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_28_uop_pc = T_34572[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49466 = debug_entry_28_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_29_uop_pc = T_46500[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49467 = debug_entry_29_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_28_exception = T_28311_T_34574_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49478 = debug_entry_28_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_29_exception = T_40239_T_46502_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49481 = debug_entry_29_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49484 = T_26182_14_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49486 = T_26182_14_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49488 = T_26182_14_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49490 = T_26182_14_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49493 = T_49490 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49494 = T_49488 ? 8'h66 : T_49493; // @[rob.scala 1050:21]
  wire [7:0] T_49495 = T_49486 ? 8'h43 : T_49494; // @[rob.scala 1049:21]
  wire [7:0] T_49496 = T_49484 ? 8'h58 : T_49495; // @[rob.scala 1048:21]
  wire  T_49499 = T_38110_14_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49501 = T_38110_14_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49503 = T_38110_14_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49505 = T_38110_14_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49508 = T_49505 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49509 = T_49503 ? 8'h66 : T_49508; // @[rob.scala 1050:21]
  wire [7:0] T_49510 = T_49501 ? 8'h43 : T_49509; // @[rob.scala 1049:21]
  wire [7:0] T_49511 = T_49499 ? 8'h58 : T_49510; // @[rob.scala 1048:21]
  wire  T_49518 = rob_head == 5'hf; // @[rob.scala 970:26]
  wire  T_49520 = rob_tail == 5'hf; // @[rob.scala 970:50]
  wire  T_49521 = T_49518 & T_49520; // @[rob.scala 970:40]
  wire [7:0] T_49530 = T_49520 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49531 = T_49518 ? 8'h48 : T_49530; // @[rob.scala 971:18]
  wire [7:0] T_49532 = T_49521 ? 8'h42 : T_49531; // @[rob.scala 970:18]
  wire [7:0] T_49542 = T_23706_15 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49545 = T_35634_15 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_30_busy = T_23710_T_34576_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49548 = debug_entry_30_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_31_busy = T_35638_T_46504_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49551 = debug_entry_31_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_30_uop_pc = T_34686[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49552 = debug_entry_30_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_31_uop_pc = T_46614[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49553 = debug_entry_31_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_30_exception = T_28311_T_34688_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49564 = debug_entry_30_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_31_exception = T_40239_T_46616_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49567 = debug_entry_31_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49570 = T_26182_15_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49572 = T_26182_15_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49574 = T_26182_15_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49576 = T_26182_15_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49579 = T_49576 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49580 = T_49574 ? 8'h66 : T_49579; // @[rob.scala 1050:21]
  wire [7:0] T_49581 = T_49572 ? 8'h43 : T_49580; // @[rob.scala 1049:21]
  wire [7:0] T_49582 = T_49570 ? 8'h58 : T_49581; // @[rob.scala 1048:21]
  wire  T_49585 = T_38110_15_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49587 = T_38110_15_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49589 = T_38110_15_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49591 = T_38110_15_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49594 = T_49591 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49595 = T_49589 ? 8'h66 : T_49594; // @[rob.scala 1050:21]
  wire [7:0] T_49596 = T_49587 ? 8'h43 : T_49595; // @[rob.scala 1049:21]
  wire [7:0] T_49597 = T_49585 ? 8'h58 : T_49596; // @[rob.scala 1048:21]
  wire  T_49604 = rob_head == 5'h10; // @[rob.scala 970:26]
  wire  T_49606 = rob_tail == 5'h10; // @[rob.scala 970:50]
  wire  T_49607 = T_49604 & T_49606; // @[rob.scala 970:40]
  wire [7:0] T_49616 = T_49606 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49617 = T_49604 ? 8'h48 : T_49616; // @[rob.scala 971:18]
  wire [7:0] T_49618 = T_49607 ? 8'h42 : T_49617; // @[rob.scala 970:18]
  wire [7:0] T_49628 = T_23706_16 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49631 = T_35634_16 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_32_busy = T_23710_T_34690_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49634 = debug_entry_32_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_33_busy = T_35638_T_46618_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49637 = debug_entry_33_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_32_uop_pc = T_34800[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49638 = debug_entry_32_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_33_uop_pc = T_46728[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49639 = debug_entry_33_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_32_exception = T_28311_T_34802_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49650 = debug_entry_32_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_33_exception = T_40239_T_46730_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49653 = debug_entry_33_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49656 = T_26182_16_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49658 = T_26182_16_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49660 = T_26182_16_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49662 = T_26182_16_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49665 = T_49662 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49666 = T_49660 ? 8'h66 : T_49665; // @[rob.scala 1050:21]
  wire [7:0] T_49667 = T_49658 ? 8'h43 : T_49666; // @[rob.scala 1049:21]
  wire [7:0] T_49668 = T_49656 ? 8'h58 : T_49667; // @[rob.scala 1048:21]
  wire  T_49671 = T_38110_16_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49673 = T_38110_16_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49675 = T_38110_16_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49677 = T_38110_16_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49680 = T_49677 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49681 = T_49675 ? 8'h66 : T_49680; // @[rob.scala 1050:21]
  wire [7:0] T_49682 = T_49673 ? 8'h43 : T_49681; // @[rob.scala 1049:21]
  wire [7:0] T_49683 = T_49671 ? 8'h58 : T_49682; // @[rob.scala 1048:21]
  wire  T_49690 = rob_head == 5'h11; // @[rob.scala 970:26]
  wire  T_49692 = rob_tail == 5'h11; // @[rob.scala 970:50]
  wire  T_49693 = T_49690 & T_49692; // @[rob.scala 970:40]
  wire [7:0] T_49702 = T_49692 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49703 = T_49690 ? 8'h48 : T_49702; // @[rob.scala 971:18]
  wire [7:0] T_49704 = T_49693 ? 8'h42 : T_49703; // @[rob.scala 970:18]
  wire [7:0] T_49714 = T_23706_17 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49717 = T_35634_17 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_34_busy = T_23710_T_34804_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49720 = debug_entry_34_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_35_busy = T_35638_T_46732_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49723 = debug_entry_35_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_34_uop_pc = T_34914[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49724 = debug_entry_34_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_35_uop_pc = T_46842[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49725 = debug_entry_35_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_34_exception = T_28311_T_34916_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49736 = debug_entry_34_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_35_exception = T_40239_T_46844_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49739 = debug_entry_35_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49742 = T_26182_17_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49744 = T_26182_17_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49746 = T_26182_17_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49748 = T_26182_17_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49751 = T_49748 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49752 = T_49746 ? 8'h66 : T_49751; // @[rob.scala 1050:21]
  wire [7:0] T_49753 = T_49744 ? 8'h43 : T_49752; // @[rob.scala 1049:21]
  wire [7:0] T_49754 = T_49742 ? 8'h58 : T_49753; // @[rob.scala 1048:21]
  wire  T_49757 = T_38110_17_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49759 = T_38110_17_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49761 = T_38110_17_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49763 = T_38110_17_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49766 = T_49763 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49767 = T_49761 ? 8'h66 : T_49766; // @[rob.scala 1050:21]
  wire [7:0] T_49768 = T_49759 ? 8'h43 : T_49767; // @[rob.scala 1049:21]
  wire [7:0] T_49769 = T_49757 ? 8'h58 : T_49768; // @[rob.scala 1048:21]
  wire  T_49776 = rob_head == 5'h12; // @[rob.scala 970:26]
  wire  T_49778 = rob_tail == 5'h12; // @[rob.scala 970:50]
  wire  T_49779 = T_49776 & T_49778; // @[rob.scala 970:40]
  wire [7:0] T_49788 = T_49778 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49789 = T_49776 ? 8'h48 : T_49788; // @[rob.scala 971:18]
  wire [7:0] T_49790 = T_49779 ? 8'h42 : T_49789; // @[rob.scala 970:18]
  wire [7:0] T_49800 = T_23706_18 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49803 = T_35634_18 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_36_busy = T_23710_T_34918_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49806 = debug_entry_36_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_37_busy = T_35638_T_46846_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49809 = debug_entry_37_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_36_uop_pc = T_35028[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49810 = debug_entry_36_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_37_uop_pc = T_46956[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49811 = debug_entry_37_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_36_exception = T_28311_T_35030_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49822 = debug_entry_36_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_37_exception = T_40239_T_46958_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49825 = debug_entry_37_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49828 = T_26182_18_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49830 = T_26182_18_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49832 = T_26182_18_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49834 = T_26182_18_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49837 = T_49834 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49838 = T_49832 ? 8'h66 : T_49837; // @[rob.scala 1050:21]
  wire [7:0] T_49839 = T_49830 ? 8'h43 : T_49838; // @[rob.scala 1049:21]
  wire [7:0] T_49840 = T_49828 ? 8'h58 : T_49839; // @[rob.scala 1048:21]
  wire  T_49843 = T_38110_18_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49845 = T_38110_18_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49847 = T_38110_18_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49849 = T_38110_18_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49852 = T_49849 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49853 = T_49847 ? 8'h66 : T_49852; // @[rob.scala 1050:21]
  wire [7:0] T_49854 = T_49845 ? 8'h43 : T_49853; // @[rob.scala 1049:21]
  wire [7:0] T_49855 = T_49843 ? 8'h58 : T_49854; // @[rob.scala 1048:21]
  wire  T_49862 = rob_head == 5'h13; // @[rob.scala 970:26]
  wire  T_49864 = rob_tail == 5'h13; // @[rob.scala 970:50]
  wire  T_49865 = T_49862 & T_49864; // @[rob.scala 970:40]
  wire [7:0] T_49874 = T_49864 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49875 = T_49862 ? 8'h48 : T_49874; // @[rob.scala 971:18]
  wire [7:0] T_49876 = T_49865 ? 8'h42 : T_49875; // @[rob.scala 970:18]
  wire [7:0] T_49886 = T_23706_19 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49889 = T_35634_19 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_38_busy = T_23710_T_35032_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49892 = debug_entry_38_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_39_busy = T_35638_T_46960_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49895 = debug_entry_39_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_38_uop_pc = T_35142[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49896 = debug_entry_38_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_39_uop_pc = T_47070[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49897 = debug_entry_39_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_38_exception = T_28311_T_35144_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49908 = debug_entry_38_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_39_exception = T_40239_T_47072_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49911 = debug_entry_39_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_49914 = T_26182_19_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49916 = T_26182_19_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49918 = T_26182_19_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49920 = T_26182_19_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49923 = T_49920 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49924 = T_49918 ? 8'h66 : T_49923; // @[rob.scala 1050:21]
  wire [7:0] T_49925 = T_49916 ? 8'h43 : T_49924; // @[rob.scala 1049:21]
  wire [7:0] T_49926 = T_49914 ? 8'h58 : T_49925; // @[rob.scala 1048:21]
  wire  T_49929 = T_38110_19_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_49931 = T_38110_19_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_49933 = T_38110_19_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_49935 = T_38110_19_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_49938 = T_49935 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_49939 = T_49933 ? 8'h66 : T_49938; // @[rob.scala 1050:21]
  wire [7:0] T_49940 = T_49931 ? 8'h43 : T_49939; // @[rob.scala 1049:21]
  wire [7:0] T_49941 = T_49929 ? 8'h58 : T_49940; // @[rob.scala 1048:21]
  wire  T_49948 = rob_head == 5'h14; // @[rob.scala 970:26]
  wire  T_49950 = rob_tail == 5'h14; // @[rob.scala 970:50]
  wire  T_49951 = T_49948 & T_49950; // @[rob.scala 970:40]
  wire [7:0] T_49960 = T_49950 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_49961 = T_49948 ? 8'h48 : T_49960; // @[rob.scala 971:18]
  wire [7:0] T_49962 = T_49951 ? 8'h42 : T_49961; // @[rob.scala 970:18]
  wire [7:0] T_49972 = T_23706_20 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_49975 = T_35634_20 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_40_busy = T_23710_T_35146_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49978 = debug_entry_40_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_41_busy = T_35638_T_47074_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_49981 = debug_entry_41_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_40_uop_pc = T_35256[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_49982 = debug_entry_40_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_41_uop_pc = T_47184[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_49983 = debug_entry_41_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_40_exception = T_28311_T_35258_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49994 = debug_entry_40_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_41_exception = T_40239_T_47186_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_49997 = debug_entry_41_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_50000 = T_26182_20_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50002 = T_26182_20_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50004 = T_26182_20_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50006 = T_26182_20_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50009 = T_50006 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50010 = T_50004 ? 8'h66 : T_50009; // @[rob.scala 1050:21]
  wire [7:0] T_50011 = T_50002 ? 8'h43 : T_50010; // @[rob.scala 1049:21]
  wire [7:0] T_50012 = T_50000 ? 8'h58 : T_50011; // @[rob.scala 1048:21]
  wire  T_50015 = T_38110_20_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50017 = T_38110_20_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50019 = T_38110_20_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50021 = T_38110_20_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50024 = T_50021 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50025 = T_50019 ? 8'h66 : T_50024; // @[rob.scala 1050:21]
  wire [7:0] T_50026 = T_50017 ? 8'h43 : T_50025; // @[rob.scala 1049:21]
  wire [7:0] T_50027 = T_50015 ? 8'h58 : T_50026; // @[rob.scala 1048:21]
  wire  T_50034 = rob_head == 5'h15; // @[rob.scala 970:26]
  wire  T_50036 = rob_tail == 5'h15; // @[rob.scala 970:50]
  wire  T_50037 = T_50034 & T_50036; // @[rob.scala 970:40]
  wire [7:0] T_50046 = T_50036 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_50047 = T_50034 ? 8'h48 : T_50046; // @[rob.scala 971:18]
  wire [7:0] T_50048 = T_50037 ? 8'h42 : T_50047; // @[rob.scala 970:18]
  wire [7:0] T_50058 = T_23706_21 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_50061 = T_35634_21 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_42_busy = T_23710_T_35260_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_50064 = debug_entry_42_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_43_busy = T_35638_T_47188_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_50067 = debug_entry_43_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_42_uop_pc = T_35370[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_50068 = debug_entry_42_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_43_uop_pc = T_47298[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_50069 = debug_entry_43_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_42_exception = T_28311_T_35372_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_50080 = debug_entry_42_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_43_exception = T_40239_T_47300_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_50083 = debug_entry_43_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_50086 = T_26182_21_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50088 = T_26182_21_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50090 = T_26182_21_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50092 = T_26182_21_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50095 = T_50092 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50096 = T_50090 ? 8'h66 : T_50095; // @[rob.scala 1050:21]
  wire [7:0] T_50097 = T_50088 ? 8'h43 : T_50096; // @[rob.scala 1049:21]
  wire [7:0] T_50098 = T_50086 ? 8'h58 : T_50097; // @[rob.scala 1048:21]
  wire  T_50101 = T_38110_21_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50103 = T_38110_21_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50105 = T_38110_21_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50107 = T_38110_21_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50110 = T_50107 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50111 = T_50105 ? 8'h66 : T_50110; // @[rob.scala 1050:21]
  wire [7:0] T_50112 = T_50103 ? 8'h43 : T_50111; // @[rob.scala 1049:21]
  wire [7:0] T_50113 = T_50101 ? 8'h58 : T_50112; // @[rob.scala 1048:21]
  wire  T_50120 = rob_head == 5'h16; // @[rob.scala 970:26]
  wire  T_50122 = rob_tail == 5'h16; // @[rob.scala 970:50]
  wire  T_50123 = T_50120 & T_50122; // @[rob.scala 970:40]
  wire [7:0] T_50132 = T_50122 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_50133 = T_50120 ? 8'h48 : T_50132; // @[rob.scala 971:18]
  wire [7:0] T_50134 = T_50123 ? 8'h42 : T_50133; // @[rob.scala 970:18]
  wire [7:0] T_50144 = T_23706_22 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_50147 = T_35634_22 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_44_busy = T_23710_T_35374_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_50150 = debug_entry_44_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_45_busy = T_35638_T_47302_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_50153 = debug_entry_45_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_44_uop_pc = T_35484[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_50154 = debug_entry_44_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_45_uop_pc = T_47412[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_50155 = debug_entry_45_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_44_exception = T_28311_T_35486_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_50166 = debug_entry_44_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_45_exception = T_40239_T_47414_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_50169 = debug_entry_45_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_50172 = T_26182_22_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50174 = T_26182_22_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50176 = T_26182_22_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50178 = T_26182_22_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50181 = T_50178 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50182 = T_50176 ? 8'h66 : T_50181; // @[rob.scala 1050:21]
  wire [7:0] T_50183 = T_50174 ? 8'h43 : T_50182; // @[rob.scala 1049:21]
  wire [7:0] T_50184 = T_50172 ? 8'h58 : T_50183; // @[rob.scala 1048:21]
  wire  T_50187 = T_38110_22_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50189 = T_38110_22_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50191 = T_38110_22_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50193 = T_38110_22_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50196 = T_50193 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50197 = T_50191 ? 8'h66 : T_50196; // @[rob.scala 1050:21]
  wire [7:0] T_50198 = T_50189 ? 8'h43 : T_50197; // @[rob.scala 1049:21]
  wire [7:0] T_50199 = T_50187 ? 8'h58 : T_50198; // @[rob.scala 1048:21]
  wire  T_50209 = T_48136 & T_48178; // @[rob.scala 970:40]
  wire [7:0] T_50218 = T_48178 ? 8'h54 : 8'h20; // @[rob.scala 972:18]
  wire [7:0] T_50219 = T_48136 ? 8'h48 : T_50218; // @[rob.scala 971:18]
  wire [7:0] T_50220 = T_50209 ? 8'h42 : T_50219; // @[rob.scala 970:18]
  wire [7:0] T_50230 = T_23706_23 ? 8'h56 : 8'h20; // @[rob.scala 996:21]
  wire [7:0] T_50233 = T_35634_23 ? 8'h56 : 8'h20; // @[rob.scala 997:21]
  wire  debug_entry_46_busy = T_23710_T_35488_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_50236 = debug_entry_46_busy ? 8'h42 : 8'h20; // @[rob.scala 998:21]
  wire  debug_entry_47_busy = T_35638_T_47416_data; // @[rob.scala 240:26 rob.scala 552:43]
  wire [7:0] T_50239 = debug_entry_47_busy ? 8'h42 : 8'h20; // @[rob.scala 999:21]
  wire [39:0] debug_entry_46_uop_pc = T_35598[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [31:0] T_50240 = debug_entry_46_uop_pc[31:0]; // @[rob.scala 1000:45]
  wire [39:0] debug_entry_47_uop_pc = T_47526[39:0]; // @[rob.scala 240:26 rob.scala 554:45]
  wire [15:0] T_50241 = debug_entry_47_uop_pc[15:0]; // @[rob.scala 1001:45]
  wire  debug_entry_46_exception = T_28311_T_35600_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_50252 = debug_entry_46_exception ? 8'h45 : 8'h2d; // @[rob.scala 1007:21]
  wire  debug_entry_47_exception = T_40239_T_47528_data; // @[rob.scala 240:26 rob.scala 555:48]
  wire [7:0] T_50255 = debug_entry_47_exception ? 8'h45 : 8'h2d; // @[rob.scala 1008:21]
  wire  T_50258 = T_26182_23_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50260 = T_26182_23_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50262 = T_26182_23_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50264 = T_26182_23_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50267 = T_50264 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50268 = T_50262 ? 8'h66 : T_50267; // @[rob.scala 1050:21]
  wire [7:0] T_50269 = T_50260 ? 8'h43 : T_50268; // @[rob.scala 1049:21]
  wire [7:0] T_50270 = T_50258 ? 8'h58 : T_50269; // @[rob.scala 1048:21]
  wire  T_50273 = T_38110_23_dst_rtype == 2'h0; // @[rob.scala 1048:58]
  wire  T_50275 = T_38110_23_dst_rtype == 2'h3; // @[rob.scala 1049:58]
  wire  T_50277 = T_38110_23_dst_rtype == 2'h1; // @[rob.scala 1050:58]
  wire  T_50279 = T_38110_23_dst_rtype == 2'h2; // @[rob.scala 1051:58]
  wire [7:0] T_50282 = T_50279 ? 8'h2d : 8'h3f; // @[rob.scala 1051:21]
  wire [7:0] T_50283 = T_50277 ? 8'h66 : T_50282; // @[rob.scala 1050:21]
  wire [7:0] T_50284 = T_50275 ? 8'h43 : T_50283; // @[rob.scala 1049:21]
  wire [7:0] T_50285 = T_50273 ? 8'h58 : T_50284; // @[rob.scala 1048:21]
  wire [5:0] new_DoPrim0 = {{1'd0}, rob_tail};
  wire  new_DoPrim1 = T_47543 & T_47545;
  wire  new_DoPrim2 = T_47560 & T_47562;
  wire  new_DoPrim4401855 = T_47635 | T_47664;
  wire [4:0] new_DoPrim4401856 = T_47637 | T_47666;
  wire  new_DoPrim4401857 = io_com_valids_0 & rob_head_is_store_0;
  wire  new_DoPrim4401858 = io_com_valids_1 & rob_head_is_store_1;
  wire  new_DoPrim4401859 = io_com_valids_0 & rob_head_is_load_0;
  wire  new_DoPrim4401860 = io_com_valids_1 & rob_head_is_load_1;
  wire  new_DoPrim4430078 = T_47568 & T_47572;
  wire  new_DoPrim4430080 = will_throw_exception | io_cxcpt_valid;
  wire  new_DoPrim4430081 = T_29099 & T_29272;
  wire  new_DoPrim4430082 = T_41027 & T_41200;
  wire [63:0] new_DoPrim4430083 = {T_47581,r_xcpt_badvaddr};
  wire [39:0] new_DoPrim4430084 = T_23619[39:0];
  wire  new_DoPrim4430086 = rob_pc_hob_next_val | T_23559;
  wire [39:0] new_DoPrim4430087 = T_23644[39:0];
  wire  new_DoPrim4430089 = T_47568 | T_47615;
  wire [39:0] new_DoPrim4430090 = T_47612[39:0];
  wire  new_DoPrim4430092 = T_23670 | T_23671;
  wire  new_DoPrim4430093 = T_48130 & T_48194;
  wire  new_DoPrim4430094 = T_48196 & T_48198;
  wire  new_DoPrim4430095 = T_48134 & row_metadata_has_brorjalr_T_23664_data;
  wire [5:0] new_DoPrim4430098 = {{1'd0}, rob_head};
  wire [63:0] new_DoPrim4430178 = {{24'd0}, r_xcpt_badvaddr};
  wire  new_DoPrim113799324 = T_47568 & T_47569;
  wire  new_DoPrim113799325 = T_47568 | T_47615;
  wire [3:0] new_DoPrim113799327 = T_23586[3:0];
  wire [3:0] new_DoPrim113799474 = T_47586[3:0];
  wire  new_DoPrim113799476 = T_23559 & T_23568;
  wire [3:0] new_DoPrim113799477 = T_23565[3:0];
  wire [36:0] new_DoPrim113799479 = T_23562[36:0];
  wire [3:0] new_DoPrim113799482 = T_23576[3:0];
  wire  new_DoPrim113799628 = rob_head[0];
  wire [3:0] new_DoPrim113799629 = T_47586[3:0];
  wire  new_DoPrim113799631 = T_23559 & T_23563;
  wire [3:0] new_DoPrim113799632 = T_23565[3:0];
  wire [36:0] new_DoPrim113799634 = T_23562[36:0];
  wire [4:0] new_DoPrim113799640 = T_23573[4:0];
  wire  new_DoPrim113799714 = T_23559 & io_dis_new_packet;
  wire  new_DoPrim113799794 = T_23559 & io_dis_new_packet;
  wire  new_DoPrim113799882 = ~(io_dis_uops_0_is_fence | io_dis_uops_0_is_fencei);
  wire  new_DoPrim113799884 = io_wb_resps_0_valid & T_28592;
  wire [4:0] new_DoPrim113799885 = T_28589[4:0];
  wire  new_DoPrim113799889 = io_wb_resps_1_valid & T_28600;
  wire [4:0] new_DoPrim113799890 = T_28597[4:0];
  wire  new_DoPrim113799894 = io_wb_resps_2_valid & T_28608;
  wire [4:0] new_DoPrim113799895 = T_28605[4:0];
  wire  new_DoPrim113799899 = io_lsu_clr_bsy_valid & T_28614;
  wire [4:0] new_DoPrim113799900 = T_28617[4:0];
  wire  new_DoPrim113799984 = io_lxcpt_valid & T_29075;
  wire [4:0] new_DoPrim113799985 = T_29078[4:0];
  wire  new_DoPrim113799989 = io_bxcpt_valid & T_29083;
  wire [4:0] new_DoPrim113799990 = T_29086[4:0];
  wire  new_DoPrim113799994 = rob_state == 2'h2;
  wire  new_DoPrim113828224 = io_fflags_0_valid & T_29061;
  wire [4:0] new_DoPrim113828225 = T_29064[4:0];
  wire  new_DoPrim113828229 = io_fflags_1_valid & T_29068;
  wire [4:0] new_DoPrim113828230 = T_29071[4:0];
  wire  new_DoPrim113828312 = ~(io_dis_uops_1_is_fence | io_dis_uops_1_is_fencei);
  wire  new_DoPrim113828314 = io_wb_resps_0_valid & T_28590;
  wire [4:0] new_DoPrim113828315 = T_28589[4:0];
  wire  new_DoPrim113828319 = io_wb_resps_1_valid & T_28598;
  wire [4:0] new_DoPrim113828320 = T_28597[4:0];
  wire  new_DoPrim113828324 = io_wb_resps_2_valid & T_28606;
  wire [4:0] new_DoPrim113828325 = T_28605[4:0];
  wire  new_DoPrim113828329 = io_lsu_clr_bsy_valid & T_28612;
  wire [4:0] new_DoPrim113828330 = T_28617[4:0];
  wire  new_DoPrim113828414 = io_lxcpt_valid & T_29073;
  wire [4:0] new_DoPrim113828415 = T_29078[4:0];
  wire  new_DoPrim113828419 = io_bxcpt_valid & T_29081;
  wire [4:0] new_DoPrim113828420 = T_29086[4:0];
  wire  new_DoPrim113828424 = rob_state == 2'h2;
  wire  new_DoPrim113856654 = io_fflags_0_valid & T_29059;
  wire [4:0] new_DoPrim113856655 = T_29064[4:0];
  wire  new_DoPrim113856659 = io_fflags_1_valid & T_29066;
  wire [4:0] new_DoPrim113856660 = T_29071[4:0];
  assign T_23555_T_23587_addr = new_DoPrim113799327;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_23587_data = T_23555[T_23555_T_23587_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_23587_data = T_23555_T_23587_addr >= 4'hc ? _RAND_1[36:0] : T_23555[T_23555_T_23587_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_32958_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_32958_data = T_23555[T_23555_T_32958_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_32958_data = T_23555_T_32958_addr >= 4'hc ? _RAND_2[36:0] : T_23555[T_23555_T_32958_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33072_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33072_data = T_23555[T_23555_T_33072_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33072_data = T_23555_T_33072_addr >= 4'hc ? _RAND_3[36:0] : T_23555[T_23555_T_33072_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33186_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33186_data = T_23555[T_23555_T_33186_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33186_data = T_23555_T_33186_addr >= 4'hc ? _RAND_4[36:0] : T_23555[T_23555_T_33186_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33300_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33300_data = T_23555[T_23555_T_33300_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33300_data = T_23555_T_33300_addr >= 4'hc ? _RAND_5[36:0] : T_23555[T_23555_T_33300_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33414_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33414_data = T_23555[T_23555_T_33414_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33414_data = T_23555_T_33414_addr >= 4'hc ? _RAND_6[36:0] : T_23555[T_23555_T_33414_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33528_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33528_data = T_23555[T_23555_T_33528_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33528_data = T_23555_T_33528_addr >= 4'hc ? _RAND_7[36:0] : T_23555[T_23555_T_33528_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33642_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33642_data = T_23555[T_23555_T_33642_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33642_data = T_23555_T_33642_addr >= 4'hc ? _RAND_8[36:0] : T_23555[T_23555_T_33642_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33756_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33756_data = T_23555[T_23555_T_33756_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33756_data = T_23555_T_33756_addr >= 4'hc ? _RAND_9[36:0] : T_23555[T_23555_T_33756_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33870_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33870_data = T_23555[T_23555_T_33870_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33870_data = T_23555_T_33870_addr >= 4'hc ? _RAND_10[36:0] : T_23555[T_23555_T_33870_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33984_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_33984_data = T_23555[T_23555_T_33984_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_33984_data = T_23555_T_33984_addr >= 4'hc ? _RAND_11[36:0] : T_23555[T_23555_T_33984_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34098_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34098_data = T_23555[T_23555_T_34098_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34098_data = T_23555_T_34098_addr >= 4'hc ? _RAND_12[36:0] : T_23555[T_23555_T_34098_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34212_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34212_data = T_23555[T_23555_T_34212_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34212_data = T_23555_T_34212_addr >= 4'hc ? _RAND_13[36:0] : T_23555[T_23555_T_34212_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34326_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34326_data = T_23555[T_23555_T_34326_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34326_data = T_23555_T_34326_addr >= 4'hc ? _RAND_14[36:0] : T_23555[T_23555_T_34326_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34440_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34440_data = T_23555[T_23555_T_34440_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34440_data = T_23555_T_34440_addr >= 4'hc ? _RAND_15[36:0] : T_23555[T_23555_T_34440_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34554_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34554_data = T_23555[T_23555_T_34554_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34554_data = T_23555_T_34554_addr >= 4'hc ? _RAND_16[36:0] : T_23555[T_23555_T_34554_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34668_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34668_data = T_23555[T_23555_T_34668_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34668_data = T_23555_T_34668_addr >= 4'hc ? _RAND_17[36:0] : T_23555[T_23555_T_34668_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34782_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34782_data = T_23555[T_23555_T_34782_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34782_data = T_23555_T_34782_addr >= 4'hc ? _RAND_18[36:0] : T_23555[T_23555_T_34782_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34896_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_34896_data = T_23555[T_23555_T_34896_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_34896_data = T_23555_T_34896_addr >= 4'hc ? _RAND_19[36:0] : T_23555[T_23555_T_34896_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35010_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35010_data = T_23555[T_23555_T_35010_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_35010_data = T_23555_T_35010_addr >= 4'hc ? _RAND_20[36:0] : T_23555[T_23555_T_35010_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35124_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35124_data = T_23555[T_23555_T_35124_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_35124_data = T_23555_T_35124_addr >= 4'hc ? _RAND_21[36:0] : T_23555[T_23555_T_35124_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35238_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35238_data = T_23555[T_23555_T_35238_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_35238_data = T_23555_T_35238_addr >= 4'hc ? _RAND_22[36:0] : T_23555[T_23555_T_35238_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35352_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35352_data = T_23555[T_23555_T_35352_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_35352_data = T_23555_T_35352_addr >= 4'hc ? _RAND_23[36:0] : T_23555[T_23555_T_35352_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35466_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35466_data = T_23555[T_23555_T_35466_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_35466_data = T_23555_T_35466_addr >= 4'hc ? _RAND_24[36:0] : T_23555[T_23555_T_35466_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35580_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_35580_data = T_23555[T_23555_T_35580_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_35580_data = T_23555_T_35580_addr >= 4'hc ? _RAND_25[36:0] : T_23555[T_23555_T_35580_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_44886_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_44886_data = T_23555[T_23555_T_44886_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_44886_data = T_23555_T_44886_addr >= 4'hc ? _RAND_26[36:0] : T_23555[T_23555_T_44886_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45000_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45000_data = T_23555[T_23555_T_45000_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45000_data = T_23555_T_45000_addr >= 4'hc ? _RAND_27[36:0] : T_23555[T_23555_T_45000_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45114_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45114_data = T_23555[T_23555_T_45114_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45114_data = T_23555_T_45114_addr >= 4'hc ? _RAND_28[36:0] : T_23555[T_23555_T_45114_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45228_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45228_data = T_23555[T_23555_T_45228_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45228_data = T_23555_T_45228_addr >= 4'hc ? _RAND_29[36:0] : T_23555[T_23555_T_45228_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45342_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45342_data = T_23555[T_23555_T_45342_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45342_data = T_23555_T_45342_addr >= 4'hc ? _RAND_30[36:0] : T_23555[T_23555_T_45342_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45456_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45456_data = T_23555[T_23555_T_45456_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45456_data = T_23555_T_45456_addr >= 4'hc ? _RAND_31[36:0] : T_23555[T_23555_T_45456_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45570_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45570_data = T_23555[T_23555_T_45570_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45570_data = T_23555_T_45570_addr >= 4'hc ? _RAND_32[36:0] : T_23555[T_23555_T_45570_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45684_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45684_data = T_23555[T_23555_T_45684_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45684_data = T_23555_T_45684_addr >= 4'hc ? _RAND_33[36:0] : T_23555[T_23555_T_45684_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45798_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45798_data = T_23555[T_23555_T_45798_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45798_data = T_23555_T_45798_addr >= 4'hc ? _RAND_34[36:0] : T_23555[T_23555_T_45798_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45912_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_45912_data = T_23555[T_23555_T_45912_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_45912_data = T_23555_T_45912_addr >= 4'hc ? _RAND_35[36:0] : T_23555[T_23555_T_45912_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46026_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46026_data = T_23555[T_23555_T_46026_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46026_data = T_23555_T_46026_addr >= 4'hc ? _RAND_36[36:0] : T_23555[T_23555_T_46026_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46140_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46140_data = T_23555[T_23555_T_46140_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46140_data = T_23555_T_46140_addr >= 4'hc ? _RAND_37[36:0] : T_23555[T_23555_T_46140_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46254_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46254_data = T_23555[T_23555_T_46254_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46254_data = T_23555_T_46254_addr >= 4'hc ? _RAND_38[36:0] : T_23555[T_23555_T_46254_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46368_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46368_data = T_23555[T_23555_T_46368_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46368_data = T_23555_T_46368_addr >= 4'hc ? _RAND_39[36:0] : T_23555[T_23555_T_46368_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46482_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46482_data = T_23555[T_23555_T_46482_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46482_data = T_23555_T_46482_addr >= 4'hc ? _RAND_40[36:0] : T_23555[T_23555_T_46482_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46596_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46596_data = T_23555[T_23555_T_46596_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46596_data = T_23555_T_46596_addr >= 4'hc ? _RAND_41[36:0] : T_23555[T_23555_T_46596_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46710_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46710_data = T_23555[T_23555_T_46710_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46710_data = T_23555_T_46710_addr >= 4'hc ? _RAND_42[36:0] : T_23555[T_23555_T_46710_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46824_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46824_data = T_23555[T_23555_T_46824_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46824_data = T_23555_T_46824_addr >= 4'hc ? _RAND_43[36:0] : T_23555[T_23555_T_46824_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46938_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_46938_data = T_23555[T_23555_T_46938_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_46938_data = T_23555_T_46938_addr >= 4'hc ? _RAND_44[36:0] : T_23555[T_23555_T_46938_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47052_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47052_data = T_23555[T_23555_T_47052_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_47052_data = T_23555_T_47052_addr >= 4'hc ? _RAND_45[36:0] : T_23555[T_23555_T_47052_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47166_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47166_data = T_23555[T_23555_T_47166_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_47166_data = T_23555_T_47166_addr >= 4'hc ? _RAND_46[36:0] : T_23555[T_23555_T_47166_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47280_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47280_data = T_23555[T_23555_T_47280_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_47280_data = T_23555_T_47280_addr >= 4'hc ? _RAND_47[36:0] : T_23555[T_23555_T_47280_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47394_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47394_data = T_23555[T_23555_T_47394_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_47394_data = T_23555_T_47394_addr >= 4'hc ? _RAND_48[36:0] : T_23555[T_23555_T_47394_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47508_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47508_data = T_23555[T_23555_T_47508_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_47508_data = T_23555_T_47508_addr >= 4'hc ? _RAND_49[36:0] : T_23555[T_23555_T_47508_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47587_addr = new_DoPrim113799474;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_47587_data = T_23555[T_23555_T_47587_addr]; // @[rob.scala 893:22]
  `else
  assign T_23555_T_47587_data = T_23555_T_47587_addr >= 4'hc ? _RAND_50[36:0] : T_23555[T_23555_T_47587_addr]; // @[rob.scala 893:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23555_T_23571_data = new_DoPrim113799479;
  assign T_23555_T_23571_addr = new_DoPrim113799477;
  assign T_23555_T_23571_mask = 1'h1;
  assign T_23555_T_23571_en = new_DoPrim113799476;
  assign T_23558_T_23592_addr = new_DoPrim113799482;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_23592_data = T_23558[T_23558_T_23592_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_23592_data = T_23558_T_23592_addr >= 4'hc ? _RAND_52[36:0] : T_23558[T_23558_T_23592_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_32964_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_32964_data = T_23558[T_23558_T_32964_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_32964_data = T_23558_T_32964_addr >= 4'hc ? _RAND_53[36:0] : T_23558[T_23558_T_32964_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33078_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33078_data = T_23558[T_23558_T_33078_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33078_data = T_23558_T_33078_addr >= 4'hc ? _RAND_54[36:0] : T_23558[T_23558_T_33078_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33192_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33192_data = T_23558[T_23558_T_33192_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33192_data = T_23558_T_33192_addr >= 4'hc ? _RAND_55[36:0] : T_23558[T_23558_T_33192_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33306_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33306_data = T_23558[T_23558_T_33306_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33306_data = T_23558_T_33306_addr >= 4'hc ? _RAND_56[36:0] : T_23558[T_23558_T_33306_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33420_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33420_data = T_23558[T_23558_T_33420_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33420_data = T_23558_T_33420_addr >= 4'hc ? _RAND_57[36:0] : T_23558[T_23558_T_33420_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33534_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33534_data = T_23558[T_23558_T_33534_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33534_data = T_23558_T_33534_addr >= 4'hc ? _RAND_58[36:0] : T_23558[T_23558_T_33534_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33648_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33648_data = T_23558[T_23558_T_33648_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33648_data = T_23558_T_33648_addr >= 4'hc ? _RAND_59[36:0] : T_23558[T_23558_T_33648_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33762_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33762_data = T_23558[T_23558_T_33762_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33762_data = T_23558_T_33762_addr >= 4'hc ? _RAND_60[36:0] : T_23558[T_23558_T_33762_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33876_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33876_data = T_23558[T_23558_T_33876_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33876_data = T_23558_T_33876_addr >= 4'hc ? _RAND_61[36:0] : T_23558[T_23558_T_33876_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33990_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_33990_data = T_23558[T_23558_T_33990_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_33990_data = T_23558_T_33990_addr >= 4'hc ? _RAND_62[36:0] : T_23558[T_23558_T_33990_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34104_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34104_data = T_23558[T_23558_T_34104_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34104_data = T_23558_T_34104_addr >= 4'hc ? _RAND_63[36:0] : T_23558[T_23558_T_34104_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34218_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34218_data = T_23558[T_23558_T_34218_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34218_data = T_23558_T_34218_addr >= 4'hc ? _RAND_64[36:0] : T_23558[T_23558_T_34218_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34332_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34332_data = T_23558[T_23558_T_34332_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34332_data = T_23558_T_34332_addr >= 4'hc ? _RAND_65[36:0] : T_23558[T_23558_T_34332_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34446_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34446_data = T_23558[T_23558_T_34446_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34446_data = T_23558_T_34446_addr >= 4'hc ? _RAND_66[36:0] : T_23558[T_23558_T_34446_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34560_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34560_data = T_23558[T_23558_T_34560_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34560_data = T_23558_T_34560_addr >= 4'hc ? _RAND_67[36:0] : T_23558[T_23558_T_34560_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34674_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34674_data = T_23558[T_23558_T_34674_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34674_data = T_23558_T_34674_addr >= 4'hc ? _RAND_68[36:0] : T_23558[T_23558_T_34674_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34788_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34788_data = T_23558[T_23558_T_34788_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34788_data = T_23558_T_34788_addr >= 4'hc ? _RAND_69[36:0] : T_23558[T_23558_T_34788_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34902_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_34902_data = T_23558[T_23558_T_34902_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_34902_data = T_23558_T_34902_addr >= 4'hc ? _RAND_70[36:0] : T_23558[T_23558_T_34902_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35016_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35016_data = T_23558[T_23558_T_35016_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_35016_data = T_23558_T_35016_addr >= 4'hc ? _RAND_71[36:0] : T_23558[T_23558_T_35016_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35130_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35130_data = T_23558[T_23558_T_35130_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_35130_data = T_23558_T_35130_addr >= 4'hc ? _RAND_72[36:0] : T_23558[T_23558_T_35130_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35244_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35244_data = T_23558[T_23558_T_35244_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_35244_data = T_23558_T_35244_addr >= 4'hc ? _RAND_73[36:0] : T_23558[T_23558_T_35244_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35358_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35358_data = T_23558[T_23558_T_35358_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_35358_data = T_23558_T_35358_addr >= 4'hc ? _RAND_74[36:0] : T_23558[T_23558_T_35358_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35472_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35472_data = T_23558[T_23558_T_35472_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_35472_data = T_23558_T_35472_addr >= 4'hc ? _RAND_75[36:0] : T_23558[T_23558_T_35472_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35586_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_35586_data = T_23558[T_23558_T_35586_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_35586_data = T_23558_T_35586_addr >= 4'hc ? _RAND_76[36:0] : T_23558[T_23558_T_35586_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_44892_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_44892_data = T_23558[T_23558_T_44892_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_44892_data = T_23558_T_44892_addr >= 4'hc ? _RAND_77[36:0] : T_23558[T_23558_T_44892_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45006_addr = 4'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45006_data = T_23558[T_23558_T_45006_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45006_data = T_23558_T_45006_addr >= 4'hc ? _RAND_78[36:0] : T_23558[T_23558_T_45006_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45120_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45120_data = T_23558[T_23558_T_45120_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45120_data = T_23558_T_45120_addr >= 4'hc ? _RAND_79[36:0] : T_23558[T_23558_T_45120_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45234_addr = 4'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45234_data = T_23558[T_23558_T_45234_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45234_data = T_23558_T_45234_addr >= 4'hc ? _RAND_80[36:0] : T_23558[T_23558_T_45234_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45348_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45348_data = T_23558[T_23558_T_45348_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45348_data = T_23558_T_45348_addr >= 4'hc ? _RAND_81[36:0] : T_23558[T_23558_T_45348_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45462_addr = 4'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45462_data = T_23558[T_23558_T_45462_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45462_data = T_23558_T_45462_addr >= 4'hc ? _RAND_82[36:0] : T_23558[T_23558_T_45462_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45576_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45576_data = T_23558[T_23558_T_45576_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45576_data = T_23558_T_45576_addr >= 4'hc ? _RAND_83[36:0] : T_23558[T_23558_T_45576_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45690_addr = 4'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45690_data = T_23558[T_23558_T_45690_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45690_data = T_23558_T_45690_addr >= 4'hc ? _RAND_84[36:0] : T_23558[T_23558_T_45690_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45804_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45804_data = T_23558[T_23558_T_45804_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45804_data = T_23558_T_45804_addr >= 4'hc ? _RAND_85[36:0] : T_23558[T_23558_T_45804_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45918_addr = 4'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_45918_data = T_23558[T_23558_T_45918_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_45918_data = T_23558_T_45918_addr >= 4'hc ? _RAND_86[36:0] : T_23558[T_23558_T_45918_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46032_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46032_data = T_23558[T_23558_T_46032_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46032_data = T_23558_T_46032_addr >= 4'hc ? _RAND_87[36:0] : T_23558[T_23558_T_46032_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46146_addr = 4'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46146_data = T_23558[T_23558_T_46146_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46146_data = T_23558_T_46146_addr >= 4'hc ? _RAND_88[36:0] : T_23558[T_23558_T_46146_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46260_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46260_data = T_23558[T_23558_T_46260_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46260_data = T_23558_T_46260_addr >= 4'hc ? _RAND_89[36:0] : T_23558[T_23558_T_46260_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46374_addr = 4'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46374_data = T_23558[T_23558_T_46374_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46374_data = T_23558_T_46374_addr >= 4'hc ? _RAND_90[36:0] : T_23558[T_23558_T_46374_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46488_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46488_data = T_23558[T_23558_T_46488_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46488_data = T_23558_T_46488_addr >= 4'hc ? _RAND_91[36:0] : T_23558[T_23558_T_46488_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46602_addr = 4'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46602_data = T_23558[T_23558_T_46602_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46602_data = T_23558_T_46602_addr >= 4'hc ? _RAND_92[36:0] : T_23558[T_23558_T_46602_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46716_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46716_data = T_23558[T_23558_T_46716_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46716_data = T_23558_T_46716_addr >= 4'hc ? _RAND_93[36:0] : T_23558[T_23558_T_46716_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46830_addr = 4'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46830_data = T_23558[T_23558_T_46830_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46830_data = T_23558_T_46830_addr >= 4'hc ? _RAND_94[36:0] : T_23558[T_23558_T_46830_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46944_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_46944_data = T_23558[T_23558_T_46944_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_46944_data = T_23558_T_46944_addr >= 4'hc ? _RAND_95[36:0] : T_23558[T_23558_T_46944_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47058_addr = 4'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47058_data = T_23558[T_23558_T_47058_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_47058_data = T_23558_T_47058_addr >= 4'hc ? _RAND_96[36:0] : T_23558[T_23558_T_47058_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47172_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47172_data = T_23558[T_23558_T_47172_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_47172_data = T_23558_T_47172_addr >= 4'hc ? _RAND_97[36:0] : T_23558[T_23558_T_47172_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47286_addr = 4'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47286_data = T_23558[T_23558_T_47286_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_47286_data = T_23558_T_47286_addr >= 4'hc ? _RAND_98[36:0] : T_23558[T_23558_T_47286_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47400_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47400_data = T_23558[T_23558_T_47400_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_47400_data = T_23558_T_47400_addr >= 4'hc ? _RAND_99[36:0] : T_23558[T_23558_T_47400_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47514_addr = 4'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47514_data = T_23558[T_23558_T_47514_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_47514_data = T_23558_T_47514_addr >= 4'hc ? _RAND_100[36:0] : T_23558[T_23558_T_47514_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47593_addr = new_DoPrim113799629;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_47593_data = T_23558[T_23558_T_47593_addr]; // @[rob.scala 894:22]
  `else
  assign T_23558_T_47593_data = T_23558_T_47593_addr >= 4'hc ? _RAND_101[36:0] : T_23558[T_23558_T_47593_addr]; // @[rob.scala 894:22]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23558_T_23566_data = new_DoPrim113799634;
  assign T_23558_T_23566_addr = new_DoPrim113799632;
  assign T_23558_T_23566_mask = 1'h1;
  assign T_23558_T_23566_en = new_DoPrim113799631;
  assign row_metadata_brob_idx_T_23666_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_23666_data = row_metadata_brob_idx[row_metadata_brob_idx_T_23666_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_23666_data = row_metadata_brob_idx_T_23666_addr >= 5'h18 ? _RAND_103[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_23666_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_23669_addr = new_DoPrim113799640;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_23669_data = row_metadata_brob_idx[row_metadata_brob_idx_T_23669_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_23669_data = row_metadata_brob_idx_T_23669_addr >= 5'h18 ? _RAND_104[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_23669_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48247_addr = 5'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48247_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48247_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48247_data = row_metadata_brob_idx_T_48247_addr >= 5'h18 ? _RAND_105[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48247_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48333_addr = 5'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48333_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48333_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48333_data = row_metadata_brob_idx_T_48333_addr >= 5'h18 ? _RAND_106[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48333_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48419_addr = 5'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48419_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48419_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48419_data = row_metadata_brob_idx_T_48419_addr >= 5'h18 ? _RAND_107[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48419_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48505_addr = 5'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48505_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48505_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48505_data = row_metadata_brob_idx_T_48505_addr >= 5'h18 ? _RAND_108[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48505_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48591_addr = 5'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48591_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48591_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48591_data = row_metadata_brob_idx_T_48591_addr >= 5'h18 ? _RAND_109[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48591_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48677_addr = 5'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48677_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48677_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48677_data = row_metadata_brob_idx_T_48677_addr >= 5'h18 ? _RAND_110[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48677_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48763_addr = 5'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48763_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48763_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48763_data = row_metadata_brob_idx_T_48763_addr >= 5'h18 ? _RAND_111[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48763_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48849_addr = 5'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48849_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48849_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48849_data = row_metadata_brob_idx_T_48849_addr >= 5'h18 ? _RAND_112[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48849_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48935_addr = 5'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_48935_data = row_metadata_brob_idx[row_metadata_brob_idx_T_48935_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_48935_data = row_metadata_brob_idx_T_48935_addr >= 5'h18 ? _RAND_113[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_48935_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49021_addr = 5'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49021_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49021_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49021_data = row_metadata_brob_idx_T_49021_addr >= 5'h18 ? _RAND_114[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49021_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49107_addr = 5'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49107_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49107_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49107_data = row_metadata_brob_idx_T_49107_addr >= 5'h18 ? _RAND_115[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49107_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49193_addr = 5'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49193_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49193_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49193_data = row_metadata_brob_idx_T_49193_addr >= 5'h18 ? _RAND_116[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49193_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49279_addr = 5'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49279_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49279_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49279_data = row_metadata_brob_idx_T_49279_addr >= 5'h18 ? _RAND_117[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49279_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49365_addr = 5'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49365_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49365_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49365_data = row_metadata_brob_idx_T_49365_addr >= 5'h18 ? _RAND_118[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49365_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49451_addr = 5'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49451_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49451_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49451_data = row_metadata_brob_idx_T_49451_addr >= 5'h18 ? _RAND_119[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49451_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49537_addr = 5'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49537_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49537_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49537_data = row_metadata_brob_idx_T_49537_addr >= 5'h18 ? _RAND_120[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49537_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49623_addr = 5'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49623_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49623_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49623_data = row_metadata_brob_idx_T_49623_addr >= 5'h18 ? _RAND_121[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49623_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49709_addr = 5'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49709_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49709_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49709_data = row_metadata_brob_idx_T_49709_addr >= 5'h18 ? _RAND_122[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49709_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49795_addr = 5'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49795_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49795_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49795_data = row_metadata_brob_idx_T_49795_addr >= 5'h18 ? _RAND_123[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49795_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49881_addr = 5'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49881_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49881_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49881_data = row_metadata_brob_idx_T_49881_addr >= 5'h18 ? _RAND_124[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49881_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49967_addr = 5'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_49967_data = row_metadata_brob_idx[row_metadata_brob_idx_T_49967_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_49967_data = row_metadata_brob_idx_T_49967_addr >= 5'h18 ? _RAND_125[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_49967_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_50053_addr = 5'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_50053_data = row_metadata_brob_idx[row_metadata_brob_idx_T_50053_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_50053_data = row_metadata_brob_idx_T_50053_addr >= 5'h18 ? _RAND_126[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_50053_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_50139_addr = 5'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_50139_data = row_metadata_brob_idx[row_metadata_brob_idx_T_50139_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_50139_data = row_metadata_brob_idx_T_50139_addr >= 5'h18 ? _RAND_127[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_50139_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_50225_addr = 5'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_50225_data = row_metadata_brob_idx[row_metadata_brob_idx_T_50225_addr]; // @[rob.scala 295:35]
  `else
  assign row_metadata_brob_idx_T_50225_data = row_metadata_brob_idx_T_50225_addr >= 5'h18 ? _RAND_128[4:0] :
    row_metadata_brob_idx[row_metadata_brob_idx_T_50225_addr]; // @[rob.scala 295:35]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx_T_23653_data = io_dis_uops_0_brob_idx;
  assign row_metadata_brob_idx_T_23653_addr = rob_tail;
  assign row_metadata_brob_idx_T_23653_mask = 1'h1;
  assign row_metadata_brob_idx_T_23653_en = new_DoPrim113799714;
  assign row_metadata_has_brorjalr_T_23664_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_23664_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_23664_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_23664_data = row_metadata_has_brorjalr_T_23664_addr >= 5'h18 ? _RAND_130[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_23664_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48249_addr = 5'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48249_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48249_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48249_data = row_metadata_has_brorjalr_T_48249_addr >= 5'h18 ? _RAND_131[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48249_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48335_addr = 5'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48335_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48335_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48335_data = row_metadata_has_brorjalr_T_48335_addr >= 5'h18 ? _RAND_132[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48335_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48421_addr = 5'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48421_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48421_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48421_data = row_metadata_has_brorjalr_T_48421_addr >= 5'h18 ? _RAND_133[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48421_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48507_addr = 5'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48507_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48507_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48507_data = row_metadata_has_brorjalr_T_48507_addr >= 5'h18 ? _RAND_134[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48507_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48593_addr = 5'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48593_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48593_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48593_data = row_metadata_has_brorjalr_T_48593_addr >= 5'h18 ? _RAND_135[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48593_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48679_addr = 5'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48679_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48679_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48679_data = row_metadata_has_brorjalr_T_48679_addr >= 5'h18 ? _RAND_136[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48679_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48765_addr = 5'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48765_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48765_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48765_data = row_metadata_has_brorjalr_T_48765_addr >= 5'h18 ? _RAND_137[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48765_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48851_addr = 5'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48851_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48851_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48851_data = row_metadata_has_brorjalr_T_48851_addr >= 5'h18 ? _RAND_138[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48851_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48937_addr = 5'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_48937_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48937_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_48937_data = row_metadata_has_brorjalr_T_48937_addr >= 5'h18 ? _RAND_139[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_48937_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49023_addr = 5'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49023_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49023_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49023_data = row_metadata_has_brorjalr_T_49023_addr >= 5'h18 ? _RAND_140[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49023_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49109_addr = 5'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49109_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49109_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49109_data = row_metadata_has_brorjalr_T_49109_addr >= 5'h18 ? _RAND_141[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49109_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49195_addr = 5'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49195_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49195_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49195_data = row_metadata_has_brorjalr_T_49195_addr >= 5'h18 ? _RAND_142[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49195_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49281_addr = 5'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49281_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49281_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49281_data = row_metadata_has_brorjalr_T_49281_addr >= 5'h18 ? _RAND_143[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49281_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49367_addr = 5'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49367_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49367_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49367_data = row_metadata_has_brorjalr_T_49367_addr >= 5'h18 ? _RAND_144[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49367_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49453_addr = 5'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49453_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49453_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49453_data = row_metadata_has_brorjalr_T_49453_addr >= 5'h18 ? _RAND_145[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49453_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49539_addr = 5'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49539_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49539_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49539_data = row_metadata_has_brorjalr_T_49539_addr >= 5'h18 ? _RAND_146[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49539_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49625_addr = 5'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49625_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49625_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49625_data = row_metadata_has_brorjalr_T_49625_addr >= 5'h18 ? _RAND_147[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49625_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49711_addr = 5'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49711_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49711_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49711_data = row_metadata_has_brorjalr_T_49711_addr >= 5'h18 ? _RAND_148[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49711_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49797_addr = 5'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49797_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49797_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49797_data = row_metadata_has_brorjalr_T_49797_addr >= 5'h18 ? _RAND_149[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49797_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49883_addr = 5'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49883_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49883_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49883_data = row_metadata_has_brorjalr_T_49883_addr >= 5'h18 ? _RAND_150[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49883_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49969_addr = 5'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_49969_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49969_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_49969_data = row_metadata_has_brorjalr_T_49969_addr >= 5'h18 ? _RAND_151[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_49969_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_50055_addr = 5'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_50055_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_50055_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_50055_data = row_metadata_has_brorjalr_T_50055_addr >= 5'h18 ? _RAND_152[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_50055_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_50141_addr = 5'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_50141_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_50141_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_50141_data = row_metadata_has_brorjalr_T_50141_addr >= 5'h18 ? _RAND_153[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_50141_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_50227_addr = 5'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_50227_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_50227_addr]; // @[rob.scala 296:38]
  `else
  assign row_metadata_has_brorjalr_T_50227_data = row_metadata_has_brorjalr_T_50227_addr >= 5'h18 ? _RAND_154[0:0] :
    row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_50227_addr]; // @[rob.scala 296:38]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr_T_23654_data = io_dis_has_br_or_jalr_in_packet;
  assign row_metadata_has_brorjalr_T_23654_addr = rob_tail;
  assign row_metadata_has_brorjalr_T_23654_mask = 1'h1;
  assign row_metadata_has_brorjalr_T_23654_en = new_DoPrim113799794;
  assign row_metadata_has_brorjalr_T_23662_data = 1'h0;
  assign row_metadata_has_brorjalr_T_23662_addr = rob_tail;
  assign row_metadata_has_brorjalr_T_23662_mask = 1'h1;
  assign row_metadata_has_brorjalr_T_23662_en = io_flush_brob;
  assign T_23710_T_29091_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_29091_data = T_23710[T_23710_T_29091_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_29091_data = T_23710_T_29091_addr >= 5'h18 ? _RAND_156[0:0] : T_23710[T_23710_T_29091_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_32866_addr = 5'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_32866_data = T_23710[T_23710_T_32866_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_32866_data = T_23710_T_32866_addr >= 5'h18 ? _RAND_157[0:0] : T_23710[T_23710_T_32866_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_32980_addr = 5'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_32980_data = T_23710[T_23710_T_32980_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_32980_data = T_23710_T_32980_addr >= 5'h18 ? _RAND_158[0:0] : T_23710[T_23710_T_32980_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33094_addr = 5'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33094_data = T_23710[T_23710_T_33094_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33094_data = T_23710_T_33094_addr >= 5'h18 ? _RAND_159[0:0] : T_23710[T_23710_T_33094_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33208_addr = 5'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33208_data = T_23710[T_23710_T_33208_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33208_data = T_23710_T_33208_addr >= 5'h18 ? _RAND_160[0:0] : T_23710[T_23710_T_33208_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33322_addr = 5'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33322_data = T_23710[T_23710_T_33322_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33322_data = T_23710_T_33322_addr >= 5'h18 ? _RAND_161[0:0] : T_23710[T_23710_T_33322_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33436_addr = 5'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33436_data = T_23710[T_23710_T_33436_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33436_data = T_23710_T_33436_addr >= 5'h18 ? _RAND_162[0:0] : T_23710[T_23710_T_33436_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33550_addr = 5'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33550_data = T_23710[T_23710_T_33550_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33550_data = T_23710_T_33550_addr >= 5'h18 ? _RAND_163[0:0] : T_23710[T_23710_T_33550_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33664_addr = 5'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33664_data = T_23710[T_23710_T_33664_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33664_data = T_23710_T_33664_addr >= 5'h18 ? _RAND_164[0:0] : T_23710[T_23710_T_33664_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33778_addr = 5'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33778_data = T_23710[T_23710_T_33778_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33778_data = T_23710_T_33778_addr >= 5'h18 ? _RAND_165[0:0] : T_23710[T_23710_T_33778_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33892_addr = 5'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_33892_data = T_23710[T_23710_T_33892_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_33892_data = T_23710_T_33892_addr >= 5'h18 ? _RAND_166[0:0] : T_23710[T_23710_T_33892_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34006_addr = 5'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34006_data = T_23710[T_23710_T_34006_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34006_data = T_23710_T_34006_addr >= 5'h18 ? _RAND_167[0:0] : T_23710[T_23710_T_34006_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34120_addr = 5'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34120_data = T_23710[T_23710_T_34120_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34120_data = T_23710_T_34120_addr >= 5'h18 ? _RAND_168[0:0] : T_23710[T_23710_T_34120_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34234_addr = 5'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34234_data = T_23710[T_23710_T_34234_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34234_data = T_23710_T_34234_addr >= 5'h18 ? _RAND_169[0:0] : T_23710[T_23710_T_34234_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34348_addr = 5'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34348_data = T_23710[T_23710_T_34348_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34348_data = T_23710_T_34348_addr >= 5'h18 ? _RAND_170[0:0] : T_23710[T_23710_T_34348_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34462_addr = 5'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34462_data = T_23710[T_23710_T_34462_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34462_data = T_23710_T_34462_addr >= 5'h18 ? _RAND_171[0:0] : T_23710[T_23710_T_34462_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34576_addr = 5'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34576_data = T_23710[T_23710_T_34576_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34576_data = T_23710_T_34576_addr >= 5'h18 ? _RAND_172[0:0] : T_23710[T_23710_T_34576_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34690_addr = 5'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34690_data = T_23710[T_23710_T_34690_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34690_data = T_23710_T_34690_addr >= 5'h18 ? _RAND_173[0:0] : T_23710[T_23710_T_34690_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34804_addr = 5'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34804_data = T_23710[T_23710_T_34804_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34804_data = T_23710_T_34804_addr >= 5'h18 ? _RAND_174[0:0] : T_23710[T_23710_T_34804_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34918_addr = 5'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_34918_data = T_23710[T_23710_T_34918_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_34918_data = T_23710_T_34918_addr >= 5'h18 ? _RAND_175[0:0] : T_23710[T_23710_T_34918_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35032_addr = 5'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35032_data = T_23710[T_23710_T_35032_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_35032_data = T_23710_T_35032_addr >= 5'h18 ? _RAND_176[0:0] : T_23710[T_23710_T_35032_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35146_addr = 5'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35146_data = T_23710[T_23710_T_35146_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_35146_data = T_23710_T_35146_addr >= 5'h18 ? _RAND_177[0:0] : T_23710[T_23710_T_35146_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35260_addr = 5'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35260_data = T_23710[T_23710_T_35260_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_35260_data = T_23710_T_35260_addr >= 5'h18 ? _RAND_178[0:0] : T_23710[T_23710_T_35260_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35374_addr = 5'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35374_data = T_23710[T_23710_T_35374_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_35374_data = T_23710_T_35374_addr >= 5'h18 ? _RAND_179[0:0] : T_23710[T_23710_T_35374_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35488_addr = 5'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_35488_data = T_23710[T_23710_T_35488_addr]; // @[rob.scala 335:30]
  `else
  assign T_23710_T_35488_data = T_23710_T_35488_addr >= 5'h18 ? _RAND_180[0:0] : T_23710[T_23710_T_35488_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_23710_T_28316_data = new_DoPrim113799882;
  assign T_23710_T_28316_addr = rob_tail;
  assign T_23710_T_28316_mask = 1'h1;
  assign T_23710_T_28316_en = io_dis_valids_0;
  assign T_23710_T_28594_data = 1'h0;
  assign T_23710_T_28594_addr = new_DoPrim113799885;
  assign T_23710_T_28594_mask = 1'h1;
  assign T_23710_T_28594_en = new_DoPrim113799884;
  assign T_23710_T_28602_data = 1'h0;
  assign T_23710_T_28602_addr = new_DoPrim113799890;
  assign T_23710_T_28602_mask = 1'h1;
  assign T_23710_T_28602_en = new_DoPrim113799889;
  assign T_23710_T_28610_data = 1'h0;
  assign T_23710_T_28610_addr = new_DoPrim113799895;
  assign T_23710_T_28610_mask = 1'h1;
  assign T_23710_T_28610_en = new_DoPrim113799894;
  assign T_23710_T_28618_data = 1'h0;
  assign T_23710_T_28618_addr = new_DoPrim113799900;
  assign T_23710_T_28618_mask = 1'h1;
  assign T_23710_T_28618_en = new_DoPrim113799899;
  assign T_28311_T_29089_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_29089_data = T_28311[T_28311_T_29089_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_29089_data = T_28311_T_29089_addr >= 5'h18 ? _RAND_182[0:0] : T_28311[T_28311_T_29089_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_32978_addr = 5'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_32978_data = T_28311[T_28311_T_32978_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_32978_data = T_28311_T_32978_addr >= 5'h18 ? _RAND_183[0:0] : T_28311[T_28311_T_32978_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33092_addr = 5'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33092_data = T_28311[T_28311_T_33092_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33092_data = T_28311_T_33092_addr >= 5'h18 ? _RAND_184[0:0] : T_28311[T_28311_T_33092_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33206_addr = 5'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33206_data = T_28311[T_28311_T_33206_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33206_data = T_28311_T_33206_addr >= 5'h18 ? _RAND_185[0:0] : T_28311[T_28311_T_33206_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33320_addr = 5'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33320_data = T_28311[T_28311_T_33320_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33320_data = T_28311_T_33320_addr >= 5'h18 ? _RAND_186[0:0] : T_28311[T_28311_T_33320_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33434_addr = 5'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33434_data = T_28311[T_28311_T_33434_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33434_data = T_28311_T_33434_addr >= 5'h18 ? _RAND_187[0:0] : T_28311[T_28311_T_33434_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33548_addr = 5'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33548_data = T_28311[T_28311_T_33548_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33548_data = T_28311_T_33548_addr >= 5'h18 ? _RAND_188[0:0] : T_28311[T_28311_T_33548_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33662_addr = 5'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33662_data = T_28311[T_28311_T_33662_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33662_data = T_28311_T_33662_addr >= 5'h18 ? _RAND_189[0:0] : T_28311[T_28311_T_33662_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33776_addr = 5'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33776_data = T_28311[T_28311_T_33776_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33776_data = T_28311_T_33776_addr >= 5'h18 ? _RAND_190[0:0] : T_28311[T_28311_T_33776_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33890_addr = 5'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_33890_data = T_28311[T_28311_T_33890_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_33890_data = T_28311_T_33890_addr >= 5'h18 ? _RAND_191[0:0] : T_28311[T_28311_T_33890_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34004_addr = 5'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34004_data = T_28311[T_28311_T_34004_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34004_data = T_28311_T_34004_addr >= 5'h18 ? _RAND_192[0:0] : T_28311[T_28311_T_34004_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34118_addr = 5'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34118_data = T_28311[T_28311_T_34118_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34118_data = T_28311_T_34118_addr >= 5'h18 ? _RAND_193[0:0] : T_28311[T_28311_T_34118_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34232_addr = 5'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34232_data = T_28311[T_28311_T_34232_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34232_data = T_28311_T_34232_addr >= 5'h18 ? _RAND_194[0:0] : T_28311[T_28311_T_34232_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34346_addr = 5'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34346_data = T_28311[T_28311_T_34346_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34346_data = T_28311_T_34346_addr >= 5'h18 ? _RAND_195[0:0] : T_28311[T_28311_T_34346_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34460_addr = 5'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34460_data = T_28311[T_28311_T_34460_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34460_data = T_28311_T_34460_addr >= 5'h18 ? _RAND_196[0:0] : T_28311[T_28311_T_34460_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34574_addr = 5'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34574_data = T_28311[T_28311_T_34574_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34574_data = T_28311_T_34574_addr >= 5'h18 ? _RAND_197[0:0] : T_28311[T_28311_T_34574_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34688_addr = 5'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34688_data = T_28311[T_28311_T_34688_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34688_data = T_28311_T_34688_addr >= 5'h18 ? _RAND_198[0:0] : T_28311[T_28311_T_34688_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34802_addr = 5'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34802_data = T_28311[T_28311_T_34802_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34802_data = T_28311_T_34802_addr >= 5'h18 ? _RAND_199[0:0] : T_28311[T_28311_T_34802_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34916_addr = 5'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_34916_data = T_28311[T_28311_T_34916_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_34916_data = T_28311_T_34916_addr >= 5'h18 ? _RAND_200[0:0] : T_28311[T_28311_T_34916_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35030_addr = 5'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35030_data = T_28311[T_28311_T_35030_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_35030_data = T_28311_T_35030_addr >= 5'h18 ? _RAND_201[0:0] : T_28311[T_28311_T_35030_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35144_addr = 5'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35144_data = T_28311[T_28311_T_35144_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_35144_data = T_28311_T_35144_addr >= 5'h18 ? _RAND_202[0:0] : T_28311[T_28311_T_35144_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35258_addr = 5'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35258_data = T_28311[T_28311_T_35258_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_35258_data = T_28311_T_35258_addr >= 5'h18 ? _RAND_203[0:0] : T_28311[T_28311_T_35258_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35372_addr = 5'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35372_data = T_28311[T_28311_T_35372_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_35372_data = T_28311_T_35372_addr >= 5'h18 ? _RAND_204[0:0] : T_28311[T_28311_T_35372_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35486_addr = 5'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35486_data = T_28311[T_28311_T_35486_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_35486_data = T_28311_T_35486_addr >= 5'h18 ? _RAND_205[0:0] : T_28311[T_28311_T_35486_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35600_addr = 5'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_35600_data = T_28311[T_28311_T_35600_addr]; // @[rob.scala 339:30]
  `else
  assign T_28311_T_35600_data = T_28311_T_35600_addr >= 5'h18 ? _RAND_206[0:0] : T_28311[T_28311_T_35600_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28311_T_28407_data = io_dis_uops_0_exception;
  assign T_28311_T_28407_addr = rob_tail;
  assign T_28311_T_28407_mask = 1'h1;
  assign T_28311_T_28407_en = io_dis_valids_0;
  assign T_28311_T_29079_data = 1'h1;
  assign T_28311_T_29079_addr = new_DoPrim113799985;
  assign T_28311_T_29079_mask = 1'h1;
  assign T_28311_T_29079_en = new_DoPrim113799984;
  assign T_28311_T_29087_data = 1'h1;
  assign T_28311_T_29087_addr = new_DoPrim113799990;
  assign T_28311_T_29087_mask = 1'h1;
  assign T_28311_T_29087_en = new_DoPrim113799989;
  assign T_28311_T_29363_data = 1'h0;
  assign T_28311_T_29363_addr = T_29097 ? rob_tail : rob_head;
  assign T_28311_T_29363_mask = 1'h1;
  assign T_28311_T_29363_en = new_DoPrim113799994;
  assign T_28314_T_31814_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_28314_T_31814_data = T_28314[T_28314_T_31814_addr]; // @[rob.scala 340:30]
  `else
  assign T_28314_T_31814_data = T_28314_T_31814_addr >= 5'h18 ? _RAND_208[4:0] : T_28314[T_28314_T_31814_addr]; // @[rob.scala 340:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_28314_T_28408_data = 5'h0;
  assign T_28314_T_28408_addr = rob_tail;
  assign T_28314_T_28408_mask = 1'h1;
  assign T_28314_T_28408_en = io_dis_valids_0;
  assign T_28314_T_29065_data = io_fflags_0_bits_flags;
  assign T_28314_T_29065_addr = new_DoPrim113828225;
  assign T_28314_T_29065_mask = 1'h1;
  assign T_28314_T_29065_en = new_DoPrim113828224;
  assign T_28314_T_29072_data = io_fflags_1_bits_flags;
  assign T_28314_T_29072_addr = new_DoPrim113828230;
  assign T_28314_T_29072_mask = 1'h1;
  assign T_28314_T_29072_en = new_DoPrim113828229;
  assign T_35638_T_41019_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_41019_data = T_35638[T_35638_T_41019_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_41019_data = T_35638_T_41019_addr >= 5'h18 ? _RAND_210[0:0] : T_35638[T_35638_T_41019_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_44794_addr = 5'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_44794_data = T_35638[T_35638_T_44794_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_44794_data = T_35638_T_44794_addr >= 5'h18 ? _RAND_211[0:0] : T_35638[T_35638_T_44794_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_44908_addr = 5'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_44908_data = T_35638[T_35638_T_44908_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_44908_data = T_35638_T_44908_addr >= 5'h18 ? _RAND_212[0:0] : T_35638[T_35638_T_44908_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45022_addr = 5'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45022_data = T_35638[T_35638_T_45022_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45022_data = T_35638_T_45022_addr >= 5'h18 ? _RAND_213[0:0] : T_35638[T_35638_T_45022_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45136_addr = 5'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45136_data = T_35638[T_35638_T_45136_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45136_data = T_35638_T_45136_addr >= 5'h18 ? _RAND_214[0:0] : T_35638[T_35638_T_45136_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45250_addr = 5'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45250_data = T_35638[T_35638_T_45250_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45250_data = T_35638_T_45250_addr >= 5'h18 ? _RAND_215[0:0] : T_35638[T_35638_T_45250_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45364_addr = 5'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45364_data = T_35638[T_35638_T_45364_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45364_data = T_35638_T_45364_addr >= 5'h18 ? _RAND_216[0:0] : T_35638[T_35638_T_45364_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45478_addr = 5'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45478_data = T_35638[T_35638_T_45478_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45478_data = T_35638_T_45478_addr >= 5'h18 ? _RAND_217[0:0] : T_35638[T_35638_T_45478_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45592_addr = 5'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45592_data = T_35638[T_35638_T_45592_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45592_data = T_35638_T_45592_addr >= 5'h18 ? _RAND_218[0:0] : T_35638[T_35638_T_45592_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45706_addr = 5'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45706_data = T_35638[T_35638_T_45706_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45706_data = T_35638_T_45706_addr >= 5'h18 ? _RAND_219[0:0] : T_35638[T_35638_T_45706_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45820_addr = 5'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45820_data = T_35638[T_35638_T_45820_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45820_data = T_35638_T_45820_addr >= 5'h18 ? _RAND_220[0:0] : T_35638[T_35638_T_45820_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45934_addr = 5'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_45934_data = T_35638[T_35638_T_45934_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_45934_data = T_35638_T_45934_addr >= 5'h18 ? _RAND_221[0:0] : T_35638[T_35638_T_45934_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46048_addr = 5'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46048_data = T_35638[T_35638_T_46048_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46048_data = T_35638_T_46048_addr >= 5'h18 ? _RAND_222[0:0] : T_35638[T_35638_T_46048_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46162_addr = 5'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46162_data = T_35638[T_35638_T_46162_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46162_data = T_35638_T_46162_addr >= 5'h18 ? _RAND_223[0:0] : T_35638[T_35638_T_46162_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46276_addr = 5'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46276_data = T_35638[T_35638_T_46276_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46276_data = T_35638_T_46276_addr >= 5'h18 ? _RAND_224[0:0] : T_35638[T_35638_T_46276_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46390_addr = 5'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46390_data = T_35638[T_35638_T_46390_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46390_data = T_35638_T_46390_addr >= 5'h18 ? _RAND_225[0:0] : T_35638[T_35638_T_46390_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46504_addr = 5'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46504_data = T_35638[T_35638_T_46504_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46504_data = T_35638_T_46504_addr >= 5'h18 ? _RAND_226[0:0] : T_35638[T_35638_T_46504_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46618_addr = 5'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46618_data = T_35638[T_35638_T_46618_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46618_data = T_35638_T_46618_addr >= 5'h18 ? _RAND_227[0:0] : T_35638[T_35638_T_46618_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46732_addr = 5'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46732_data = T_35638[T_35638_T_46732_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46732_data = T_35638_T_46732_addr >= 5'h18 ? _RAND_228[0:0] : T_35638[T_35638_T_46732_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46846_addr = 5'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46846_data = T_35638[T_35638_T_46846_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46846_data = T_35638_T_46846_addr >= 5'h18 ? _RAND_229[0:0] : T_35638[T_35638_T_46846_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46960_addr = 5'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_46960_data = T_35638[T_35638_T_46960_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_46960_data = T_35638_T_46960_addr >= 5'h18 ? _RAND_230[0:0] : T_35638[T_35638_T_46960_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47074_addr = 5'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47074_data = T_35638[T_35638_T_47074_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_47074_data = T_35638_T_47074_addr >= 5'h18 ? _RAND_231[0:0] : T_35638[T_35638_T_47074_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47188_addr = 5'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47188_data = T_35638[T_35638_T_47188_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_47188_data = T_35638_T_47188_addr >= 5'h18 ? _RAND_232[0:0] : T_35638[T_35638_T_47188_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47302_addr = 5'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47302_data = T_35638[T_35638_T_47302_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_47302_data = T_35638_T_47302_addr >= 5'h18 ? _RAND_233[0:0] : T_35638[T_35638_T_47302_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47416_addr = 5'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_47416_data = T_35638[T_35638_T_47416_addr]; // @[rob.scala 335:30]
  `else
  assign T_35638_T_47416_data = T_35638_T_47416_addr >= 5'h18 ? _RAND_234[0:0] : T_35638[T_35638_T_47416_addr]; // @[rob.scala 335:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_35638_T_40244_data = new_DoPrim113828312;
  assign T_35638_T_40244_addr = rob_tail;
  assign T_35638_T_40244_mask = 1'h1;
  assign T_35638_T_40244_en = io_dis_valids_1;
  assign T_35638_T_40522_data = 1'h0;
  assign T_35638_T_40522_addr = new_DoPrim113828315;
  assign T_35638_T_40522_mask = 1'h1;
  assign T_35638_T_40522_en = new_DoPrim113828314;
  assign T_35638_T_40530_data = 1'h0;
  assign T_35638_T_40530_addr = new_DoPrim113828320;
  assign T_35638_T_40530_mask = 1'h1;
  assign T_35638_T_40530_en = new_DoPrim113828319;
  assign T_35638_T_40538_data = 1'h0;
  assign T_35638_T_40538_addr = new_DoPrim113828325;
  assign T_35638_T_40538_mask = 1'h1;
  assign T_35638_T_40538_en = new_DoPrim113828324;
  assign T_35638_T_40546_data = 1'h0;
  assign T_35638_T_40546_addr = new_DoPrim113828330;
  assign T_35638_T_40546_mask = 1'h1;
  assign T_35638_T_40546_en = new_DoPrim113828329;
  assign T_40239_T_41017_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_41017_data = T_40239[T_40239_T_41017_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_41017_data = T_40239_T_41017_addr >= 5'h18 ? _RAND_236[0:0] : T_40239[T_40239_T_41017_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_44906_addr = 5'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_44906_data = T_40239[T_40239_T_44906_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_44906_data = T_40239_T_44906_addr >= 5'h18 ? _RAND_237[0:0] : T_40239[T_40239_T_44906_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45020_addr = 5'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45020_data = T_40239[T_40239_T_45020_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45020_data = T_40239_T_45020_addr >= 5'h18 ? _RAND_238[0:0] : T_40239[T_40239_T_45020_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45134_addr = 5'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45134_data = T_40239[T_40239_T_45134_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45134_data = T_40239_T_45134_addr >= 5'h18 ? _RAND_239[0:0] : T_40239[T_40239_T_45134_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45248_addr = 5'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45248_data = T_40239[T_40239_T_45248_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45248_data = T_40239_T_45248_addr >= 5'h18 ? _RAND_240[0:0] : T_40239[T_40239_T_45248_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45362_addr = 5'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45362_data = T_40239[T_40239_T_45362_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45362_data = T_40239_T_45362_addr >= 5'h18 ? _RAND_241[0:0] : T_40239[T_40239_T_45362_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45476_addr = 5'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45476_data = T_40239[T_40239_T_45476_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45476_data = T_40239_T_45476_addr >= 5'h18 ? _RAND_242[0:0] : T_40239[T_40239_T_45476_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45590_addr = 5'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45590_data = T_40239[T_40239_T_45590_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45590_data = T_40239_T_45590_addr >= 5'h18 ? _RAND_243[0:0] : T_40239[T_40239_T_45590_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45704_addr = 5'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45704_data = T_40239[T_40239_T_45704_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45704_data = T_40239_T_45704_addr >= 5'h18 ? _RAND_244[0:0] : T_40239[T_40239_T_45704_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45818_addr = 5'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45818_data = T_40239[T_40239_T_45818_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45818_data = T_40239_T_45818_addr >= 5'h18 ? _RAND_245[0:0] : T_40239[T_40239_T_45818_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45932_addr = 5'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_45932_data = T_40239[T_40239_T_45932_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_45932_data = T_40239_T_45932_addr >= 5'h18 ? _RAND_246[0:0] : T_40239[T_40239_T_45932_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46046_addr = 5'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46046_data = T_40239[T_40239_T_46046_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46046_data = T_40239_T_46046_addr >= 5'h18 ? _RAND_247[0:0] : T_40239[T_40239_T_46046_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46160_addr = 5'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46160_data = T_40239[T_40239_T_46160_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46160_data = T_40239_T_46160_addr >= 5'h18 ? _RAND_248[0:0] : T_40239[T_40239_T_46160_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46274_addr = 5'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46274_data = T_40239[T_40239_T_46274_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46274_data = T_40239_T_46274_addr >= 5'h18 ? _RAND_249[0:0] : T_40239[T_40239_T_46274_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46388_addr = 5'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46388_data = T_40239[T_40239_T_46388_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46388_data = T_40239_T_46388_addr >= 5'h18 ? _RAND_250[0:0] : T_40239[T_40239_T_46388_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46502_addr = 5'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46502_data = T_40239[T_40239_T_46502_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46502_data = T_40239_T_46502_addr >= 5'h18 ? _RAND_251[0:0] : T_40239[T_40239_T_46502_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46616_addr = 5'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46616_data = T_40239[T_40239_T_46616_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46616_data = T_40239_T_46616_addr >= 5'h18 ? _RAND_252[0:0] : T_40239[T_40239_T_46616_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46730_addr = 5'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46730_data = T_40239[T_40239_T_46730_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46730_data = T_40239_T_46730_addr >= 5'h18 ? _RAND_253[0:0] : T_40239[T_40239_T_46730_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46844_addr = 5'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46844_data = T_40239[T_40239_T_46844_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46844_data = T_40239_T_46844_addr >= 5'h18 ? _RAND_254[0:0] : T_40239[T_40239_T_46844_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46958_addr = 5'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_46958_data = T_40239[T_40239_T_46958_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_46958_data = T_40239_T_46958_addr >= 5'h18 ? _RAND_255[0:0] : T_40239[T_40239_T_46958_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47072_addr = 5'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47072_data = T_40239[T_40239_T_47072_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_47072_data = T_40239_T_47072_addr >= 5'h18 ? _RAND_256[0:0] : T_40239[T_40239_T_47072_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47186_addr = 5'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47186_data = T_40239[T_40239_T_47186_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_47186_data = T_40239_T_47186_addr >= 5'h18 ? _RAND_257[0:0] : T_40239[T_40239_T_47186_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47300_addr = 5'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47300_data = T_40239[T_40239_T_47300_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_47300_data = T_40239_T_47300_addr >= 5'h18 ? _RAND_258[0:0] : T_40239[T_40239_T_47300_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47414_addr = 5'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47414_data = T_40239[T_40239_T_47414_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_47414_data = T_40239_T_47414_addr >= 5'h18 ? _RAND_259[0:0] : T_40239[T_40239_T_47414_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47528_addr = 5'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_47528_data = T_40239[T_40239_T_47528_addr]; // @[rob.scala 339:30]
  `else
  assign T_40239_T_47528_data = T_40239_T_47528_addr >= 5'h18 ? _RAND_260[0:0] : T_40239[T_40239_T_47528_addr]; // @[rob.scala 339:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40239_T_40335_data = io_dis_uops_1_exception;
  assign T_40239_T_40335_addr = rob_tail;
  assign T_40239_T_40335_mask = 1'h1;
  assign T_40239_T_40335_en = io_dis_valids_1;
  assign T_40239_T_41007_data = 1'h1;
  assign T_40239_T_41007_addr = new_DoPrim113828415;
  assign T_40239_T_41007_mask = 1'h1;
  assign T_40239_T_41007_en = new_DoPrim113828414;
  assign T_40239_T_41015_data = 1'h1;
  assign T_40239_T_41015_addr = new_DoPrim113828420;
  assign T_40239_T_41015_mask = 1'h1;
  assign T_40239_T_41015_en = new_DoPrim113828419;
  assign T_40239_T_41291_data = 1'h0;
  assign T_40239_T_41291_addr = T_29097 ? rob_tail : rob_head;
  assign T_40239_T_41291_mask = 1'h1;
  assign T_40239_T_41291_en = new_DoPrim113828424;
  assign T_40242_T_43742_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_40242_T_43742_data = T_40242[T_40242_T_43742_addr]; // @[rob.scala 340:30]
  `else
  assign T_40242_T_43742_data = T_40242_T_43742_addr >= 5'h18 ? _RAND_262[4:0] : T_40242[T_40242_T_43742_addr]; // @[rob.scala 340:30]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign T_40242_T_40336_data = 5'h0;
  assign T_40242_T_40336_addr = rob_tail;
  assign T_40242_T_40336_mask = 1'h1;
  assign T_40242_T_40336_en = io_dis_valids_1;
  assign T_40242_T_40993_data = io_fflags_0_bits_flags;
  assign T_40242_T_40993_addr = new_DoPrim113856655;
  assign T_40242_T_40993_mask = 1'h1;
  assign T_40242_T_40993_en = new_DoPrim113856654;
  assign T_40242_T_41000_data = io_fflags_1_bits_flags;
  assign T_40242_T_41000_addr = new_DoPrim113856660;
  assign T_40242_T_41000_mask = 1'h1;
  assign T_40242_T_41000_en = new_DoPrim113856659;
  assign io_curr_rob_tail = new_DoPrim0; // @[rob.scala 761:21]
  assign io_com_valids_0 = new_DoPrim1; // @[rob.scala 585:72]
  assign io_com_valids_1 = new_DoPrim2; // @[rob.scala 585:72]
  assign io_com_uops_0_valid = 5'h17 == T_29096 ? T_26182_23_valid : _GEN_5971; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_iw_state = 5'h17 == T_29096 ? T_26182_23_iw_state : _GEN_5972; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_uopc = 5'h17 == T_29096 ? T_26182_23_uopc : _GEN_5973; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_inst = 5'h17 == T_29096 ? T_26182_23_inst : _GEN_5974; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_pc = 5'h17 == T_29096 ? T_26182_23_pc : _GEN_5975; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_fu_code = 5'h17 == T_29096 ? T_26182_23_fu_code : _GEN_5976; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_br_type = 5'h17 == T_29096 ? T_26182_23_ctrl_br_type : _GEN_5977; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_op1_sel = 5'h17 == T_29096 ? T_26182_23_ctrl_op1_sel : _GEN_5978; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_op2_sel = 5'h17 == T_29096 ? T_26182_23_ctrl_op2_sel : _GEN_5979; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_imm_sel = 5'h17 == T_29096 ? T_26182_23_ctrl_imm_sel : _GEN_5980; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_op_fcn = 5'h17 == T_29096 ? T_26182_23_ctrl_op_fcn : _GEN_5981; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_fcn_dw = 5'h17 == T_29096 ? T_26182_23_ctrl_fcn_dw : _GEN_5982; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_rf_wen = 5'h17 == T_29096 ? T_26182_23_ctrl_rf_wen : _GEN_5983; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_csr_cmd = 5'h17 == T_29096 ? T_26182_23_ctrl_csr_cmd : _GEN_5984; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_is_load = 5'h17 == T_29096 ? T_26182_23_ctrl_is_load : _GEN_5985; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_is_sta = 5'h17 == T_29096 ? T_26182_23_ctrl_is_sta : _GEN_5986; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ctrl_is_std = 5'h17 == T_29096 ? T_26182_23_ctrl_is_std : _GEN_5987; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_wakeup_delay = 5'h17 == T_29096 ? T_26182_23_wakeup_delay : _GEN_5988; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_allocate_brtag = 5'h17 == T_29096 ? T_26182_23_allocate_brtag : _GEN_5989; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_br_or_jmp = 5'h17 == T_29096 ? T_26182_23_is_br_or_jmp : _GEN_5990; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_jump = 5'h17 == T_29096 ? T_26182_23_is_jump : _GEN_5991; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_jal = 5'h17 == T_29096 ? T_26182_23_is_jal : _GEN_5992; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_ret = 5'h17 == T_29096 ? T_26182_23_is_ret : _GEN_5993; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_call = 5'h17 == T_29096 ? T_26182_23_is_call : _GEN_5994; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_mask = 5'h17 == T_29096 ? T_26182_23_br_mask : _GEN_5995; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_tag = 5'h17 == T_29096 ? T_26182_23_br_tag : _GEN_5996; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_prediction_bpd_predict_val = 5'h17 == T_29096 ? T_26182_23_br_prediction_bpd_predict_val :
    _GEN_5997; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_prediction_bpd_predict_taken = 5'h17 == T_29096 ? T_26182_23_br_prediction_bpd_predict_taken
     : _GEN_5998; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_prediction_btb_hit = 5'h17 == T_29096 ? T_26182_23_br_prediction_btb_hit : _GEN_5999; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_prediction_btb_predicted = 5'h17 == T_29096 ? T_26182_23_br_prediction_btb_predicted :
    _GEN_6000; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_br_prediction_is_br_or_jalr = 5'h17 == T_29096 ? T_26182_23_br_prediction_is_br_or_jalr :
    _GEN_6001; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stat_brjmp_mispredicted = 5'h17 == T_29096 ? T_26182_23_stat_brjmp_mispredicted : _GEN_6002; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stat_btb_made_pred = 5'h17 == T_29096 ? T_26182_23_stat_btb_made_pred : _GEN_6003; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stat_btb_mispredicted = 5'h17 == T_29096 ? T_26182_23_stat_btb_mispredicted : _GEN_6004; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stat_bpd_made_pred = 5'h17 == T_29096 ? T_26182_23_stat_bpd_made_pred : _GEN_6005; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stat_bpd_mispredicted = 5'h17 == T_29096 ? T_26182_23_stat_bpd_mispredicted : _GEN_6006; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_fetch_pc_lob = 5'h17 == T_29096 ? T_26182_23_fetch_pc_lob : _GEN_6007; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_imm_packed = 5'h17 == T_29096 ? T_26182_23_imm_packed : _GEN_6008; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_csr_addr = 5'h17 == T_29096 ? T_26182_23_csr_addr : _GEN_6009; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_rob_idx = 5'h17 == T_29096 ? T_26182_23_rob_idx : _GEN_6010; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ldq_idx = 5'h17 == T_29096 ? T_26182_23_ldq_idx : _GEN_6011; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stq_idx = 5'h17 == T_29096 ? T_26182_23_stq_idx : _GEN_6012; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_brob_idx = 5'h17 == T_29096 ? T_26182_23_brob_idx : _GEN_6013; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_pdst = 5'h17 == T_29096 ? T_26182_23_pdst : _GEN_6014; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_pop1 = 5'h17 == T_29096 ? T_26182_23_pop1 : _GEN_6015; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_pop2 = 5'h17 == T_29096 ? T_26182_23_pop2 : _GEN_6016; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_pop3 = 5'h17 == T_29096 ? T_26182_23_pop3 : _GEN_6017; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_prs1_busy = 5'h17 == T_29096 ? T_26182_23_prs1_busy : _GEN_6018; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_prs2_busy = 5'h17 == T_29096 ? T_26182_23_prs2_busy : _GEN_6019; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_prs3_busy = 5'h17 == T_29096 ? T_26182_23_prs3_busy : _GEN_6020; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_stale_pdst = 5'h17 == T_29096 ? T_26182_23_stale_pdst : _GEN_6021; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_exception = 5'h17 == T_29096 ? T_26182_23_exception : _GEN_6022; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_exc_cause = 5'h17 == T_29096 ? T_26182_23_exc_cause : _GEN_6023; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_bypassable = 5'h17 == T_29096 ? T_26182_23_bypassable : _GEN_6024; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_mem_cmd = 5'h17 == T_29096 ? T_26182_23_mem_cmd : _GEN_6025; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_mem_typ = 5'h17 == T_29096 ? T_26182_23_mem_typ : _GEN_6026; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_fence = 5'h17 == T_29096 ? T_26182_23_is_fence : _GEN_6027; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_fencei = 5'h17 == T_29096 ? T_26182_23_is_fencei : _GEN_6028; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_store = 5'h17 == T_29096 ? T_26182_23_is_store : _GEN_6029; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_amo = 5'h17 == T_29096 ? T_26182_23_is_amo : _GEN_6030; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_load = 5'h17 == T_29096 ? T_26182_23_is_load : _GEN_6031; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_is_unique = 5'h17 == T_29096 ? T_26182_23_is_unique : _GEN_6032; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_flush_on_commit = 5'h17 == T_29096 ? T_26182_23_flush_on_commit : _GEN_6033; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ldst = 5'h17 == T_29096 ? T_26182_23_ldst : _GEN_6034; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_lrs1 = 5'h17 == T_29096 ? T_26182_23_lrs1 : _GEN_6035; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_lrs2 = 5'h17 == T_29096 ? T_26182_23_lrs2 : _GEN_6036; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_lrs3 = 5'h17 == T_29096 ? T_26182_23_lrs3 : _GEN_6037; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_ldst_val = 5'h17 == T_29096 ? T_26182_23_ldst_val : _GEN_6038; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_dst_rtype = 5'h17 == T_29096 ? T_26182_23_dst_rtype : _GEN_6039; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_lrs1_rtype = 5'h17 == T_29096 ? T_26182_23_lrs1_rtype : _GEN_6040; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_lrs2_rtype = 5'h17 == T_29096 ? T_26182_23_lrs2_rtype : _GEN_6041; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_frs3_en = 5'h17 == T_29096 ? T_26182_23_frs3_en : _GEN_6042; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_fp_val = 5'h17 == T_29096 ? T_26182_23_fp_val : _GEN_6043; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_fp_single = 5'h17 == T_29096 ? T_26182_23_fp_single : _GEN_6044; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_xcpt_if = 5'h17 == T_29096 ? T_26182_23_xcpt_if : _GEN_6045; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_replay_if = 5'h17 == T_29096 ? T_26182_23_replay_if : _GEN_6046; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_0_debug_wdata = 5'h17 == rob_head ? T_26182_23_debug_wdata : _GEN_8092; // @[rob.scala 507:28 rob.scala 507:28]
  assign io_com_uops_0_debug_events_fetch_seq = 5'h17 == T_29096 ? T_26182_23_debug_events_fetch_seq : _GEN_6048; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_valid = 5'h17 == T_29096 ? T_38110_23_valid : _GEN_20114; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_iw_state = 5'h17 == T_29096 ? T_38110_23_iw_state : _GEN_20115; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_uopc = 5'h17 == T_29096 ? T_38110_23_uopc : _GEN_20116; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_inst = 5'h17 == T_29096 ? T_38110_23_inst : _GEN_20117; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_pc = 5'h17 == T_29096 ? T_38110_23_pc : _GEN_20118; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_fu_code = 5'h17 == T_29096 ? T_38110_23_fu_code : _GEN_20119; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_br_type = 5'h17 == T_29096 ? T_38110_23_ctrl_br_type : _GEN_20120; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_op1_sel = 5'h17 == T_29096 ? T_38110_23_ctrl_op1_sel : _GEN_20121; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_op2_sel = 5'h17 == T_29096 ? T_38110_23_ctrl_op2_sel : _GEN_20122; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_imm_sel = 5'h17 == T_29096 ? T_38110_23_ctrl_imm_sel : _GEN_20123; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_op_fcn = 5'h17 == T_29096 ? T_38110_23_ctrl_op_fcn : _GEN_20124; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_fcn_dw = 5'h17 == T_29096 ? T_38110_23_ctrl_fcn_dw : _GEN_20125; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_rf_wen = 5'h17 == T_29096 ? T_38110_23_ctrl_rf_wen : _GEN_20126; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_csr_cmd = 5'h17 == T_29096 ? T_38110_23_ctrl_csr_cmd : _GEN_20127; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_is_load = 5'h17 == T_29096 ? T_38110_23_ctrl_is_load : _GEN_20128; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_is_sta = 5'h17 == T_29096 ? T_38110_23_ctrl_is_sta : _GEN_20129; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ctrl_is_std = 5'h17 == T_29096 ? T_38110_23_ctrl_is_std : _GEN_20130; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_wakeup_delay = 5'h17 == T_29096 ? T_38110_23_wakeup_delay : _GEN_20131; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_allocate_brtag = 5'h17 == T_29096 ? T_38110_23_allocate_brtag : _GEN_20132; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_br_or_jmp = 5'h17 == T_29096 ? T_38110_23_is_br_or_jmp : _GEN_20133; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_jump = 5'h17 == T_29096 ? T_38110_23_is_jump : _GEN_20134; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_jal = 5'h17 == T_29096 ? T_38110_23_is_jal : _GEN_20135; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_ret = 5'h17 == T_29096 ? T_38110_23_is_ret : _GEN_20136; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_call = 5'h17 == T_29096 ? T_38110_23_is_call : _GEN_20137; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_mask = 5'h17 == T_29096 ? T_38110_23_br_mask : _GEN_20138; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_tag = 5'h17 == T_29096 ? T_38110_23_br_tag : _GEN_20139; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_prediction_bpd_predict_val = 5'h17 == T_29096 ? T_38110_23_br_prediction_bpd_predict_val :
    _GEN_20140; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_prediction_bpd_predict_taken = 5'h17 == T_29096 ? T_38110_23_br_prediction_bpd_predict_taken
     : _GEN_20141; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_prediction_btb_hit = 5'h17 == T_29096 ? T_38110_23_br_prediction_btb_hit : _GEN_20142; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_prediction_btb_predicted = 5'h17 == T_29096 ? T_38110_23_br_prediction_btb_predicted :
    _GEN_20143; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_br_prediction_is_br_or_jalr = 5'h17 == T_29096 ? T_38110_23_br_prediction_is_br_or_jalr :
    _GEN_20144; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stat_brjmp_mispredicted = 5'h17 == T_29096 ? T_38110_23_stat_brjmp_mispredicted : _GEN_20145; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stat_btb_made_pred = 5'h17 == T_29096 ? T_38110_23_stat_btb_made_pred : _GEN_20146; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stat_btb_mispredicted = 5'h17 == T_29096 ? T_38110_23_stat_btb_mispredicted : _GEN_20147; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stat_bpd_made_pred = 5'h17 == T_29096 ? T_38110_23_stat_bpd_made_pred : _GEN_20148; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stat_bpd_mispredicted = 5'h17 == T_29096 ? T_38110_23_stat_bpd_mispredicted : _GEN_20149; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_fetch_pc_lob = 5'h17 == T_29096 ? T_38110_23_fetch_pc_lob : _GEN_20150; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_imm_packed = 5'h17 == T_29096 ? T_38110_23_imm_packed : _GEN_20151; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_csr_addr = 5'h17 == T_29096 ? T_38110_23_csr_addr : _GEN_20152; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_rob_idx = 5'h17 == T_29096 ? T_38110_23_rob_idx : _GEN_20153; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ldq_idx = 5'h17 == T_29096 ? T_38110_23_ldq_idx : _GEN_20154; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stq_idx = 5'h17 == T_29096 ? T_38110_23_stq_idx : _GEN_20155; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_brob_idx = 5'h17 == T_29096 ? T_38110_23_brob_idx : _GEN_20156; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_pdst = 5'h17 == T_29096 ? T_38110_23_pdst : _GEN_20157; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_pop1 = 5'h17 == T_29096 ? T_38110_23_pop1 : _GEN_20158; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_pop2 = 5'h17 == T_29096 ? T_38110_23_pop2 : _GEN_20159; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_pop3 = 5'h17 == T_29096 ? T_38110_23_pop3 : _GEN_20160; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_prs1_busy = 5'h17 == T_29096 ? T_38110_23_prs1_busy : _GEN_20161; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_prs2_busy = 5'h17 == T_29096 ? T_38110_23_prs2_busy : _GEN_20162; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_prs3_busy = 5'h17 == T_29096 ? T_38110_23_prs3_busy : _GEN_20163; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_stale_pdst = 5'h17 == T_29096 ? T_38110_23_stale_pdst : _GEN_20164; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_exception = 5'h17 == T_29096 ? T_38110_23_exception : _GEN_20165; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_exc_cause = 5'h17 == T_29096 ? T_38110_23_exc_cause : _GEN_20166; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_bypassable = 5'h17 == T_29096 ? T_38110_23_bypassable : _GEN_20167; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_mem_cmd = 5'h17 == T_29096 ? T_38110_23_mem_cmd : _GEN_20168; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_mem_typ = 5'h17 == T_29096 ? T_38110_23_mem_typ : _GEN_20169; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_fence = 5'h17 == T_29096 ? T_38110_23_is_fence : _GEN_20170; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_fencei = 5'h17 == T_29096 ? T_38110_23_is_fencei : _GEN_20171; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_store = 5'h17 == T_29096 ? T_38110_23_is_store : _GEN_20172; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_amo = 5'h17 == T_29096 ? T_38110_23_is_amo : _GEN_20173; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_load = 5'h17 == T_29096 ? T_38110_23_is_load : _GEN_20174; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_is_unique = 5'h17 == T_29096 ? T_38110_23_is_unique : _GEN_20175; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_flush_on_commit = 5'h17 == T_29096 ? T_38110_23_flush_on_commit : _GEN_20176; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ldst = 5'h17 == T_29096 ? T_38110_23_ldst : _GEN_20177; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_lrs1 = 5'h17 == T_29096 ? T_38110_23_lrs1 : _GEN_20178; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_lrs2 = 5'h17 == T_29096 ? T_38110_23_lrs2 : _GEN_20179; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_lrs3 = 5'h17 == T_29096 ? T_38110_23_lrs3 : _GEN_20180; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_ldst_val = 5'h17 == T_29096 ? T_38110_23_ldst_val : _GEN_20181; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_dst_rtype = 5'h17 == T_29096 ? T_38110_23_dst_rtype : _GEN_20182; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_lrs1_rtype = 5'h17 == T_29096 ? T_38110_23_lrs1_rtype : _GEN_20183; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_lrs2_rtype = 5'h17 == T_29096 ? T_38110_23_lrs2_rtype : _GEN_20184; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_frs3_en = 5'h17 == T_29096 ? T_38110_23_frs3_en : _GEN_20185; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_fp_val = 5'h17 == T_29096 ? T_38110_23_fp_val : _GEN_20186; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_fp_single = 5'h17 == T_29096 ? T_38110_23_fp_single : _GEN_20187; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_xcpt_if = 5'h17 == T_29096 ? T_38110_23_xcpt_if : _GEN_20188; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_replay_if = 5'h17 == T_29096 ? T_38110_23_replay_if : _GEN_20189; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_uops_1_debug_wdata = 5'h17 == rob_head ? T_38110_23_debug_wdata : _GEN_22235; // @[rob.scala 507:28 rob.scala 507:28]
  assign io_com_uops_1_debug_events_fetch_seq = 5'h17 == T_29096 ? T_38110_23_debug_events_fetch_seq : _GEN_20191; // @[rob.scala 453:59 rob.scala 453:59]
  assign io_com_fflags_val = new_DoPrim4401855; // @[rob.scala 640:44]
  assign io_com_fflags = new_DoPrim4401856; // @[rob.scala 641:40]
  assign io_com_st_mask_0 = new_DoPrim4401857; // @[rob.scala 869:45]
  assign io_com_st_mask_1 = new_DoPrim4401858; // @[rob.scala 869:45]
  assign io_com_ld_mask_0 = new_DoPrim4401859; // @[rob.scala 870:45]
  assign io_com_ld_mask_1 = new_DoPrim4401860; // @[rob.scala 870:45]
  assign io_com_load_is_at_rob_head = T_48220 ? rob_head_is_load_1 : rob_head_is_load_0; // @[rob.scala 873:31 rob.scala 873:31]
  assign io_com_exception = new_DoPrim4430078; // @[rob.scala 596:44]
  assign io_com_exc_cause = r_xcpt_uop_exc_cause; // @[rob.scala 597:24]
  assign io_com_handling_exc = new_DoPrim4430080; // @[rob.scala 593:48]
  assign io_com_rbk_valids_0 = new_DoPrim4430081; // @[rob.scala 452:48]
  assign io_com_rbk_valids_1 = new_DoPrim4430082; // @[rob.scala 452:48]
  assign io_com_badvaddr = new_DoPrim4430083; // @[Cat.scala 20:58]
  assign io_get_pc_curr_pc = new_DoPrim4430084; // @[rob.scala 268:22]
  assign io_get_pc_curr_brob_idx = row_metadata_brob_idx_T_23669_data; // @[rob.scala 318:28]
  assign io_get_pc_next_val = new_DoPrim4430086; // @[rob.scala 279:46]
  assign io_get_pc_next_pc = new_DoPrim4430087; // @[rob.scala 280:22]
  assign io_lsu_misspec = T_47576; // @[rob.scala 601:19]
  assign io_flush_take_pc = new_DoPrim4430089; // @[rob.scala 608:37]
  assign io_flush_pc = new_DoPrim4430090; // @[rob.scala 605:17]
  assign io_flush_pipeline = T_47616; // @[rob.scala 612:22]
  assign io_flush_brob = new_DoPrim4430092; // @[rob.scala 322:61]
  assign io_empty = new_DoPrim4430093; // @[rob.scala 759:40]
  assign io_ready = new_DoPrim4430094; // @[rob.scala 764:41]
  assign io_brob_deallocate_valid = new_DoPrim4430095; // @[rob.scala 315:56]
  assign io_brob_deallocate_bits_brob_idx = row_metadata_brob_idx_T_23666_data; // @[rob.scala 316:37]
  assign io_debug_state = rob_state; // @[rob.scala 878:22]
  assign io_debug_rob_head = new_DoPrim4430098; // @[rob.scala 879:22]
  assign io_debug_xcpt_val = r_xcpt_val; // @[rob.scala 880:22]
  assign io_debug_xcpt_uop_valid = r_xcpt_uop_valid; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_iw_state = r_xcpt_uop_iw_state; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_uopc = r_xcpt_uop_uopc; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_inst = r_xcpt_uop_inst; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_pc = r_xcpt_uop_pc; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_fu_code = r_xcpt_uop_fu_code; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_br_type = r_xcpt_uop_ctrl_br_type; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_op1_sel = r_xcpt_uop_ctrl_op1_sel; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_op2_sel = r_xcpt_uop_ctrl_op2_sel; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_imm_sel = r_xcpt_uop_ctrl_imm_sel; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_op_fcn = r_xcpt_uop_ctrl_op_fcn; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_fcn_dw = r_xcpt_uop_ctrl_fcn_dw; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_rf_wen = r_xcpt_uop_ctrl_rf_wen; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_csr_cmd = r_xcpt_uop_ctrl_csr_cmd; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_is_load = r_xcpt_uop_ctrl_is_load; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_is_sta = r_xcpt_uop_ctrl_is_sta; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ctrl_is_std = r_xcpt_uop_ctrl_is_std; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_wakeup_delay = r_xcpt_uop_wakeup_delay; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_allocate_brtag = r_xcpt_uop_allocate_brtag; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_br_or_jmp = r_xcpt_uop_is_br_or_jmp; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_jump = r_xcpt_uop_is_jump; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_jal = r_xcpt_uop_is_jal; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_ret = r_xcpt_uop_is_ret; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_call = r_xcpt_uop_is_call; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_mask = r_xcpt_uop_br_mask; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_tag = r_xcpt_uop_br_tag; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_prediction_bpd_predict_val = r_xcpt_uop_br_prediction_bpd_predict_val; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_prediction_bpd_predict_taken = r_xcpt_uop_br_prediction_bpd_predict_taken; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_prediction_btb_hit = r_xcpt_uop_br_prediction_btb_hit; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_prediction_btb_predicted = r_xcpt_uop_br_prediction_btb_predicted; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_br_prediction_is_br_or_jalr = r_xcpt_uop_br_prediction_is_br_or_jalr; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stat_brjmp_mispredicted = r_xcpt_uop_stat_brjmp_mispredicted; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stat_btb_made_pred = r_xcpt_uop_stat_btb_made_pred; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stat_btb_mispredicted = r_xcpt_uop_stat_btb_mispredicted; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stat_bpd_made_pred = r_xcpt_uop_stat_bpd_made_pred; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stat_bpd_mispredicted = r_xcpt_uop_stat_bpd_mispredicted; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_fetch_pc_lob = r_xcpt_uop_fetch_pc_lob; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_imm_packed = r_xcpt_uop_imm_packed; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_csr_addr = r_xcpt_uop_csr_addr; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_rob_idx = r_xcpt_uop_rob_idx; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ldq_idx = r_xcpt_uop_ldq_idx; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stq_idx = r_xcpt_uop_stq_idx; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_brob_idx = r_xcpt_uop_brob_idx; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_pdst = r_xcpt_uop_pdst; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_pop1 = r_xcpt_uop_pop1; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_pop2 = r_xcpt_uop_pop2; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_pop3 = r_xcpt_uop_pop3; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_prs1_busy = r_xcpt_uop_prs1_busy; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_prs2_busy = r_xcpt_uop_prs2_busy; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_prs3_busy = r_xcpt_uop_prs3_busy; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_stale_pdst = r_xcpt_uop_stale_pdst; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_exception = r_xcpt_uop_exception; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_exc_cause = r_xcpt_uop_exc_cause; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_bypassable = r_xcpt_uop_bypassable; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_mem_cmd = r_xcpt_uop_mem_cmd; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_mem_typ = r_xcpt_uop_mem_typ; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_fence = r_xcpt_uop_is_fence; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_fencei = r_xcpt_uop_is_fencei; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_store = r_xcpt_uop_is_store; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_amo = r_xcpt_uop_is_amo; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_load = r_xcpt_uop_is_load; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_is_unique = r_xcpt_uop_is_unique; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_flush_on_commit = r_xcpt_uop_flush_on_commit; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ldst = r_xcpt_uop_ldst; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_lrs1 = r_xcpt_uop_lrs1; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_lrs2 = r_xcpt_uop_lrs2; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_lrs3 = r_xcpt_uop_lrs3; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_ldst_val = r_xcpt_uop_ldst_val; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_dst_rtype = r_xcpt_uop_dst_rtype; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_lrs1_rtype = r_xcpt_uop_lrs1_rtype; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_lrs2_rtype = r_xcpt_uop_lrs2_rtype; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_frs3_en = r_xcpt_uop_frs3_en; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_fp_val = r_xcpt_uop_fp_val; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_fp_single = r_xcpt_uop_fp_single; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_xcpt_if = r_xcpt_uop_xcpt_if; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_replay_if = r_xcpt_uop_replay_if; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_debug_wdata = r_xcpt_uop_debug_wdata; // @[rob.scala 881:22]
  assign io_debug_xcpt_uop_debug_events_fetch_seq = r_xcpt_uop_debug_events_fetch_seq; // @[rob.scala 881:22]
  assign io_debug_xcpt_badvaddr = new_DoPrim4430178; // @[rob.scala 882:27]
  always @(posedge clk) begin
    if(T_23555_T_23571_en & T_23555_T_23571_mask) begin
      T_23555[T_23555_T_23571_addr] <= T_23555_T_23571_data; // @[rob.scala 893:22]
    end
    if(T_23558_T_23566_en & T_23558_T_23566_mask) begin
      T_23558[T_23558_T_23566_addr] <= T_23558_T_23566_data; // @[rob.scala 894:22]
    end
    if(row_metadata_brob_idx_T_23653_en & row_metadata_brob_idx_T_23653_mask) begin
      row_metadata_brob_idx[row_metadata_brob_idx_T_23653_addr] <= row_metadata_brob_idx_T_23653_data; // @[rob.scala 295:35]
    end
    if(row_metadata_has_brorjalr_T_23654_en & row_metadata_has_brorjalr_T_23654_mask) begin
      row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_23654_addr] <= row_metadata_has_brorjalr_T_23654_data; // @[rob.scala 296:38]
    end
    if(row_metadata_has_brorjalr_T_23662_en & row_metadata_has_brorjalr_T_23662_mask) begin
      row_metadata_has_brorjalr[row_metadata_has_brorjalr_T_23662_addr] <= row_metadata_has_brorjalr_T_23662_data; // @[rob.scala 296:38]
    end
    if(T_23710_T_28316_en & T_23710_T_28316_mask) begin
      T_23710[T_23710_T_28316_addr] <= T_23710_T_28316_data; // @[rob.scala 335:30]
    end
    if(T_23710_T_28594_en & T_23710_T_28594_mask) begin
      T_23710[T_23710_T_28594_addr] <= T_23710_T_28594_data; // @[rob.scala 335:30]
    end
    if(T_23710_T_28602_en & T_23710_T_28602_mask) begin
      T_23710[T_23710_T_28602_addr] <= T_23710_T_28602_data; // @[rob.scala 335:30]
    end
    if(T_23710_T_28610_en & T_23710_T_28610_mask) begin
      T_23710[T_23710_T_28610_addr] <= T_23710_T_28610_data; // @[rob.scala 335:30]
    end
    if(T_23710_T_28618_en & T_23710_T_28618_mask) begin
      T_23710[T_23710_T_28618_addr] <= T_23710_T_28618_data; // @[rob.scala 335:30]
    end
    if(T_28311_T_28407_en & T_28311_T_28407_mask) begin
      T_28311[T_28311_T_28407_addr] <= T_28311_T_28407_data; // @[rob.scala 339:30]
    end
    if(T_28311_T_29079_en & T_28311_T_29079_mask) begin
      T_28311[T_28311_T_29079_addr] <= T_28311_T_29079_data; // @[rob.scala 339:30]
    end
    if(T_28311_T_29087_en & T_28311_T_29087_mask) begin
      T_28311[T_28311_T_29087_addr] <= T_28311_T_29087_data; // @[rob.scala 339:30]
    end
    if(T_28311_T_29363_en & T_28311_T_29363_mask) begin
      T_28311[T_28311_T_29363_addr] <= T_28311_T_29363_data; // @[rob.scala 339:30]
    end
    if(T_28314_T_28408_en & T_28314_T_28408_mask) begin
      T_28314[T_28314_T_28408_addr] <= T_28314_T_28408_data; // @[rob.scala 340:30]
    end
    if(T_28314_T_29065_en & T_28314_T_29065_mask) begin
      T_28314[T_28314_T_29065_addr] <= T_28314_T_29065_data; // @[rob.scala 340:30]
    end
    if(T_28314_T_29072_en & T_28314_T_29072_mask) begin
      T_28314[T_28314_T_29072_addr] <= T_28314_T_29072_data; // @[rob.scala 340:30]
    end
    if(T_35638_T_40244_en & T_35638_T_40244_mask) begin
      T_35638[T_35638_T_40244_addr] <= T_35638_T_40244_data; // @[rob.scala 335:30]
    end
    if(T_35638_T_40522_en & T_35638_T_40522_mask) begin
      T_35638[T_35638_T_40522_addr] <= T_35638_T_40522_data; // @[rob.scala 335:30]
    end
    if(T_35638_T_40530_en & T_35638_T_40530_mask) begin
      T_35638[T_35638_T_40530_addr] <= T_35638_T_40530_data; // @[rob.scala 335:30]
    end
    if(T_35638_T_40538_en & T_35638_T_40538_mask) begin
      T_35638[T_35638_T_40538_addr] <= T_35638_T_40538_data; // @[rob.scala 335:30]
    end
    if(T_35638_T_40546_en & T_35638_T_40546_mask) begin
      T_35638[T_35638_T_40546_addr] <= T_35638_T_40546_data; // @[rob.scala 335:30]
    end
    if(T_40239_T_40335_en & T_40239_T_40335_mask) begin
      T_40239[T_40239_T_40335_addr] <= T_40239_T_40335_data; // @[rob.scala 339:30]
    end
    if(T_40239_T_41007_en & T_40239_T_41007_mask) begin
      T_40239[T_40239_T_41007_addr] <= T_40239_T_41007_data; // @[rob.scala 339:30]
    end
    if(T_40239_T_41015_en & T_40239_T_41015_mask) begin
      T_40239[T_40239_T_41015_addr] <= T_40239_T_41015_data; // @[rob.scala 339:30]
    end
    if(T_40239_T_41291_en & T_40239_T_41291_mask) begin
      T_40239[T_40239_T_41291_addr] <= T_40239_T_41291_data; // @[rob.scala 339:30]
    end
    if(T_40242_T_40336_en & T_40242_T_40336_mask) begin
      T_40242[T_40242_T_40336_addr] <= T_40242_T_40336_data; // @[rob.scala 340:30]
    end
    if(T_40242_T_40993_en & T_40242_T_40993_mask) begin
      T_40242[T_40242_T_40993_addr] <= T_40242_T_40993_data; // @[rob.scala 340:30]
    end
    if(T_40242_T_41000_en & T_40242_T_41000_mask) begin
      T_40242[T_40242_T_41000_addr] <= T_40242_T_41000_data; // @[rob.scala 340:30]
    end
    if (reset) begin
      rob_state <= 2'h0;
    end else if (T_48207) begin // @[Conditional.scala 24:73]
      if (T_48210) begin // @[rob.scala 810:13]
        rob_state <= 2'h1; // @[rob.scala 811:26]
      end else if (T_47568) begin // @[rob.scala 806:13]
        rob_state <= 2'h2; // @[rob.scala 807:26]
      end else begin
        rob_state <= _GEN_28807;
      end
    end else begin
      rob_state <= _GEN_28807;
    end
    if (reset) begin
      rob_head <= 5'h0;
    end else if (T_48134) begin // @[rob.scala 719:4]
      if (T_48136) begin // @[util.scala 76:13]
        rob_head <= 5'h0;
      end else begin
        rob_head <= T_48140;
      end
    end
    if (reset) begin
      rob_tail <= 5'h0;
    end else begin
      rob_tail <= _GEN_28799[4:0];
    end
    if (reset) begin
      r_xcpt_val <= 1'h0;
    end else if (T_48093) begin // @[rob.scala 689:4]
      r_xcpt_val <= 1'h0; // @[rob.scala 690:18]
    end else if (T_47875) begin // @[rob.scala 660:4]
      r_xcpt_val <= _GEN_28635;
    end
    r_xcpt_uop_valid <= next_xcpt_uop_valid; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_iw_state <= next_xcpt_uop_iw_state; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_uopc <= next_xcpt_uop_uopc; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_inst <= next_xcpt_uop_inst; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_pc <= next_xcpt_uop_pc; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_fu_code <= next_xcpt_uop_fu_code; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_br_type <= next_xcpt_uop_ctrl_br_type; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_op1_sel <= next_xcpt_uop_ctrl_op1_sel; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_op2_sel <= next_xcpt_uop_ctrl_op2_sel; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_imm_sel <= next_xcpt_uop_ctrl_imm_sel; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_op_fcn <= next_xcpt_uop_ctrl_op_fcn; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_fcn_dw <= next_xcpt_uop_ctrl_fcn_dw; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_rf_wen <= next_xcpt_uop_ctrl_rf_wen; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_csr_cmd <= next_xcpt_uop_ctrl_csr_cmd; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_is_load <= next_xcpt_uop_ctrl_is_load; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_is_sta <= next_xcpt_uop_ctrl_is_sta; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ctrl_is_std <= next_xcpt_uop_ctrl_is_std; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_wakeup_delay <= next_xcpt_uop_wakeup_delay; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_allocate_brtag <= next_xcpt_uop_allocate_brtag; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_br_or_jmp <= next_xcpt_uop_is_br_or_jmp; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_jump <= next_xcpt_uop_is_jump; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_jal <= next_xcpt_uop_is_jal; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_ret <= next_xcpt_uop_is_ret; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_call <= next_xcpt_uop_is_call; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_br_mask <= T_48087; // @[util.scala 32:17]
    r_xcpt_uop_br_tag <= next_xcpt_uop_br_tag; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_br_prediction_bpd_predict_val <= next_xcpt_uop_br_prediction_bpd_predict_val; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_br_prediction_bpd_predict_taken <= next_xcpt_uop_br_prediction_bpd_predict_taken; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_br_prediction_btb_hit <= next_xcpt_uop_br_prediction_btb_hit; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_br_prediction_btb_predicted <= next_xcpt_uop_br_prediction_btb_predicted; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_br_prediction_is_br_or_jalr <= next_xcpt_uop_br_prediction_is_br_or_jalr; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stat_brjmp_mispredicted <= next_xcpt_uop_stat_brjmp_mispredicted; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stat_btb_made_pred <= next_xcpt_uop_stat_btb_made_pred; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stat_btb_mispredicted <= next_xcpt_uop_stat_btb_mispredicted; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stat_bpd_made_pred <= next_xcpt_uop_stat_bpd_made_pred; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stat_bpd_mispredicted <= next_xcpt_uop_stat_bpd_mispredicted; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_fetch_pc_lob <= next_xcpt_uop_fetch_pc_lob; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_imm_packed <= next_xcpt_uop_imm_packed; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_csr_addr <= next_xcpt_uop_csr_addr; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_rob_idx <= next_xcpt_uop_rob_idx; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ldq_idx <= next_xcpt_uop_ldq_idx; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stq_idx <= next_xcpt_uop_stq_idx; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_brob_idx <= next_xcpt_uop_brob_idx; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_pdst <= next_xcpt_uop_pdst; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_pop1 <= next_xcpt_uop_pop1; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_pop2 <= next_xcpt_uop_pop2; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_pop3 <= next_xcpt_uop_pop3; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_prs1_busy <= next_xcpt_uop_prs1_busy; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_prs2_busy <= next_xcpt_uop_prs2_busy; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_prs3_busy <= next_xcpt_uop_prs3_busy; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_stale_pdst <= next_xcpt_uop_stale_pdst; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_exception <= next_xcpt_uop_exception; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_exc_cause <= next_xcpt_uop_exc_cause; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_bypassable <= next_xcpt_uop_bypassable; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_mem_cmd <= next_xcpt_uop_mem_cmd; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_mem_typ <= next_xcpt_uop_mem_typ; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_fence <= next_xcpt_uop_is_fence; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_fencei <= next_xcpt_uop_is_fencei; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_store <= next_xcpt_uop_is_store; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_amo <= next_xcpt_uop_is_amo; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_load <= next_xcpt_uop_is_load; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_is_unique <= next_xcpt_uop_is_unique; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_flush_on_commit <= next_xcpt_uop_flush_on_commit; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ldst <= next_xcpt_uop_ldst; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_lrs1 <= next_xcpt_uop_lrs1; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_lrs2 <= next_xcpt_uop_lrs2; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_lrs3 <= next_xcpt_uop_lrs3; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_ldst_val <= next_xcpt_uop_ldst_val; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_dst_rtype <= next_xcpt_uop_dst_rtype; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_lrs1_rtype <= next_xcpt_uop_lrs1_rtype; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_lrs2_rtype <= next_xcpt_uop_lrs2_rtype; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_frs3_en <= next_xcpt_uop_frs3_en; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_fp_val <= next_xcpt_uop_fp_val; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_fp_single <= next_xcpt_uop_fp_single; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_xcpt_if <= next_xcpt_uop_xcpt_if; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_replay_if <= next_xcpt_uop_replay_if; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_debug_wdata <= next_xcpt_uop_debug_wdata; // @[rob.scala 660:4 rob.scala 652:18]
    r_xcpt_uop_debug_events_fetch_seq <= next_xcpt_uop_debug_events_fetch_seq; // @[rob.scala 660:4 rob.scala 652:18]
    if (T_47875) begin // @[rob.scala 660:4]
      if (T_47991) begin // @[rob.scala 676:7]
        r_xcpt_badvaddr <= T_48084; // @[rob.scala 682:26]
      end else if (T_47876) begin // @[rob.scala 662:7]
        if (T_47981) begin // @[rob.scala 668:10]
          r_xcpt_badvaddr <= T_47984; // @[rob.scala 672:37]
        end
      end
    end
    if (reset) begin
      T_35634_23 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h17 == rob_head) begin // @[rob.scala 500:28]
        T_35634_23 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_23 <= _GEN_20392;
      end
    end else begin
      T_35634_23 <= _GEN_20392;
    end
    if (reset) begin
      T_35634_22 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h16 == rob_head) begin // @[rob.scala 500:28]
        T_35634_22 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_22 <= _GEN_20389;
      end
    end else begin
      T_35634_22 <= _GEN_20389;
    end
    if (reset) begin
      T_35634_21 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h15 == rob_head) begin // @[rob.scala 500:28]
        T_35634_21 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_21 <= _GEN_20386;
      end
    end else begin
      T_35634_21 <= _GEN_20386;
    end
    if (reset) begin
      T_35634_20 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h14 == rob_head) begin // @[rob.scala 500:28]
        T_35634_20 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_20 <= _GEN_20383;
      end
    end else begin
      T_35634_20 <= _GEN_20383;
    end
    if (reset) begin
      T_35634_19 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h13 == rob_head) begin // @[rob.scala 500:28]
        T_35634_19 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_19 <= _GEN_20380;
      end
    end else begin
      T_35634_19 <= _GEN_20380;
    end
    if (reset) begin
      T_35634_18 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h12 == rob_head) begin // @[rob.scala 500:28]
        T_35634_18 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_18 <= _GEN_20377;
      end
    end else begin
      T_35634_18 <= _GEN_20377;
    end
    if (reset) begin
      T_35634_17 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h11 == rob_head) begin // @[rob.scala 500:28]
        T_35634_17 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_17 <= _GEN_20374;
      end
    end else begin
      T_35634_17 <= _GEN_20374;
    end
    if (reset) begin
      T_35634_16 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h10 == rob_head) begin // @[rob.scala 500:28]
        T_35634_16 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_16 <= _GEN_20371;
      end
    end else begin
      T_35634_16 <= _GEN_20371;
    end
    if (reset) begin
      T_35634_15 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'hf == rob_head) begin // @[rob.scala 500:28]
        T_35634_15 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_15 <= _GEN_20368;
      end
    end else begin
      T_35634_15 <= _GEN_20368;
    end
    if (reset) begin
      T_35634_14 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'he == rob_head) begin // @[rob.scala 500:28]
        T_35634_14 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_14 <= _GEN_20365;
      end
    end else begin
      T_35634_14 <= _GEN_20365;
    end
    if (reset) begin
      T_35634_13 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'hd == rob_head) begin // @[rob.scala 500:28]
        T_35634_13 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_13 <= _GEN_20362;
      end
    end else begin
      T_35634_13 <= _GEN_20362;
    end
    if (reset) begin
      T_35634_12 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'hc == rob_head) begin // @[rob.scala 500:28]
        T_35634_12 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_12 <= _GEN_20359;
      end
    end else begin
      T_35634_12 <= _GEN_20359;
    end
    if (reset) begin
      T_35634_11 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'hb == rob_head) begin // @[rob.scala 500:28]
        T_35634_11 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_11 <= _GEN_20356;
      end
    end else begin
      T_35634_11 <= _GEN_20356;
    end
    if (reset) begin
      T_35634_10 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'ha == rob_head) begin // @[rob.scala 500:28]
        T_35634_10 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_10 <= _GEN_20353;
      end
    end else begin
      T_35634_10 <= _GEN_20353;
    end
    if (reset) begin
      T_35634_9 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h9 == rob_head) begin // @[rob.scala 500:28]
        T_35634_9 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_9 <= _GEN_20350;
      end
    end else begin
      T_35634_9 <= _GEN_20350;
    end
    if (reset) begin
      T_35634_8 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h8 == rob_head) begin // @[rob.scala 500:28]
        T_35634_8 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_8 <= _GEN_20347;
      end
    end else begin
      T_35634_8 <= _GEN_20347;
    end
    if (reset) begin
      T_35634_7 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h7 == rob_head) begin // @[rob.scala 500:28]
        T_35634_7 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_7 <= _GEN_20344;
      end
    end else begin
      T_35634_7 <= _GEN_20344;
    end
    if (reset) begin
      T_35634_6 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h6 == rob_head) begin // @[rob.scala 500:28]
        T_35634_6 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_6 <= _GEN_20341;
      end
    end else begin
      T_35634_6 <= _GEN_20341;
    end
    if (reset) begin
      T_35634_5 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h5 == rob_head) begin // @[rob.scala 500:28]
        T_35634_5 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_5 <= _GEN_20338;
      end
    end else begin
      T_35634_5 <= _GEN_20338;
    end
    if (reset) begin
      T_35634_4 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h4 == rob_head) begin // @[rob.scala 500:28]
        T_35634_4 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_4 <= _GEN_20335;
      end
    end else begin
      T_35634_4 <= _GEN_20335;
    end
    if (reset) begin
      T_35634_3 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h3 == rob_head) begin // @[rob.scala 500:28]
        T_35634_3 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_3 <= _GEN_20332;
      end
    end else begin
      T_35634_3 <= _GEN_20332;
    end
    if (reset) begin
      T_35634_2 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h2 == rob_head) begin // @[rob.scala 500:28]
        T_35634_2 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_2 <= _GEN_20329;
      end
    end else begin
      T_35634_2 <= _GEN_20329;
    end
    if (reset) begin
      T_35634_1 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h1 == rob_head) begin // @[rob.scala 500:28]
        T_35634_1 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_1 <= _GEN_20326;
      end
    end else begin
      T_35634_1 <= _GEN_20326;
    end
    if (reset) begin
      T_35634_0 <= 1'h0;
    end else if (T_47563) begin // @[rob.scala 499:7]
      if (5'h0 == rob_head) begin // @[rob.scala 500:28]
        T_35634_0 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_35634_0 <= _GEN_20323;
      end
    end else begin
      T_35634_0 <= _GEN_20323;
    end
    if (reset) begin
      T_23706_23 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h17 == rob_head) begin // @[rob.scala 500:28]
        T_23706_23 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_23 <= _GEN_6249;
      end
    end else begin
      T_23706_23 <= _GEN_6249;
    end
    if (reset) begin
      T_23706_22 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h16 == rob_head) begin // @[rob.scala 500:28]
        T_23706_22 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_22 <= _GEN_6246;
      end
    end else begin
      T_23706_22 <= _GEN_6246;
    end
    if (reset) begin
      T_23706_21 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h15 == rob_head) begin // @[rob.scala 500:28]
        T_23706_21 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_21 <= _GEN_6243;
      end
    end else begin
      T_23706_21 <= _GEN_6243;
    end
    if (reset) begin
      T_23706_20 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h14 == rob_head) begin // @[rob.scala 500:28]
        T_23706_20 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_20 <= _GEN_6240;
      end
    end else begin
      T_23706_20 <= _GEN_6240;
    end
    if (reset) begin
      T_23706_19 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h13 == rob_head) begin // @[rob.scala 500:28]
        T_23706_19 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_19 <= _GEN_6237;
      end
    end else begin
      T_23706_19 <= _GEN_6237;
    end
    if (reset) begin
      T_23706_18 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h12 == rob_head) begin // @[rob.scala 500:28]
        T_23706_18 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_18 <= _GEN_6234;
      end
    end else begin
      T_23706_18 <= _GEN_6234;
    end
    if (reset) begin
      T_23706_17 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h11 == rob_head) begin // @[rob.scala 500:28]
        T_23706_17 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_17 <= _GEN_6231;
      end
    end else begin
      T_23706_17 <= _GEN_6231;
    end
    if (reset) begin
      T_23706_16 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h10 == rob_head) begin // @[rob.scala 500:28]
        T_23706_16 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_16 <= _GEN_6228;
      end
    end else begin
      T_23706_16 <= _GEN_6228;
    end
    if (reset) begin
      T_23706_15 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'hf == rob_head) begin // @[rob.scala 500:28]
        T_23706_15 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_15 <= _GEN_6225;
      end
    end else begin
      T_23706_15 <= _GEN_6225;
    end
    if (reset) begin
      T_23706_14 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'he == rob_head) begin // @[rob.scala 500:28]
        T_23706_14 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_14 <= _GEN_6222;
      end
    end else begin
      T_23706_14 <= _GEN_6222;
    end
    if (reset) begin
      T_23706_13 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'hd == rob_head) begin // @[rob.scala 500:28]
        T_23706_13 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_13 <= _GEN_6219;
      end
    end else begin
      T_23706_13 <= _GEN_6219;
    end
    if (reset) begin
      T_23706_12 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'hc == rob_head) begin // @[rob.scala 500:28]
        T_23706_12 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_12 <= _GEN_6216;
      end
    end else begin
      T_23706_12 <= _GEN_6216;
    end
    if (reset) begin
      T_23706_11 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'hb == rob_head) begin // @[rob.scala 500:28]
        T_23706_11 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_11 <= _GEN_6213;
      end
    end else begin
      T_23706_11 <= _GEN_6213;
    end
    if (reset) begin
      T_23706_10 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'ha == rob_head) begin // @[rob.scala 500:28]
        T_23706_10 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_10 <= _GEN_6210;
      end
    end else begin
      T_23706_10 <= _GEN_6210;
    end
    if (reset) begin
      T_23706_9 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h9 == rob_head) begin // @[rob.scala 500:28]
        T_23706_9 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_9 <= _GEN_6207;
      end
    end else begin
      T_23706_9 <= _GEN_6207;
    end
    if (reset) begin
      T_23706_8 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h8 == rob_head) begin // @[rob.scala 500:28]
        T_23706_8 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_8 <= _GEN_6204;
      end
    end else begin
      T_23706_8 <= _GEN_6204;
    end
    if (reset) begin
      T_23706_7 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h7 == rob_head) begin // @[rob.scala 500:28]
        T_23706_7 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_7 <= _GEN_6201;
      end
    end else begin
      T_23706_7 <= _GEN_6201;
    end
    if (reset) begin
      T_23706_6 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h6 == rob_head) begin // @[rob.scala 500:28]
        T_23706_6 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_6 <= _GEN_6198;
      end
    end else begin
      T_23706_6 <= _GEN_6198;
    end
    if (reset) begin
      T_23706_5 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h5 == rob_head) begin // @[rob.scala 500:28]
        T_23706_5 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_5 <= _GEN_6195;
      end
    end else begin
      T_23706_5 <= _GEN_6195;
    end
    if (reset) begin
      T_23706_4 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h4 == rob_head) begin // @[rob.scala 500:28]
        T_23706_4 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_4 <= _GEN_6192;
      end
    end else begin
      T_23706_4 <= _GEN_6192;
    end
    if (reset) begin
      T_23706_3 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h3 == rob_head) begin // @[rob.scala 500:28]
        T_23706_3 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_3 <= _GEN_6189;
      end
    end else begin
      T_23706_3 <= _GEN_6189;
    end
    if (reset) begin
      T_23706_2 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h2 == rob_head) begin // @[rob.scala 500:28]
        T_23706_2 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_2 <= _GEN_6186;
      end
    end else begin
      T_23706_2 <= _GEN_6186;
    end
    if (reset) begin
      T_23706_1 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h1 == rob_head) begin // @[rob.scala 500:28]
        T_23706_1 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_1 <= _GEN_6183;
      end
    end else begin
      T_23706_1 <= _GEN_6183;
    end
    if (reset) begin
      T_23706_0 <= 1'h0;
    end else if (T_47546) begin // @[rob.scala 499:7]
      if (5'h0 == rob_head) begin // @[rob.scala 500:28]
        T_23706_0 <= 1'h0; // @[rob.scala 500:28]
      end else begin
        T_23706_0 <= _GEN_6180;
      end
    end else begin
      T_23706_0 <= _GEN_6180;
    end
    if (reset) begin
      r_partial_row <= 1'h0;
    end else if (T_23661) begin // @[rob.scala 304:4]
      r_partial_row <= io_dis_partial_stall; // @[rob.scala 305:21]
    end else if (T_23652) begin // @[rob.scala 298:4]
      r_partial_row <= io_dis_partial_stall; // @[rob.scala 301:21]
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_0_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_0_inst <= _GEN_8220;
      end
    end else begin
      T_26182_0_inst <= _GEN_8220;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_29464) begin // @[rob.scala 490:10]
      T_26182_0_br_mask <= T_29466; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 402:72]
        T_26182_0_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_0_stat_brjmp_mispredicted <= _GEN_2726;
      end
    end else begin
      T_26182_0_stat_brjmp_mispredicted <= _GEN_2726;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 404:72]
        T_26182_0_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_0_stat_btb_made_pred <= _GEN_2750;
      end
    end else begin
      T_26182_0_stat_btb_made_pred <= _GEN_2750;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 403:72]
        T_26182_0_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_0_stat_btb_mispredicted <= _GEN_2774;
      end
    end else begin
      T_26182_0_stat_btb_mispredicted <= _GEN_2774;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 406:72]
        T_26182_0_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_0_stat_bpd_made_pred <= _GEN_2798;
      end
    end else begin
      T_26182_0_stat_bpd_made_pred <= _GEN_2798;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 405:72]
        T_26182_0_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_0_stat_bpd_mispredicted <= _GEN_2822;
      end
    end else begin
      T_26182_0_stat_bpd_mispredicted <= _GEN_2822;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h0 == T_28605) begin // @[rob.scala 531:53]
        T_26182_0_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_0_debug_wdata <= _GEN_10260;
      end
    end else begin
      T_26182_0_debug_wdata <= _GEN_10260;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_0_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_1_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_1_inst <= _GEN_8221;
      end
    end else begin
      T_26182_1_inst <= _GEN_8221;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_29566) begin // @[rob.scala 490:10]
      T_26182_1_br_mask <= T_29568; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 402:72]
        T_26182_1_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_1_stat_brjmp_mispredicted <= _GEN_2727;
      end
    end else begin
      T_26182_1_stat_brjmp_mispredicted <= _GEN_2727;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 404:72]
        T_26182_1_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_1_stat_btb_made_pred <= _GEN_2751;
      end
    end else begin
      T_26182_1_stat_btb_made_pred <= _GEN_2751;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 403:72]
        T_26182_1_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_1_stat_btb_mispredicted <= _GEN_2775;
      end
    end else begin
      T_26182_1_stat_btb_mispredicted <= _GEN_2775;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 406:72]
        T_26182_1_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_1_stat_bpd_made_pred <= _GEN_2799;
      end
    end else begin
      T_26182_1_stat_bpd_made_pred <= _GEN_2799;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 405:72]
        T_26182_1_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_1_stat_bpd_mispredicted <= _GEN_2823;
      end
    end else begin
      T_26182_1_stat_bpd_mispredicted <= _GEN_2823;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h1 == T_28605) begin // @[rob.scala 531:53]
        T_26182_1_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_1_debug_wdata <= _GEN_10261;
      end
    end else begin
      T_26182_1_debug_wdata <= _GEN_10261;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_1_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_2_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_2_inst <= _GEN_8222;
      end
    end else begin
      T_26182_2_inst <= _GEN_8222;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_29668) begin // @[rob.scala 490:10]
      T_26182_2_br_mask <= T_29670; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 402:72]
        T_26182_2_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_2_stat_brjmp_mispredicted <= _GEN_2728;
      end
    end else begin
      T_26182_2_stat_brjmp_mispredicted <= _GEN_2728;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 404:72]
        T_26182_2_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_2_stat_btb_made_pred <= _GEN_2752;
      end
    end else begin
      T_26182_2_stat_btb_made_pred <= _GEN_2752;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 403:72]
        T_26182_2_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_2_stat_btb_mispredicted <= _GEN_2776;
      end
    end else begin
      T_26182_2_stat_btb_mispredicted <= _GEN_2776;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 406:72]
        T_26182_2_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_2_stat_bpd_made_pred <= _GEN_2800;
      end
    end else begin
      T_26182_2_stat_bpd_made_pred <= _GEN_2800;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 405:72]
        T_26182_2_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_2_stat_bpd_mispredicted <= _GEN_2824;
      end
    end else begin
      T_26182_2_stat_bpd_mispredicted <= _GEN_2824;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h2 == T_28605) begin // @[rob.scala 531:53]
        T_26182_2_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_2_debug_wdata <= _GEN_10262;
      end
    end else begin
      T_26182_2_debug_wdata <= _GEN_10262;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_2_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_3_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_3_inst <= _GEN_8223;
      end
    end else begin
      T_26182_3_inst <= _GEN_8223;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_29770) begin // @[rob.scala 490:10]
      T_26182_3_br_mask <= T_29772; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 402:72]
        T_26182_3_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_3_stat_brjmp_mispredicted <= _GEN_2729;
      end
    end else begin
      T_26182_3_stat_brjmp_mispredicted <= _GEN_2729;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 404:72]
        T_26182_3_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_3_stat_btb_made_pred <= _GEN_2753;
      end
    end else begin
      T_26182_3_stat_btb_made_pred <= _GEN_2753;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 403:72]
        T_26182_3_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_3_stat_btb_mispredicted <= _GEN_2777;
      end
    end else begin
      T_26182_3_stat_btb_mispredicted <= _GEN_2777;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 406:72]
        T_26182_3_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_3_stat_bpd_made_pred <= _GEN_2801;
      end
    end else begin
      T_26182_3_stat_bpd_made_pred <= _GEN_2801;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 405:72]
        T_26182_3_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_3_stat_bpd_mispredicted <= _GEN_2825;
      end
    end else begin
      T_26182_3_stat_bpd_mispredicted <= _GEN_2825;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h3 == T_28605) begin // @[rob.scala 531:53]
        T_26182_3_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_3_debug_wdata <= _GEN_10263;
      end
    end else begin
      T_26182_3_debug_wdata <= _GEN_10263;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_3_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_4_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_4_inst <= _GEN_8224;
      end
    end else begin
      T_26182_4_inst <= _GEN_8224;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_29872) begin // @[rob.scala 490:10]
      T_26182_4_br_mask <= T_29874; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 402:72]
        T_26182_4_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_4_stat_brjmp_mispredicted <= _GEN_2730;
      end
    end else begin
      T_26182_4_stat_brjmp_mispredicted <= _GEN_2730;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 404:72]
        T_26182_4_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_4_stat_btb_made_pred <= _GEN_2754;
      end
    end else begin
      T_26182_4_stat_btb_made_pred <= _GEN_2754;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 403:72]
        T_26182_4_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_4_stat_btb_mispredicted <= _GEN_2778;
      end
    end else begin
      T_26182_4_stat_btb_mispredicted <= _GEN_2778;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 406:72]
        T_26182_4_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_4_stat_bpd_made_pred <= _GEN_2802;
      end
    end else begin
      T_26182_4_stat_bpd_made_pred <= _GEN_2802;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 405:72]
        T_26182_4_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_4_stat_bpd_mispredicted <= _GEN_2826;
      end
    end else begin
      T_26182_4_stat_bpd_mispredicted <= _GEN_2826;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h4 == T_28605) begin // @[rob.scala 531:53]
        T_26182_4_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_4_debug_wdata <= _GEN_10264;
      end
    end else begin
      T_26182_4_debug_wdata <= _GEN_10264;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_4_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_5_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_5_inst <= _GEN_8225;
      end
    end else begin
      T_26182_5_inst <= _GEN_8225;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_29974) begin // @[rob.scala 490:10]
      T_26182_5_br_mask <= T_29976; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 402:72]
        T_26182_5_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_5_stat_brjmp_mispredicted <= _GEN_2731;
      end
    end else begin
      T_26182_5_stat_brjmp_mispredicted <= _GEN_2731;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 404:72]
        T_26182_5_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_5_stat_btb_made_pred <= _GEN_2755;
      end
    end else begin
      T_26182_5_stat_btb_made_pred <= _GEN_2755;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 403:72]
        T_26182_5_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_5_stat_btb_mispredicted <= _GEN_2779;
      end
    end else begin
      T_26182_5_stat_btb_mispredicted <= _GEN_2779;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 406:72]
        T_26182_5_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_5_stat_bpd_made_pred <= _GEN_2803;
      end
    end else begin
      T_26182_5_stat_bpd_made_pred <= _GEN_2803;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 405:72]
        T_26182_5_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_5_stat_bpd_mispredicted <= _GEN_2827;
      end
    end else begin
      T_26182_5_stat_bpd_mispredicted <= _GEN_2827;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h5 == T_28605) begin // @[rob.scala 531:53]
        T_26182_5_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_5_debug_wdata <= _GEN_10265;
      end
    end else begin
      T_26182_5_debug_wdata <= _GEN_10265;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_5_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_6_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_6_inst <= _GEN_8226;
      end
    end else begin
      T_26182_6_inst <= _GEN_8226;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30076) begin // @[rob.scala 490:10]
      T_26182_6_br_mask <= T_30078; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 402:72]
        T_26182_6_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_6_stat_brjmp_mispredicted <= _GEN_2732;
      end
    end else begin
      T_26182_6_stat_brjmp_mispredicted <= _GEN_2732;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 404:72]
        T_26182_6_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_6_stat_btb_made_pred <= _GEN_2756;
      end
    end else begin
      T_26182_6_stat_btb_made_pred <= _GEN_2756;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 403:72]
        T_26182_6_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_6_stat_btb_mispredicted <= _GEN_2780;
      end
    end else begin
      T_26182_6_stat_btb_mispredicted <= _GEN_2780;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 406:72]
        T_26182_6_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_6_stat_bpd_made_pred <= _GEN_2804;
      end
    end else begin
      T_26182_6_stat_bpd_made_pred <= _GEN_2804;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 405:72]
        T_26182_6_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_6_stat_bpd_mispredicted <= _GEN_2828;
      end
    end else begin
      T_26182_6_stat_bpd_mispredicted <= _GEN_2828;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h6 == T_28605) begin // @[rob.scala 531:53]
        T_26182_6_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_6_debug_wdata <= _GEN_10266;
      end
    end else begin
      T_26182_6_debug_wdata <= _GEN_10266;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_6_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_7_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_7_inst <= _GEN_8227;
      end
    end else begin
      T_26182_7_inst <= _GEN_8227;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30178) begin // @[rob.scala 490:10]
      T_26182_7_br_mask <= T_30180; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 402:72]
        T_26182_7_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_7_stat_brjmp_mispredicted <= _GEN_2733;
      end
    end else begin
      T_26182_7_stat_brjmp_mispredicted <= _GEN_2733;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 404:72]
        T_26182_7_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_7_stat_btb_made_pred <= _GEN_2757;
      end
    end else begin
      T_26182_7_stat_btb_made_pred <= _GEN_2757;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 403:72]
        T_26182_7_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_7_stat_btb_mispredicted <= _GEN_2781;
      end
    end else begin
      T_26182_7_stat_btb_mispredicted <= _GEN_2781;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 406:72]
        T_26182_7_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_7_stat_bpd_made_pred <= _GEN_2805;
      end
    end else begin
      T_26182_7_stat_bpd_made_pred <= _GEN_2805;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 405:72]
        T_26182_7_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_7_stat_bpd_mispredicted <= _GEN_2829;
      end
    end else begin
      T_26182_7_stat_bpd_mispredicted <= _GEN_2829;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h7 == T_28605) begin // @[rob.scala 531:53]
        T_26182_7_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_7_debug_wdata <= _GEN_10267;
      end
    end else begin
      T_26182_7_debug_wdata <= _GEN_10267;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_7_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_8_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_8_inst <= _GEN_8228;
      end
    end else begin
      T_26182_8_inst <= _GEN_8228;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30280) begin // @[rob.scala 490:10]
      T_26182_8_br_mask <= T_30282; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 402:72]
        T_26182_8_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_8_stat_brjmp_mispredicted <= _GEN_2734;
      end
    end else begin
      T_26182_8_stat_brjmp_mispredicted <= _GEN_2734;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 404:72]
        T_26182_8_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_8_stat_btb_made_pred <= _GEN_2758;
      end
    end else begin
      T_26182_8_stat_btb_made_pred <= _GEN_2758;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 403:72]
        T_26182_8_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_8_stat_btb_mispredicted <= _GEN_2782;
      end
    end else begin
      T_26182_8_stat_btb_mispredicted <= _GEN_2782;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 406:72]
        T_26182_8_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_8_stat_bpd_made_pred <= _GEN_2806;
      end
    end else begin
      T_26182_8_stat_bpd_made_pred <= _GEN_2806;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 405:72]
        T_26182_8_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_8_stat_bpd_mispredicted <= _GEN_2830;
      end
    end else begin
      T_26182_8_stat_bpd_mispredicted <= _GEN_2830;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h8 == T_28605) begin // @[rob.scala 531:53]
        T_26182_8_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_8_debug_wdata <= _GEN_10268;
      end
    end else begin
      T_26182_8_debug_wdata <= _GEN_10268;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_8_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_9_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_9_inst <= _GEN_8229;
      end
    end else begin
      T_26182_9_inst <= _GEN_8229;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30382) begin // @[rob.scala 490:10]
      T_26182_9_br_mask <= T_30384; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 402:72]
        T_26182_9_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_9_stat_brjmp_mispredicted <= _GEN_2735;
      end
    end else begin
      T_26182_9_stat_brjmp_mispredicted <= _GEN_2735;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 404:72]
        T_26182_9_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_9_stat_btb_made_pred <= _GEN_2759;
      end
    end else begin
      T_26182_9_stat_btb_made_pred <= _GEN_2759;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 403:72]
        T_26182_9_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_9_stat_btb_mispredicted <= _GEN_2783;
      end
    end else begin
      T_26182_9_stat_btb_mispredicted <= _GEN_2783;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 406:72]
        T_26182_9_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_9_stat_bpd_made_pred <= _GEN_2807;
      end
    end else begin
      T_26182_9_stat_bpd_made_pred <= _GEN_2807;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 405:72]
        T_26182_9_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_9_stat_bpd_mispredicted <= _GEN_2831;
      end
    end else begin
      T_26182_9_stat_bpd_mispredicted <= _GEN_2831;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h9 == T_28605) begin // @[rob.scala 531:53]
        T_26182_9_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_9_debug_wdata <= _GEN_10269;
      end
    end else begin
      T_26182_9_debug_wdata <= _GEN_10269;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_9_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'ha == rob_tail) begin // @[rob.scala 519:33]
        T_26182_10_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_10_inst <= _GEN_8230;
      end
    end else begin
      T_26182_10_inst <= _GEN_8230;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30484) begin // @[rob.scala 490:10]
      T_26182_10_br_mask <= T_30486; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 402:72]
        T_26182_10_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_10_stat_brjmp_mispredicted <= _GEN_2736;
      end
    end else begin
      T_26182_10_stat_brjmp_mispredicted <= _GEN_2736;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 404:72]
        T_26182_10_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_10_stat_btb_made_pred <= _GEN_2760;
      end
    end else begin
      T_26182_10_stat_btb_made_pred <= _GEN_2760;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 403:72]
        T_26182_10_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_10_stat_btb_mispredicted <= _GEN_2784;
      end
    end else begin
      T_26182_10_stat_btb_mispredicted <= _GEN_2784;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 406:72]
        T_26182_10_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_10_stat_bpd_made_pred <= _GEN_2808;
      end
    end else begin
      T_26182_10_stat_bpd_made_pred <= _GEN_2808;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 405:72]
        T_26182_10_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_10_stat_bpd_mispredicted <= _GEN_2832;
      end
    end else begin
      T_26182_10_stat_bpd_mispredicted <= _GEN_2832;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'ha == T_28605) begin // @[rob.scala 531:53]
        T_26182_10_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_10_debug_wdata <= _GEN_10270;
      end
    end else begin
      T_26182_10_debug_wdata <= _GEN_10270;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_26182_10_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'hb == rob_tail) begin // @[rob.scala 519:33]
        T_26182_11_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_11_inst <= _GEN_8231;
      end
    end else begin
      T_26182_11_inst <= _GEN_8231;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30586) begin // @[rob.scala 490:10]
      T_26182_11_br_mask <= T_30588; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 402:72]
        T_26182_11_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_11_stat_brjmp_mispredicted <= _GEN_2737;
      end
    end else begin
      T_26182_11_stat_brjmp_mispredicted <= _GEN_2737;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 404:72]
        T_26182_11_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_11_stat_btb_made_pred <= _GEN_2761;
      end
    end else begin
      T_26182_11_stat_btb_made_pred <= _GEN_2761;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 403:72]
        T_26182_11_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_11_stat_btb_mispredicted <= _GEN_2785;
      end
    end else begin
      T_26182_11_stat_btb_mispredicted <= _GEN_2785;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 406:72]
        T_26182_11_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_11_stat_bpd_made_pred <= _GEN_2809;
      end
    end else begin
      T_26182_11_stat_bpd_made_pred <= _GEN_2809;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 405:72]
        T_26182_11_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_11_stat_bpd_mispredicted <= _GEN_2833;
      end
    end else begin
      T_26182_11_stat_bpd_mispredicted <= _GEN_2833;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'hb == T_28605) begin // @[rob.scala 531:53]
        T_26182_11_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_11_debug_wdata <= _GEN_10271;
      end
    end else begin
      T_26182_11_debug_wdata <= _GEN_10271;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_26182_11_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'hc == rob_tail) begin // @[rob.scala 519:33]
        T_26182_12_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_12_inst <= _GEN_8232;
      end
    end else begin
      T_26182_12_inst <= _GEN_8232;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30688) begin // @[rob.scala 490:10]
      T_26182_12_br_mask <= T_30690; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 402:72]
        T_26182_12_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_12_stat_brjmp_mispredicted <= _GEN_2738;
      end
    end else begin
      T_26182_12_stat_brjmp_mispredicted <= _GEN_2738;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 404:72]
        T_26182_12_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_12_stat_btb_made_pred <= _GEN_2762;
      end
    end else begin
      T_26182_12_stat_btb_made_pred <= _GEN_2762;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 403:72]
        T_26182_12_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_12_stat_btb_mispredicted <= _GEN_2786;
      end
    end else begin
      T_26182_12_stat_btb_mispredicted <= _GEN_2786;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 406:72]
        T_26182_12_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_12_stat_bpd_made_pred <= _GEN_2810;
      end
    end else begin
      T_26182_12_stat_bpd_made_pred <= _GEN_2810;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 405:72]
        T_26182_12_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_12_stat_bpd_mispredicted <= _GEN_2834;
      end
    end else begin
      T_26182_12_stat_bpd_mispredicted <= _GEN_2834;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'hc == T_28605) begin // @[rob.scala 531:53]
        T_26182_12_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_12_debug_wdata <= _GEN_10272;
      end
    end else begin
      T_26182_12_debug_wdata <= _GEN_10272;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_26182_12_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'hd == rob_tail) begin // @[rob.scala 519:33]
        T_26182_13_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_13_inst <= _GEN_8233;
      end
    end else begin
      T_26182_13_inst <= _GEN_8233;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30790) begin // @[rob.scala 490:10]
      T_26182_13_br_mask <= T_30792; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 402:72]
        T_26182_13_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_13_stat_brjmp_mispredicted <= _GEN_2739;
      end
    end else begin
      T_26182_13_stat_brjmp_mispredicted <= _GEN_2739;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 404:72]
        T_26182_13_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_13_stat_btb_made_pred <= _GEN_2763;
      end
    end else begin
      T_26182_13_stat_btb_made_pred <= _GEN_2763;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 403:72]
        T_26182_13_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_13_stat_btb_mispredicted <= _GEN_2787;
      end
    end else begin
      T_26182_13_stat_btb_mispredicted <= _GEN_2787;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 406:72]
        T_26182_13_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_13_stat_bpd_made_pred <= _GEN_2811;
      end
    end else begin
      T_26182_13_stat_bpd_made_pred <= _GEN_2811;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 405:72]
        T_26182_13_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_13_stat_bpd_mispredicted <= _GEN_2835;
      end
    end else begin
      T_26182_13_stat_bpd_mispredicted <= _GEN_2835;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'hd == T_28605) begin // @[rob.scala 531:53]
        T_26182_13_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_13_debug_wdata <= _GEN_10273;
      end
    end else begin
      T_26182_13_debug_wdata <= _GEN_10273;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_26182_13_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'he == rob_tail) begin // @[rob.scala 519:33]
        T_26182_14_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_14_inst <= _GEN_8234;
      end
    end else begin
      T_26182_14_inst <= _GEN_8234;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30892) begin // @[rob.scala 490:10]
      T_26182_14_br_mask <= T_30894; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 402:72]
        T_26182_14_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_14_stat_brjmp_mispredicted <= _GEN_2740;
      end
    end else begin
      T_26182_14_stat_brjmp_mispredicted <= _GEN_2740;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 404:72]
        T_26182_14_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_14_stat_btb_made_pred <= _GEN_2764;
      end
    end else begin
      T_26182_14_stat_btb_made_pred <= _GEN_2764;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 403:72]
        T_26182_14_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_14_stat_btb_mispredicted <= _GEN_2788;
      end
    end else begin
      T_26182_14_stat_btb_mispredicted <= _GEN_2788;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 406:72]
        T_26182_14_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_14_stat_bpd_made_pred <= _GEN_2812;
      end
    end else begin
      T_26182_14_stat_bpd_made_pred <= _GEN_2812;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 405:72]
        T_26182_14_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_14_stat_bpd_mispredicted <= _GEN_2836;
      end
    end else begin
      T_26182_14_stat_bpd_mispredicted <= _GEN_2836;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'he == T_28605) begin // @[rob.scala 531:53]
        T_26182_14_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_14_debug_wdata <= _GEN_10274;
      end
    end else begin
      T_26182_14_debug_wdata <= _GEN_10274;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_26182_14_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'hf == rob_tail) begin // @[rob.scala 519:33]
        T_26182_15_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_15_inst <= _GEN_8235;
      end
    end else begin
      T_26182_15_inst <= _GEN_8235;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_30994) begin // @[rob.scala 490:10]
      T_26182_15_br_mask <= T_30996; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 402:72]
        T_26182_15_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_15_stat_brjmp_mispredicted <= _GEN_2741;
      end
    end else begin
      T_26182_15_stat_brjmp_mispredicted <= _GEN_2741;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 404:72]
        T_26182_15_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_15_stat_btb_made_pred <= _GEN_2765;
      end
    end else begin
      T_26182_15_stat_btb_made_pred <= _GEN_2765;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 403:72]
        T_26182_15_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_15_stat_btb_mispredicted <= _GEN_2789;
      end
    end else begin
      T_26182_15_stat_btb_mispredicted <= _GEN_2789;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 406:72]
        T_26182_15_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_15_stat_bpd_made_pred <= _GEN_2813;
      end
    end else begin
      T_26182_15_stat_bpd_made_pred <= _GEN_2813;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 405:72]
        T_26182_15_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_15_stat_bpd_mispredicted <= _GEN_2837;
      end
    end else begin
      T_26182_15_stat_bpd_mispredicted <= _GEN_2837;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'hf == T_28605) begin // @[rob.scala 531:53]
        T_26182_15_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_15_debug_wdata <= _GEN_10275;
      end
    end else begin
      T_26182_15_debug_wdata <= _GEN_10275;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_26182_15_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_16_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_16_inst <= _GEN_8236;
      end
    end else begin
      T_26182_16_inst <= _GEN_8236;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31096) begin // @[rob.scala 490:10]
      T_26182_16_br_mask <= T_31098; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 402:72]
        T_26182_16_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_16_stat_brjmp_mispredicted <= _GEN_2742;
      end
    end else begin
      T_26182_16_stat_brjmp_mispredicted <= _GEN_2742;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 404:72]
        T_26182_16_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_16_stat_btb_made_pred <= _GEN_2766;
      end
    end else begin
      T_26182_16_stat_btb_made_pred <= _GEN_2766;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 403:72]
        T_26182_16_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_16_stat_btb_mispredicted <= _GEN_2790;
      end
    end else begin
      T_26182_16_stat_btb_mispredicted <= _GEN_2790;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 406:72]
        T_26182_16_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_16_stat_bpd_made_pred <= _GEN_2814;
      end
    end else begin
      T_26182_16_stat_bpd_made_pred <= _GEN_2814;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 405:72]
        T_26182_16_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_16_stat_bpd_mispredicted <= _GEN_2838;
      end
    end else begin
      T_26182_16_stat_bpd_mispredicted <= _GEN_2838;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h10 == T_28605) begin // @[rob.scala 531:53]
        T_26182_16_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_16_debug_wdata <= _GEN_10276;
      end
    end else begin
      T_26182_16_debug_wdata <= _GEN_10276;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_16_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_17_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_17_inst <= _GEN_8237;
      end
    end else begin
      T_26182_17_inst <= _GEN_8237;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31198) begin // @[rob.scala 490:10]
      T_26182_17_br_mask <= T_31200; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 402:72]
        T_26182_17_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_17_stat_brjmp_mispredicted <= _GEN_2743;
      end
    end else begin
      T_26182_17_stat_brjmp_mispredicted <= _GEN_2743;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 404:72]
        T_26182_17_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_17_stat_btb_made_pred <= _GEN_2767;
      end
    end else begin
      T_26182_17_stat_btb_made_pred <= _GEN_2767;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 403:72]
        T_26182_17_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_17_stat_btb_mispredicted <= _GEN_2791;
      end
    end else begin
      T_26182_17_stat_btb_mispredicted <= _GEN_2791;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 406:72]
        T_26182_17_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_17_stat_bpd_made_pred <= _GEN_2815;
      end
    end else begin
      T_26182_17_stat_bpd_made_pred <= _GEN_2815;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 405:72]
        T_26182_17_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_17_stat_bpd_mispredicted <= _GEN_2839;
      end
    end else begin
      T_26182_17_stat_bpd_mispredicted <= _GEN_2839;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h11 == T_28605) begin // @[rob.scala 531:53]
        T_26182_17_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_17_debug_wdata <= _GEN_10277;
      end
    end else begin
      T_26182_17_debug_wdata <= _GEN_10277;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_17_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_18_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_18_inst <= _GEN_8238;
      end
    end else begin
      T_26182_18_inst <= _GEN_8238;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31300) begin // @[rob.scala 490:10]
      T_26182_18_br_mask <= T_31302; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 402:72]
        T_26182_18_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_18_stat_brjmp_mispredicted <= _GEN_2744;
      end
    end else begin
      T_26182_18_stat_brjmp_mispredicted <= _GEN_2744;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 404:72]
        T_26182_18_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_18_stat_btb_made_pred <= _GEN_2768;
      end
    end else begin
      T_26182_18_stat_btb_made_pred <= _GEN_2768;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 403:72]
        T_26182_18_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_18_stat_btb_mispredicted <= _GEN_2792;
      end
    end else begin
      T_26182_18_stat_btb_mispredicted <= _GEN_2792;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 406:72]
        T_26182_18_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_18_stat_bpd_made_pred <= _GEN_2816;
      end
    end else begin
      T_26182_18_stat_bpd_made_pred <= _GEN_2816;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 405:72]
        T_26182_18_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_18_stat_bpd_mispredicted <= _GEN_2840;
      end
    end else begin
      T_26182_18_stat_bpd_mispredicted <= _GEN_2840;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h12 == T_28605) begin // @[rob.scala 531:53]
        T_26182_18_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_18_debug_wdata <= _GEN_10278;
      end
    end else begin
      T_26182_18_debug_wdata <= _GEN_10278;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_18_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_19_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_19_inst <= _GEN_8239;
      end
    end else begin
      T_26182_19_inst <= _GEN_8239;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31402) begin // @[rob.scala 490:10]
      T_26182_19_br_mask <= T_31404; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 402:72]
        T_26182_19_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_19_stat_brjmp_mispredicted <= _GEN_2745;
      end
    end else begin
      T_26182_19_stat_brjmp_mispredicted <= _GEN_2745;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 404:72]
        T_26182_19_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_19_stat_btb_made_pred <= _GEN_2769;
      end
    end else begin
      T_26182_19_stat_btb_made_pred <= _GEN_2769;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 403:72]
        T_26182_19_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_19_stat_btb_mispredicted <= _GEN_2793;
      end
    end else begin
      T_26182_19_stat_btb_mispredicted <= _GEN_2793;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 406:72]
        T_26182_19_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_19_stat_bpd_made_pred <= _GEN_2817;
      end
    end else begin
      T_26182_19_stat_bpd_made_pred <= _GEN_2817;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 405:72]
        T_26182_19_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_19_stat_bpd_mispredicted <= _GEN_2841;
      end
    end else begin
      T_26182_19_stat_bpd_mispredicted <= _GEN_2841;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h13 == T_28605) begin // @[rob.scala 531:53]
        T_26182_19_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_19_debug_wdata <= _GEN_10279;
      end
    end else begin
      T_26182_19_debug_wdata <= _GEN_10279;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_19_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_20_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_20_inst <= _GEN_8240;
      end
    end else begin
      T_26182_20_inst <= _GEN_8240;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31504) begin // @[rob.scala 490:10]
      T_26182_20_br_mask <= T_31506; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 402:72]
        T_26182_20_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_20_stat_brjmp_mispredicted <= _GEN_2746;
      end
    end else begin
      T_26182_20_stat_brjmp_mispredicted <= _GEN_2746;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 404:72]
        T_26182_20_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_20_stat_btb_made_pred <= _GEN_2770;
      end
    end else begin
      T_26182_20_stat_btb_made_pred <= _GEN_2770;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 403:72]
        T_26182_20_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_20_stat_btb_mispredicted <= _GEN_2794;
      end
    end else begin
      T_26182_20_stat_btb_mispredicted <= _GEN_2794;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 406:72]
        T_26182_20_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_20_stat_bpd_made_pred <= _GEN_2818;
      end
    end else begin
      T_26182_20_stat_bpd_made_pred <= _GEN_2818;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 405:72]
        T_26182_20_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_20_stat_bpd_mispredicted <= _GEN_2842;
      end
    end else begin
      T_26182_20_stat_bpd_mispredicted <= _GEN_2842;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h14 == T_28605) begin // @[rob.scala 531:53]
        T_26182_20_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_20_debug_wdata <= _GEN_10280;
      end
    end else begin
      T_26182_20_debug_wdata <= _GEN_10280;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_20_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_21_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_21_inst <= _GEN_8241;
      end
    end else begin
      T_26182_21_inst <= _GEN_8241;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31606) begin // @[rob.scala 490:10]
      T_26182_21_br_mask <= T_31608; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 402:72]
        T_26182_21_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_21_stat_brjmp_mispredicted <= _GEN_2747;
      end
    end else begin
      T_26182_21_stat_brjmp_mispredicted <= _GEN_2747;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 404:72]
        T_26182_21_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_21_stat_btb_made_pred <= _GEN_2771;
      end
    end else begin
      T_26182_21_stat_btb_made_pred <= _GEN_2771;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 403:72]
        T_26182_21_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_21_stat_btb_mispredicted <= _GEN_2795;
      end
    end else begin
      T_26182_21_stat_btb_mispredicted <= _GEN_2795;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 406:72]
        T_26182_21_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_21_stat_bpd_made_pred <= _GEN_2819;
      end
    end else begin
      T_26182_21_stat_bpd_made_pred <= _GEN_2819;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 405:72]
        T_26182_21_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_21_stat_bpd_mispredicted <= _GEN_2843;
      end
    end else begin
      T_26182_21_stat_bpd_mispredicted <= _GEN_2843;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h15 == T_28605) begin // @[rob.scala 531:53]
        T_26182_21_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_21_debug_wdata <= _GEN_10281;
      end
    end else begin
      T_26182_21_debug_wdata <= _GEN_10281;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_21_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_22_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_22_inst <= _GEN_8242;
      end
    end else begin
      T_26182_22_inst <= _GEN_8242;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31708) begin // @[rob.scala 490:10]
      T_26182_22_br_mask <= T_31710; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 402:72]
        T_26182_22_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_22_stat_brjmp_mispredicted <= _GEN_2748;
      end
    end else begin
      T_26182_22_stat_brjmp_mispredicted <= _GEN_2748;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 404:72]
        T_26182_22_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_22_stat_btb_made_pred <= _GEN_2772;
      end
    end else begin
      T_26182_22_stat_btb_made_pred <= _GEN_2772;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 403:72]
        T_26182_22_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_22_stat_btb_mispredicted <= _GEN_2796;
      end
    end else begin
      T_26182_22_stat_btb_mispredicted <= _GEN_2796;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 406:72]
        T_26182_22_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_22_stat_bpd_made_pred <= _GEN_2820;
      end
    end else begin
      T_26182_22_stat_bpd_made_pred <= _GEN_2820;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 405:72]
        T_26182_22_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_22_stat_bpd_mispredicted <= _GEN_2844;
      end
    end else begin
      T_26182_22_stat_bpd_mispredicted <= _GEN_2844;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h16 == T_28605) begin // @[rob.scala 531:53]
        T_26182_22_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_22_debug_wdata <= _GEN_10282;
      end
    end else begin
      T_26182_22_debug_wdata <= _GEN_10282;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_22_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_valid <= io_dis_uops_0_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_iw_state <= io_dis_uops_0_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_uopc <= io_dis_uops_0_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_32082) begin // @[rob.scala 518:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 519:33]
        T_26182_23_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_26182_23_inst <= _GEN_8243;
      end
    end else begin
      T_26182_23_inst <= _GEN_8243;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_pc <= io_dis_uops_0_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_fu_code <= io_dis_uops_0_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_br_type <= io_dis_uops_0_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_is_load <= io_dis_uops_0_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ctrl_is_std <= io_dis_uops_0_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_wakeup_delay <= io_dis_uops_0_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_allocate_brtag <= io_dis_uops_0_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_jump <= io_dis_uops_0_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_jal <= io_dis_uops_0_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_ret <= io_dis_uops_0_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_call <= io_dis_uops_0_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_31810) begin // @[rob.scala 490:10]
      T_26182_23_br_mask <= T_31812; // @[rob.scala 492:32]
    end else if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_mask <= io_dis_uops_0_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_tag <= io_dis_uops_0_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 402:72]
        T_26182_23_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_26182_23_stat_brjmp_mispredicted <= _GEN_2749;
      end
    end else begin
      T_26182_23_stat_brjmp_mispredicted <= _GEN_2749;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 404:72]
        T_26182_23_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_26182_23_stat_btb_made_pred <= _GEN_2773;
      end
    end else begin
      T_26182_23_stat_btb_made_pred <= _GEN_2773;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 403:72]
        T_26182_23_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_26182_23_stat_btb_mispredicted <= _GEN_2797;
      end
    end else begin
      T_26182_23_stat_btb_mispredicted <= _GEN_2797;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 406:72]
        T_26182_23_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_26182_23_stat_bpd_made_pred <= _GEN_2821;
      end
    end else begin
      T_26182_23_stat_bpd_made_pred <= _GEN_2821;
    end
    if (T_28623) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 405:72]
        T_26182_23_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_26182_23_stat_bpd_mispredicted <= _GEN_2845;
      end
    end else begin
      T_26182_23_stat_bpd_mispredicted <= _GEN_2845;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_imm_packed <= io_dis_uops_0_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_csr_addr <= io_dis_uops_0_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_rob_idx <= io_dis_uops_0_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ldq_idx <= io_dis_uops_0_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_stq_idx <= io_dis_uops_0_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_brob_idx <= io_dis_uops_0_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_pdst <= io_dis_uops_0_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_pop1 <= io_dis_uops_0_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_pop2 <= io_dis_uops_0_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_pop3 <= io_dis_uops_0_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_prs1_busy <= io_dis_uops_0_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_prs2_busy <= io_dis_uops_0_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_prs3_busy <= io_dis_uops_0_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_stale_pdst <= io_dis_uops_0_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_exception <= io_dis_uops_0_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_exc_cause <= io_dis_uops_0_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_bypassable <= io_dis_uops_0_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_mem_cmd <= io_dis_uops_0_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_mem_typ <= io_dis_uops_0_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_fence <= io_dis_uops_0_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_fencei <= io_dis_uops_0_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_store <= io_dis_uops_0_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_amo <= io_dis_uops_0_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_load <= io_dis_uops_0_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_is_unique <= io_dis_uops_0_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_flush_on_commit <= io_dis_uops_0_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ldst <= io_dis_uops_0_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_lrs1 <= io_dis_uops_0_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_lrs2 <= io_dis_uops_0_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_lrs3 <= io_dis_uops_0_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_ldst_val <= io_dis_uops_0_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_dst_rtype <= io_dis_uops_0_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_lrs1_rtype <= io_dis_uops_0_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_lrs2_rtype <= io_dis_uops_0_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_frs3_en <= io_dis_uops_0_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_fp_val <= io_dis_uops_0_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_fp_single <= io_dis_uops_0_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_xcpt_if <= io_dis_uops_0_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_replay_if <= io_dis_uops_0_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_32579) begin // @[rob.scala 530:10]
      if (6'h17 == T_28605) begin // @[rob.scala 531:53]
        T_26182_23_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_26182_23_debug_wdata <= _GEN_10283;
      end
    end else begin
      T_26182_23_debug_wdata <= _GEN_10283;
    end
    if (io_dis_valids_0) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_26182_23_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_0_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_0_inst <= _GEN_22363;
      end
    end else begin
      T_38110_0_inst <= _GEN_22363;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_41392) begin // @[rob.scala 490:10]
      T_38110_0_br_mask <= T_41394; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 402:72]
        T_38110_0_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_0_stat_brjmp_mispredicted <= _GEN_16869;
      end
    end else begin
      T_38110_0_stat_brjmp_mispredicted <= _GEN_16869;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 404:72]
        T_38110_0_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_0_stat_btb_made_pred <= _GEN_16893;
      end
    end else begin
      T_38110_0_stat_btb_made_pred <= _GEN_16893;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 403:72]
        T_38110_0_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_0_stat_btb_mispredicted <= _GEN_16917;
      end
    end else begin
      T_38110_0_stat_btb_mispredicted <= _GEN_16917;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 406:72]
        T_38110_0_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_0_stat_bpd_made_pred <= _GEN_16941;
      end
    end else begin
      T_38110_0_stat_bpd_made_pred <= _GEN_16941;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h0 == T_28625) begin // @[rob.scala 405:72]
        T_38110_0_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_0_stat_bpd_mispredicted <= _GEN_16965;
      end
    end else begin
      T_38110_0_stat_bpd_mispredicted <= _GEN_16965;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h0 == T_28605) begin // @[rob.scala 531:53]
        T_38110_0_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_0_debug_wdata <= _GEN_24403;
      end
    end else begin
      T_38110_0_debug_wdata <= _GEN_24403;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h0 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_0_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_1_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_1_inst <= _GEN_22364;
      end
    end else begin
      T_38110_1_inst <= _GEN_22364;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_41494) begin // @[rob.scala 490:10]
      T_38110_1_br_mask <= T_41496; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 402:72]
        T_38110_1_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_1_stat_brjmp_mispredicted <= _GEN_16870;
      end
    end else begin
      T_38110_1_stat_brjmp_mispredicted <= _GEN_16870;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 404:72]
        T_38110_1_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_1_stat_btb_made_pred <= _GEN_16894;
      end
    end else begin
      T_38110_1_stat_btb_made_pred <= _GEN_16894;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 403:72]
        T_38110_1_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_1_stat_btb_mispredicted <= _GEN_16918;
      end
    end else begin
      T_38110_1_stat_btb_mispredicted <= _GEN_16918;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 406:72]
        T_38110_1_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_1_stat_bpd_made_pred <= _GEN_16942;
      end
    end else begin
      T_38110_1_stat_bpd_made_pred <= _GEN_16942;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h1 == T_28625) begin // @[rob.scala 405:72]
        T_38110_1_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_1_stat_bpd_mispredicted <= _GEN_16966;
      end
    end else begin
      T_38110_1_stat_bpd_mispredicted <= _GEN_16966;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h1 == T_28605) begin // @[rob.scala 531:53]
        T_38110_1_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_1_debug_wdata <= _GEN_24404;
      end
    end else begin
      T_38110_1_debug_wdata <= _GEN_24404;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h1 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_1_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_2_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_2_inst <= _GEN_22365;
      end
    end else begin
      T_38110_2_inst <= _GEN_22365;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_41596) begin // @[rob.scala 490:10]
      T_38110_2_br_mask <= T_41598; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 402:72]
        T_38110_2_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_2_stat_brjmp_mispredicted <= _GEN_16871;
      end
    end else begin
      T_38110_2_stat_brjmp_mispredicted <= _GEN_16871;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 404:72]
        T_38110_2_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_2_stat_btb_made_pred <= _GEN_16895;
      end
    end else begin
      T_38110_2_stat_btb_made_pred <= _GEN_16895;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 403:72]
        T_38110_2_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_2_stat_btb_mispredicted <= _GEN_16919;
      end
    end else begin
      T_38110_2_stat_btb_mispredicted <= _GEN_16919;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 406:72]
        T_38110_2_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_2_stat_bpd_made_pred <= _GEN_16943;
      end
    end else begin
      T_38110_2_stat_bpd_made_pred <= _GEN_16943;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h2 == T_28625) begin // @[rob.scala 405:72]
        T_38110_2_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_2_stat_bpd_mispredicted <= _GEN_16967;
      end
    end else begin
      T_38110_2_stat_bpd_mispredicted <= _GEN_16967;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h2 == T_28605) begin // @[rob.scala 531:53]
        T_38110_2_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_2_debug_wdata <= _GEN_24405;
      end
    end else begin
      T_38110_2_debug_wdata <= _GEN_24405;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h2 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_2_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_3_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_3_inst <= _GEN_22366;
      end
    end else begin
      T_38110_3_inst <= _GEN_22366;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_41698) begin // @[rob.scala 490:10]
      T_38110_3_br_mask <= T_41700; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 402:72]
        T_38110_3_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_3_stat_brjmp_mispredicted <= _GEN_16872;
      end
    end else begin
      T_38110_3_stat_brjmp_mispredicted <= _GEN_16872;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 404:72]
        T_38110_3_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_3_stat_btb_made_pred <= _GEN_16896;
      end
    end else begin
      T_38110_3_stat_btb_made_pred <= _GEN_16896;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 403:72]
        T_38110_3_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_3_stat_btb_mispredicted <= _GEN_16920;
      end
    end else begin
      T_38110_3_stat_btb_mispredicted <= _GEN_16920;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 406:72]
        T_38110_3_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_3_stat_bpd_made_pred <= _GEN_16944;
      end
    end else begin
      T_38110_3_stat_bpd_made_pred <= _GEN_16944;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h3 == T_28625) begin // @[rob.scala 405:72]
        T_38110_3_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_3_stat_bpd_mispredicted <= _GEN_16968;
      end
    end else begin
      T_38110_3_stat_bpd_mispredicted <= _GEN_16968;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h3 == T_28605) begin // @[rob.scala 531:53]
        T_38110_3_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_3_debug_wdata <= _GEN_24406;
      end
    end else begin
      T_38110_3_debug_wdata <= _GEN_24406;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h3 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_3_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_4_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_4_inst <= _GEN_22367;
      end
    end else begin
      T_38110_4_inst <= _GEN_22367;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_41800) begin // @[rob.scala 490:10]
      T_38110_4_br_mask <= T_41802; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 402:72]
        T_38110_4_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_4_stat_brjmp_mispredicted <= _GEN_16873;
      end
    end else begin
      T_38110_4_stat_brjmp_mispredicted <= _GEN_16873;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 404:72]
        T_38110_4_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_4_stat_btb_made_pred <= _GEN_16897;
      end
    end else begin
      T_38110_4_stat_btb_made_pred <= _GEN_16897;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 403:72]
        T_38110_4_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_4_stat_btb_mispredicted <= _GEN_16921;
      end
    end else begin
      T_38110_4_stat_btb_mispredicted <= _GEN_16921;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 406:72]
        T_38110_4_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_4_stat_bpd_made_pred <= _GEN_16945;
      end
    end else begin
      T_38110_4_stat_bpd_made_pred <= _GEN_16945;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h4 == T_28625) begin // @[rob.scala 405:72]
        T_38110_4_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_4_stat_bpd_mispredicted <= _GEN_16969;
      end
    end else begin
      T_38110_4_stat_bpd_mispredicted <= _GEN_16969;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h4 == T_28605) begin // @[rob.scala 531:53]
        T_38110_4_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_4_debug_wdata <= _GEN_24407;
      end
    end else begin
      T_38110_4_debug_wdata <= _GEN_24407;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h4 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_4_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_5_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_5_inst <= _GEN_22368;
      end
    end else begin
      T_38110_5_inst <= _GEN_22368;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_41902) begin // @[rob.scala 490:10]
      T_38110_5_br_mask <= T_41904; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 402:72]
        T_38110_5_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_5_stat_brjmp_mispredicted <= _GEN_16874;
      end
    end else begin
      T_38110_5_stat_brjmp_mispredicted <= _GEN_16874;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 404:72]
        T_38110_5_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_5_stat_btb_made_pred <= _GEN_16898;
      end
    end else begin
      T_38110_5_stat_btb_made_pred <= _GEN_16898;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 403:72]
        T_38110_5_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_5_stat_btb_mispredicted <= _GEN_16922;
      end
    end else begin
      T_38110_5_stat_btb_mispredicted <= _GEN_16922;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 406:72]
        T_38110_5_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_5_stat_bpd_made_pred <= _GEN_16946;
      end
    end else begin
      T_38110_5_stat_bpd_made_pred <= _GEN_16946;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h5 == T_28625) begin // @[rob.scala 405:72]
        T_38110_5_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_5_stat_bpd_mispredicted <= _GEN_16970;
      end
    end else begin
      T_38110_5_stat_bpd_mispredicted <= _GEN_16970;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h5 == T_28605) begin // @[rob.scala 531:53]
        T_38110_5_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_5_debug_wdata <= _GEN_24408;
      end
    end else begin
      T_38110_5_debug_wdata <= _GEN_24408;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h5 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_5_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_6_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_6_inst <= _GEN_22369;
      end
    end else begin
      T_38110_6_inst <= _GEN_22369;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42004) begin // @[rob.scala 490:10]
      T_38110_6_br_mask <= T_42006; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 402:72]
        T_38110_6_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_6_stat_brjmp_mispredicted <= _GEN_16875;
      end
    end else begin
      T_38110_6_stat_brjmp_mispredicted <= _GEN_16875;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 404:72]
        T_38110_6_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_6_stat_btb_made_pred <= _GEN_16899;
      end
    end else begin
      T_38110_6_stat_btb_made_pred <= _GEN_16899;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 403:72]
        T_38110_6_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_6_stat_btb_mispredicted <= _GEN_16923;
      end
    end else begin
      T_38110_6_stat_btb_mispredicted <= _GEN_16923;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 406:72]
        T_38110_6_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_6_stat_bpd_made_pred <= _GEN_16947;
      end
    end else begin
      T_38110_6_stat_bpd_made_pred <= _GEN_16947;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h6 == T_28625) begin // @[rob.scala 405:72]
        T_38110_6_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_6_stat_bpd_mispredicted <= _GEN_16971;
      end
    end else begin
      T_38110_6_stat_bpd_mispredicted <= _GEN_16971;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h6 == T_28605) begin // @[rob.scala 531:53]
        T_38110_6_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_6_debug_wdata <= _GEN_24409;
      end
    end else begin
      T_38110_6_debug_wdata <= _GEN_24409;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h6 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_6_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_7_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_7_inst <= _GEN_22370;
      end
    end else begin
      T_38110_7_inst <= _GEN_22370;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42106) begin // @[rob.scala 490:10]
      T_38110_7_br_mask <= T_42108; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 402:72]
        T_38110_7_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_7_stat_brjmp_mispredicted <= _GEN_16876;
      end
    end else begin
      T_38110_7_stat_brjmp_mispredicted <= _GEN_16876;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 404:72]
        T_38110_7_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_7_stat_btb_made_pred <= _GEN_16900;
      end
    end else begin
      T_38110_7_stat_btb_made_pred <= _GEN_16900;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 403:72]
        T_38110_7_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_7_stat_btb_mispredicted <= _GEN_16924;
      end
    end else begin
      T_38110_7_stat_btb_mispredicted <= _GEN_16924;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 406:72]
        T_38110_7_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_7_stat_bpd_made_pred <= _GEN_16948;
      end
    end else begin
      T_38110_7_stat_bpd_made_pred <= _GEN_16948;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h7 == T_28625) begin // @[rob.scala 405:72]
        T_38110_7_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_7_stat_bpd_mispredicted <= _GEN_16972;
      end
    end else begin
      T_38110_7_stat_bpd_mispredicted <= _GEN_16972;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h7 == T_28605) begin // @[rob.scala 531:53]
        T_38110_7_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_7_debug_wdata <= _GEN_24410;
      end
    end else begin
      T_38110_7_debug_wdata <= _GEN_24410;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h7 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_7_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_8_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_8_inst <= _GEN_22371;
      end
    end else begin
      T_38110_8_inst <= _GEN_22371;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42208) begin // @[rob.scala 490:10]
      T_38110_8_br_mask <= T_42210; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 402:72]
        T_38110_8_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_8_stat_brjmp_mispredicted <= _GEN_16877;
      end
    end else begin
      T_38110_8_stat_brjmp_mispredicted <= _GEN_16877;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 404:72]
        T_38110_8_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_8_stat_btb_made_pred <= _GEN_16901;
      end
    end else begin
      T_38110_8_stat_btb_made_pred <= _GEN_16901;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 403:72]
        T_38110_8_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_8_stat_btb_mispredicted <= _GEN_16925;
      end
    end else begin
      T_38110_8_stat_btb_mispredicted <= _GEN_16925;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 406:72]
        T_38110_8_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_8_stat_bpd_made_pred <= _GEN_16949;
      end
    end else begin
      T_38110_8_stat_bpd_made_pred <= _GEN_16949;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h8 == T_28625) begin // @[rob.scala 405:72]
        T_38110_8_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_8_stat_bpd_mispredicted <= _GEN_16973;
      end
    end else begin
      T_38110_8_stat_bpd_mispredicted <= _GEN_16973;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h8 == T_28605) begin // @[rob.scala 531:53]
        T_38110_8_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_8_debug_wdata <= _GEN_24411;
      end
    end else begin
      T_38110_8_debug_wdata <= _GEN_24411;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h8 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_8_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_9_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_9_inst <= _GEN_22372;
      end
    end else begin
      T_38110_9_inst <= _GEN_22372;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42310) begin // @[rob.scala 490:10]
      T_38110_9_br_mask <= T_42312; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 402:72]
        T_38110_9_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_9_stat_brjmp_mispredicted <= _GEN_16878;
      end
    end else begin
      T_38110_9_stat_brjmp_mispredicted <= _GEN_16878;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 404:72]
        T_38110_9_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_9_stat_btb_made_pred <= _GEN_16902;
      end
    end else begin
      T_38110_9_stat_btb_made_pred <= _GEN_16902;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 403:72]
        T_38110_9_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_9_stat_btb_mispredicted <= _GEN_16926;
      end
    end else begin
      T_38110_9_stat_btb_mispredicted <= _GEN_16926;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 406:72]
        T_38110_9_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_9_stat_bpd_made_pred <= _GEN_16950;
      end
    end else begin
      T_38110_9_stat_bpd_made_pred <= _GEN_16950;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h9 == T_28625) begin // @[rob.scala 405:72]
        T_38110_9_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_9_stat_bpd_mispredicted <= _GEN_16974;
      end
    end else begin
      T_38110_9_stat_bpd_mispredicted <= _GEN_16974;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h9 == T_28605) begin // @[rob.scala 531:53]
        T_38110_9_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_9_debug_wdata <= _GEN_24412;
      end
    end else begin
      T_38110_9_debug_wdata <= _GEN_24412;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h9 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_9_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'ha == rob_tail) begin // @[rob.scala 519:33]
        T_38110_10_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_10_inst <= _GEN_22373;
      end
    end else begin
      T_38110_10_inst <= _GEN_22373;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42412) begin // @[rob.scala 490:10]
      T_38110_10_br_mask <= T_42414; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 402:72]
        T_38110_10_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_10_stat_brjmp_mispredicted <= _GEN_16879;
      end
    end else begin
      T_38110_10_stat_brjmp_mispredicted <= _GEN_16879;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 404:72]
        T_38110_10_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_10_stat_btb_made_pred <= _GEN_16903;
      end
    end else begin
      T_38110_10_stat_btb_made_pred <= _GEN_16903;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 403:72]
        T_38110_10_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_10_stat_btb_mispredicted <= _GEN_16927;
      end
    end else begin
      T_38110_10_stat_btb_mispredicted <= _GEN_16927;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 406:72]
        T_38110_10_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_10_stat_bpd_made_pred <= _GEN_16951;
      end
    end else begin
      T_38110_10_stat_bpd_made_pred <= _GEN_16951;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'ha == T_28625) begin // @[rob.scala 405:72]
        T_38110_10_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_10_stat_bpd_mispredicted <= _GEN_16975;
      end
    end else begin
      T_38110_10_stat_bpd_mispredicted <= _GEN_16975;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'ha == T_28605) begin // @[rob.scala 531:53]
        T_38110_10_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_10_debug_wdata <= _GEN_24413;
      end
    end else begin
      T_38110_10_debug_wdata <= _GEN_24413;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'ha == rob_tail) begin // @[rob.scala 350:34]
        T_38110_10_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'hb == rob_tail) begin // @[rob.scala 519:33]
        T_38110_11_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_11_inst <= _GEN_22374;
      end
    end else begin
      T_38110_11_inst <= _GEN_22374;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42514) begin // @[rob.scala 490:10]
      T_38110_11_br_mask <= T_42516; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 402:72]
        T_38110_11_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_11_stat_brjmp_mispredicted <= _GEN_16880;
      end
    end else begin
      T_38110_11_stat_brjmp_mispredicted <= _GEN_16880;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 404:72]
        T_38110_11_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_11_stat_btb_made_pred <= _GEN_16904;
      end
    end else begin
      T_38110_11_stat_btb_made_pred <= _GEN_16904;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 403:72]
        T_38110_11_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_11_stat_btb_mispredicted <= _GEN_16928;
      end
    end else begin
      T_38110_11_stat_btb_mispredicted <= _GEN_16928;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 406:72]
        T_38110_11_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_11_stat_bpd_made_pred <= _GEN_16952;
      end
    end else begin
      T_38110_11_stat_bpd_made_pred <= _GEN_16952;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hb == T_28625) begin // @[rob.scala 405:72]
        T_38110_11_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_11_stat_bpd_mispredicted <= _GEN_16976;
      end
    end else begin
      T_38110_11_stat_bpd_mispredicted <= _GEN_16976;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'hb == T_28605) begin // @[rob.scala 531:53]
        T_38110_11_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_11_debug_wdata <= _GEN_24414;
      end
    end else begin
      T_38110_11_debug_wdata <= _GEN_24414;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hb == rob_tail) begin // @[rob.scala 350:34]
        T_38110_11_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'hc == rob_tail) begin // @[rob.scala 519:33]
        T_38110_12_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_12_inst <= _GEN_22375;
      end
    end else begin
      T_38110_12_inst <= _GEN_22375;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42616) begin // @[rob.scala 490:10]
      T_38110_12_br_mask <= T_42618; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 402:72]
        T_38110_12_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_12_stat_brjmp_mispredicted <= _GEN_16881;
      end
    end else begin
      T_38110_12_stat_brjmp_mispredicted <= _GEN_16881;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 404:72]
        T_38110_12_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_12_stat_btb_made_pred <= _GEN_16905;
      end
    end else begin
      T_38110_12_stat_btb_made_pred <= _GEN_16905;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 403:72]
        T_38110_12_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_12_stat_btb_mispredicted <= _GEN_16929;
      end
    end else begin
      T_38110_12_stat_btb_mispredicted <= _GEN_16929;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 406:72]
        T_38110_12_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_12_stat_bpd_made_pred <= _GEN_16953;
      end
    end else begin
      T_38110_12_stat_bpd_made_pred <= _GEN_16953;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hc == T_28625) begin // @[rob.scala 405:72]
        T_38110_12_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_12_stat_bpd_mispredicted <= _GEN_16977;
      end
    end else begin
      T_38110_12_stat_bpd_mispredicted <= _GEN_16977;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'hc == T_28605) begin // @[rob.scala 531:53]
        T_38110_12_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_12_debug_wdata <= _GEN_24415;
      end
    end else begin
      T_38110_12_debug_wdata <= _GEN_24415;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hc == rob_tail) begin // @[rob.scala 350:34]
        T_38110_12_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'hd == rob_tail) begin // @[rob.scala 519:33]
        T_38110_13_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_13_inst <= _GEN_22376;
      end
    end else begin
      T_38110_13_inst <= _GEN_22376;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42718) begin // @[rob.scala 490:10]
      T_38110_13_br_mask <= T_42720; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 402:72]
        T_38110_13_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_13_stat_brjmp_mispredicted <= _GEN_16882;
      end
    end else begin
      T_38110_13_stat_brjmp_mispredicted <= _GEN_16882;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 404:72]
        T_38110_13_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_13_stat_btb_made_pred <= _GEN_16906;
      end
    end else begin
      T_38110_13_stat_btb_made_pred <= _GEN_16906;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 403:72]
        T_38110_13_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_13_stat_btb_mispredicted <= _GEN_16930;
      end
    end else begin
      T_38110_13_stat_btb_mispredicted <= _GEN_16930;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 406:72]
        T_38110_13_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_13_stat_bpd_made_pred <= _GEN_16954;
      end
    end else begin
      T_38110_13_stat_bpd_made_pred <= _GEN_16954;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hd == T_28625) begin // @[rob.scala 405:72]
        T_38110_13_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_13_stat_bpd_mispredicted <= _GEN_16978;
      end
    end else begin
      T_38110_13_stat_bpd_mispredicted <= _GEN_16978;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'hd == T_28605) begin // @[rob.scala 531:53]
        T_38110_13_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_13_debug_wdata <= _GEN_24416;
      end
    end else begin
      T_38110_13_debug_wdata <= _GEN_24416;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hd == rob_tail) begin // @[rob.scala 350:34]
        T_38110_13_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'he == rob_tail) begin // @[rob.scala 519:33]
        T_38110_14_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_14_inst <= _GEN_22377;
      end
    end else begin
      T_38110_14_inst <= _GEN_22377;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42820) begin // @[rob.scala 490:10]
      T_38110_14_br_mask <= T_42822; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 402:72]
        T_38110_14_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_14_stat_brjmp_mispredicted <= _GEN_16883;
      end
    end else begin
      T_38110_14_stat_brjmp_mispredicted <= _GEN_16883;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 404:72]
        T_38110_14_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_14_stat_btb_made_pred <= _GEN_16907;
      end
    end else begin
      T_38110_14_stat_btb_made_pred <= _GEN_16907;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 403:72]
        T_38110_14_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_14_stat_btb_mispredicted <= _GEN_16931;
      end
    end else begin
      T_38110_14_stat_btb_mispredicted <= _GEN_16931;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 406:72]
        T_38110_14_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_14_stat_bpd_made_pred <= _GEN_16955;
      end
    end else begin
      T_38110_14_stat_bpd_made_pred <= _GEN_16955;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'he == T_28625) begin // @[rob.scala 405:72]
        T_38110_14_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_14_stat_bpd_mispredicted <= _GEN_16979;
      end
    end else begin
      T_38110_14_stat_bpd_mispredicted <= _GEN_16979;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'he == T_28605) begin // @[rob.scala 531:53]
        T_38110_14_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_14_debug_wdata <= _GEN_24417;
      end
    end else begin
      T_38110_14_debug_wdata <= _GEN_24417;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'he == rob_tail) begin // @[rob.scala 350:34]
        T_38110_14_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'hf == rob_tail) begin // @[rob.scala 519:33]
        T_38110_15_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_15_inst <= _GEN_22378;
      end
    end else begin
      T_38110_15_inst <= _GEN_22378;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_42922) begin // @[rob.scala 490:10]
      T_38110_15_br_mask <= T_42924; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 402:72]
        T_38110_15_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_15_stat_brjmp_mispredicted <= _GEN_16884;
      end
    end else begin
      T_38110_15_stat_brjmp_mispredicted <= _GEN_16884;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 404:72]
        T_38110_15_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_15_stat_btb_made_pred <= _GEN_16908;
      end
    end else begin
      T_38110_15_stat_btb_made_pred <= _GEN_16908;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 403:72]
        T_38110_15_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_15_stat_btb_mispredicted <= _GEN_16932;
      end
    end else begin
      T_38110_15_stat_btb_mispredicted <= _GEN_16932;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 406:72]
        T_38110_15_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_15_stat_bpd_made_pred <= _GEN_16956;
      end
    end else begin
      T_38110_15_stat_bpd_made_pred <= _GEN_16956;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'hf == T_28625) begin // @[rob.scala 405:72]
        T_38110_15_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_15_stat_bpd_mispredicted <= _GEN_16980;
      end
    end else begin
      T_38110_15_stat_bpd_mispredicted <= _GEN_16980;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'hf == T_28605) begin // @[rob.scala 531:53]
        T_38110_15_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_15_debug_wdata <= _GEN_24418;
      end
    end else begin
      T_38110_15_debug_wdata <= _GEN_24418;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'hf == rob_tail) begin // @[rob.scala 350:34]
        T_38110_15_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_16_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_16_inst <= _GEN_22379;
      end
    end else begin
      T_38110_16_inst <= _GEN_22379;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43024) begin // @[rob.scala 490:10]
      T_38110_16_br_mask <= T_43026; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 402:72]
        T_38110_16_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_16_stat_brjmp_mispredicted <= _GEN_16885;
      end
    end else begin
      T_38110_16_stat_brjmp_mispredicted <= _GEN_16885;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 404:72]
        T_38110_16_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_16_stat_btb_made_pred <= _GEN_16909;
      end
    end else begin
      T_38110_16_stat_btb_made_pred <= _GEN_16909;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 403:72]
        T_38110_16_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_16_stat_btb_mispredicted <= _GEN_16933;
      end
    end else begin
      T_38110_16_stat_btb_mispredicted <= _GEN_16933;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 406:72]
        T_38110_16_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_16_stat_bpd_made_pred <= _GEN_16957;
      end
    end else begin
      T_38110_16_stat_bpd_made_pred <= _GEN_16957;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h10 == T_28625) begin // @[rob.scala 405:72]
        T_38110_16_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_16_stat_bpd_mispredicted <= _GEN_16981;
      end
    end else begin
      T_38110_16_stat_bpd_mispredicted <= _GEN_16981;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h10 == T_28605) begin // @[rob.scala 531:53]
        T_38110_16_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_16_debug_wdata <= _GEN_24419;
      end
    end else begin
      T_38110_16_debug_wdata <= _GEN_24419;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h10 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_16_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_17_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_17_inst <= _GEN_22380;
      end
    end else begin
      T_38110_17_inst <= _GEN_22380;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43126) begin // @[rob.scala 490:10]
      T_38110_17_br_mask <= T_43128; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 402:72]
        T_38110_17_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_17_stat_brjmp_mispredicted <= _GEN_16886;
      end
    end else begin
      T_38110_17_stat_brjmp_mispredicted <= _GEN_16886;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 404:72]
        T_38110_17_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_17_stat_btb_made_pred <= _GEN_16910;
      end
    end else begin
      T_38110_17_stat_btb_made_pred <= _GEN_16910;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 403:72]
        T_38110_17_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_17_stat_btb_mispredicted <= _GEN_16934;
      end
    end else begin
      T_38110_17_stat_btb_mispredicted <= _GEN_16934;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 406:72]
        T_38110_17_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_17_stat_bpd_made_pred <= _GEN_16958;
      end
    end else begin
      T_38110_17_stat_bpd_made_pred <= _GEN_16958;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h11 == T_28625) begin // @[rob.scala 405:72]
        T_38110_17_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_17_stat_bpd_mispredicted <= _GEN_16982;
      end
    end else begin
      T_38110_17_stat_bpd_mispredicted <= _GEN_16982;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h11 == T_28605) begin // @[rob.scala 531:53]
        T_38110_17_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_17_debug_wdata <= _GEN_24420;
      end
    end else begin
      T_38110_17_debug_wdata <= _GEN_24420;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h11 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_17_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_18_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_18_inst <= _GEN_22381;
      end
    end else begin
      T_38110_18_inst <= _GEN_22381;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43228) begin // @[rob.scala 490:10]
      T_38110_18_br_mask <= T_43230; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 402:72]
        T_38110_18_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_18_stat_brjmp_mispredicted <= _GEN_16887;
      end
    end else begin
      T_38110_18_stat_brjmp_mispredicted <= _GEN_16887;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 404:72]
        T_38110_18_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_18_stat_btb_made_pred <= _GEN_16911;
      end
    end else begin
      T_38110_18_stat_btb_made_pred <= _GEN_16911;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 403:72]
        T_38110_18_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_18_stat_btb_mispredicted <= _GEN_16935;
      end
    end else begin
      T_38110_18_stat_btb_mispredicted <= _GEN_16935;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 406:72]
        T_38110_18_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_18_stat_bpd_made_pred <= _GEN_16959;
      end
    end else begin
      T_38110_18_stat_bpd_made_pred <= _GEN_16959;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h12 == T_28625) begin // @[rob.scala 405:72]
        T_38110_18_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_18_stat_bpd_mispredicted <= _GEN_16983;
      end
    end else begin
      T_38110_18_stat_bpd_mispredicted <= _GEN_16983;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h12 == T_28605) begin // @[rob.scala 531:53]
        T_38110_18_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_18_debug_wdata <= _GEN_24421;
      end
    end else begin
      T_38110_18_debug_wdata <= _GEN_24421;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h12 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_18_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_19_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_19_inst <= _GEN_22382;
      end
    end else begin
      T_38110_19_inst <= _GEN_22382;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43330) begin // @[rob.scala 490:10]
      T_38110_19_br_mask <= T_43332; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 402:72]
        T_38110_19_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_19_stat_brjmp_mispredicted <= _GEN_16888;
      end
    end else begin
      T_38110_19_stat_brjmp_mispredicted <= _GEN_16888;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 404:72]
        T_38110_19_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_19_stat_btb_made_pred <= _GEN_16912;
      end
    end else begin
      T_38110_19_stat_btb_made_pred <= _GEN_16912;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 403:72]
        T_38110_19_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_19_stat_btb_mispredicted <= _GEN_16936;
      end
    end else begin
      T_38110_19_stat_btb_mispredicted <= _GEN_16936;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 406:72]
        T_38110_19_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_19_stat_bpd_made_pred <= _GEN_16960;
      end
    end else begin
      T_38110_19_stat_bpd_made_pred <= _GEN_16960;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h13 == T_28625) begin // @[rob.scala 405:72]
        T_38110_19_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_19_stat_bpd_mispredicted <= _GEN_16984;
      end
    end else begin
      T_38110_19_stat_bpd_mispredicted <= _GEN_16984;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h13 == T_28605) begin // @[rob.scala 531:53]
        T_38110_19_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_19_debug_wdata <= _GEN_24422;
      end
    end else begin
      T_38110_19_debug_wdata <= _GEN_24422;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h13 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_19_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_20_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_20_inst <= _GEN_22383;
      end
    end else begin
      T_38110_20_inst <= _GEN_22383;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43432) begin // @[rob.scala 490:10]
      T_38110_20_br_mask <= T_43434; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 402:72]
        T_38110_20_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_20_stat_brjmp_mispredicted <= _GEN_16889;
      end
    end else begin
      T_38110_20_stat_brjmp_mispredicted <= _GEN_16889;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 404:72]
        T_38110_20_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_20_stat_btb_made_pred <= _GEN_16913;
      end
    end else begin
      T_38110_20_stat_btb_made_pred <= _GEN_16913;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 403:72]
        T_38110_20_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_20_stat_btb_mispredicted <= _GEN_16937;
      end
    end else begin
      T_38110_20_stat_btb_mispredicted <= _GEN_16937;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 406:72]
        T_38110_20_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_20_stat_bpd_made_pred <= _GEN_16961;
      end
    end else begin
      T_38110_20_stat_bpd_made_pred <= _GEN_16961;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h14 == T_28625) begin // @[rob.scala 405:72]
        T_38110_20_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_20_stat_bpd_mispredicted <= _GEN_16985;
      end
    end else begin
      T_38110_20_stat_bpd_mispredicted <= _GEN_16985;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h14 == T_28605) begin // @[rob.scala 531:53]
        T_38110_20_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_20_debug_wdata <= _GEN_24423;
      end
    end else begin
      T_38110_20_debug_wdata <= _GEN_24423;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h14 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_20_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_21_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_21_inst <= _GEN_22384;
      end
    end else begin
      T_38110_21_inst <= _GEN_22384;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43534) begin // @[rob.scala 490:10]
      T_38110_21_br_mask <= T_43536; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 402:72]
        T_38110_21_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_21_stat_brjmp_mispredicted <= _GEN_16890;
      end
    end else begin
      T_38110_21_stat_brjmp_mispredicted <= _GEN_16890;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 404:72]
        T_38110_21_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_21_stat_btb_made_pred <= _GEN_16914;
      end
    end else begin
      T_38110_21_stat_btb_made_pred <= _GEN_16914;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 403:72]
        T_38110_21_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_21_stat_btb_mispredicted <= _GEN_16938;
      end
    end else begin
      T_38110_21_stat_btb_mispredicted <= _GEN_16938;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 406:72]
        T_38110_21_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_21_stat_bpd_made_pred <= _GEN_16962;
      end
    end else begin
      T_38110_21_stat_bpd_made_pred <= _GEN_16962;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h15 == T_28625) begin // @[rob.scala 405:72]
        T_38110_21_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_21_stat_bpd_mispredicted <= _GEN_16986;
      end
    end else begin
      T_38110_21_stat_bpd_mispredicted <= _GEN_16986;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h15 == T_28605) begin // @[rob.scala 531:53]
        T_38110_21_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_21_debug_wdata <= _GEN_24424;
      end
    end else begin
      T_38110_21_debug_wdata <= _GEN_24424;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h15 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_21_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_22_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_22_inst <= _GEN_22385;
      end
    end else begin
      T_38110_22_inst <= _GEN_22385;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43636) begin // @[rob.scala 490:10]
      T_38110_22_br_mask <= T_43638; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 402:72]
        T_38110_22_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_22_stat_brjmp_mispredicted <= _GEN_16891;
      end
    end else begin
      T_38110_22_stat_brjmp_mispredicted <= _GEN_16891;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 404:72]
        T_38110_22_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_22_stat_btb_made_pred <= _GEN_16915;
      end
    end else begin
      T_38110_22_stat_btb_made_pred <= _GEN_16915;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 403:72]
        T_38110_22_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_22_stat_btb_mispredicted <= _GEN_16939;
      end
    end else begin
      T_38110_22_stat_btb_mispredicted <= _GEN_16939;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 406:72]
        T_38110_22_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_22_stat_bpd_made_pred <= _GEN_16963;
      end
    end else begin
      T_38110_22_stat_bpd_made_pred <= _GEN_16963;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h16 == T_28625) begin // @[rob.scala 405:72]
        T_38110_22_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_22_stat_bpd_mispredicted <= _GEN_16987;
      end
    end else begin
      T_38110_22_stat_bpd_mispredicted <= _GEN_16987;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h16 == T_28605) begin // @[rob.scala 531:53]
        T_38110_22_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_22_debug_wdata <= _GEN_24425;
      end
    end else begin
      T_38110_22_debug_wdata <= _GEN_24425;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h16 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_22_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_valid <= io_dis_uops_1_valid; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_iw_state <= io_dis_uops_1_iw_state; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_uopc <= io_dis_uops_1_uopc; // @[rob.scala 350:34]
      end
    end
    if (T_44010) begin // @[rob.scala 518:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 519:33]
        T_38110_23_inst <= 32'h4033; // @[rob.scala 519:33]
      end else begin
        T_38110_23_inst <= _GEN_22386;
      end
    end else begin
      T_38110_23_inst <= _GEN_22386;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_pc <= io_dis_uops_1_pc; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_fu_code <= io_dis_uops_1_fu_code; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_br_type <= io_dis_uops_1_ctrl_br_type; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_is_load <= io_dis_uops_1_ctrl_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ctrl_is_std <= io_dis_uops_1_ctrl_is_std; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_wakeup_delay <= io_dis_uops_1_wakeup_delay; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_allocate_brtag <= io_dis_uops_1_allocate_brtag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_jump <= io_dis_uops_1_is_jump; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_jal <= io_dis_uops_1_is_jal; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_ret <= io_dis_uops_1_is_ret; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_call <= io_dis_uops_1_is_call; // @[rob.scala 350:34]
      end
    end
    if (T_43738) begin // @[rob.scala 490:10]
      T_38110_23_br_mask <= T_43740; // @[rob.scala 492:32]
    end else if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_mask <= io_dis_uops_1_br_mask; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_tag <= io_dis_uops_1_br_tag; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr; // @[rob.scala 350:34]
      end
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 402:72]
        T_38110_23_stat_brjmp_mispredicted <= io_brinfo_mispredict; // @[rob.scala 402:72]
      end else begin
        T_38110_23_stat_brjmp_mispredicted <= _GEN_16892;
      end
    end else begin
      T_38110_23_stat_brjmp_mispredicted <= _GEN_16892;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 404:72]
        T_38110_23_stat_btb_made_pred <= io_brinfo_btb_made_pred; // @[rob.scala 404:72]
      end else begin
        T_38110_23_stat_btb_made_pred <= _GEN_16916;
      end
    end else begin
      T_38110_23_stat_btb_made_pred <= _GEN_16916;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 403:72]
        T_38110_23_stat_btb_mispredicted <= io_brinfo_btb_mispredict; // @[rob.scala 403:72]
      end else begin
        T_38110_23_stat_btb_mispredicted <= _GEN_16940;
      end
    end else begin
      T_38110_23_stat_btb_mispredicted <= _GEN_16940;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 406:72]
        T_38110_23_stat_bpd_made_pred <= io_brinfo_bpd_made_pred; // @[rob.scala 406:72]
      end else begin
        T_38110_23_stat_bpd_made_pred <= _GEN_16964;
      end
    end else begin
      T_38110_23_stat_bpd_made_pred <= _GEN_16964;
    end
    if (T_40551) begin // @[rob.scala 401:7]
      if (6'h17 == T_28625) begin // @[rob.scala 405:72]
        T_38110_23_stat_bpd_mispredicted <= io_brinfo_bpd_mispredict; // @[rob.scala 405:72]
      end else begin
        T_38110_23_stat_bpd_mispredicted <= _GEN_16988;
      end
    end else begin
      T_38110_23_stat_bpd_mispredicted <= _GEN_16988;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_imm_packed <= io_dis_uops_1_imm_packed; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_csr_addr <= io_dis_uops_1_csr_addr; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_rob_idx <= io_dis_uops_1_rob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ldq_idx <= io_dis_uops_1_ldq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_stq_idx <= io_dis_uops_1_stq_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_brob_idx <= io_dis_uops_1_brob_idx; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_pdst <= io_dis_uops_1_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_pop1 <= io_dis_uops_1_pop1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_pop2 <= io_dis_uops_1_pop2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_pop3 <= io_dis_uops_1_pop3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_prs1_busy <= io_dis_uops_1_prs1_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_prs2_busy <= io_dis_uops_1_prs2_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_prs3_busy <= io_dis_uops_1_prs3_busy; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_stale_pdst <= io_dis_uops_1_stale_pdst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_exception <= io_dis_uops_1_exception; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_exc_cause <= io_dis_uops_1_exc_cause; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_bypassable <= io_dis_uops_1_bypassable; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_mem_cmd <= io_dis_uops_1_mem_cmd; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_mem_typ <= io_dis_uops_1_mem_typ; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_fence <= io_dis_uops_1_is_fence; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_fencei <= io_dis_uops_1_is_fencei; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_store <= io_dis_uops_1_is_store; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_amo <= io_dis_uops_1_is_amo; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_load <= io_dis_uops_1_is_load; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_is_unique <= io_dis_uops_1_is_unique; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_flush_on_commit <= io_dis_uops_1_flush_on_commit; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ldst <= io_dis_uops_1_ldst; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_lrs1 <= io_dis_uops_1_lrs1; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_lrs2 <= io_dis_uops_1_lrs2; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_lrs3 <= io_dis_uops_1_lrs3; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_ldst_val <= io_dis_uops_1_ldst_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_dst_rtype <= io_dis_uops_1_dst_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_lrs1_rtype <= io_dis_uops_1_lrs1_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_lrs2_rtype <= io_dis_uops_1_lrs2_rtype; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_frs3_en <= io_dis_uops_1_frs3_en; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_fp_val <= io_dis_uops_1_fp_val; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_fp_single <= io_dis_uops_1_fp_single; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_xcpt_if <= io_dis_uops_1_xcpt_if; // @[rob.scala 350:34]
      end
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_replay_if <= io_dis_uops_1_replay_if; // @[rob.scala 350:34]
      end
    end
    if (T_44507) begin // @[rob.scala 530:10]
      if (6'h17 == T_28605) begin // @[rob.scala 531:53]
        T_38110_23_debug_wdata <= io_debug_wb_wdata_2; // @[rob.scala 531:53]
      end else begin
        T_38110_23_debug_wdata <= _GEN_24426;
      end
    end else begin
      T_38110_23_debug_wdata <= _GEN_24426;
    end
    if (io_dis_valids_1) begin // @[rob.scala 346:7]
      if (5'h17 == rob_tail) begin // @[rob.scala 350:34]
        T_38110_23_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq; // @[rob.scala 350:34]
      end
    end
    T_47576 <= new_DoPrim113799324; // @[rob.scala 601:48]
    T_47616 <= new_DoPrim113799325; // @[rob.scala 608:37]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_32359) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 535:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_32359) begin
          $fatal; // @[rob.scala 535:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_32371) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 538:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_32371) begin
          $fatal; // @[rob.scala 538:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_32563) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 535:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_32563) begin
          $fatal; // @[rob.scala 535:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_32575) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 538:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_32575) begin
          $fatal; // @[rob.scala 538:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_32767) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 535:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_32767) begin
          $fatal; // @[rob.scala 535:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_32779) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 538:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_32779) begin
          $fatal; // @[rob.scala 538:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_44287) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 535:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_44287) begin
          $fatal; // @[rob.scala 535:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_44299) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 538:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_44299) begin
          $fatal; // @[rob.scala 538:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_44491) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 535:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_44491) begin
          $fatal; // @[rob.scala 535:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_44503) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 538:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_44503) begin
          $fatal; // @[rob.scala 538:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_44695) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 535:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_44695) begin
          $fatal; // @[rob.scala 535:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_44707) begin
          $fwrite(32'h80000002,
            "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n"
            ); // @[rob.scala 538:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_44707) begin
          $fatal; // @[rob.scala 538:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_47648) begin
          $fwrite(32'h80000002,
            "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:630 assert (!(io.com_valids(w) &&\n"
            ); // @[rob.scala 630:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_47648) begin
          $fatal; // @[rob.scala 630:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_47659) begin
          $fwrite(32'h80000002,
            "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:634 assert (!(io.com_valids(w) &&\n"
            ); // @[rob.scala 634:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_47659) begin
          $fatal; // @[rob.scala 634:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_47677) begin
          $fwrite(32'h80000002,
            "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:630 assert (!(io.com_valids(w) &&\n"
            ); // @[rob.scala 630:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_47677) begin
          $fatal; // @[rob.scala 630:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_47688) begin
          $fwrite(32'h80000002,
            "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:634 assert (!(io.com_valids(w) &&\n"
            ); // @[rob.scala 634:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_47688) begin
          $fatal; // @[rob.scala 634:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48105) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:693 assert (!(exception_thrown && !io.cxcpt.valid && !r_xcpt_val),\n"
            ); // @[rob.scala 693:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_48105) begin
          $fatal; // @[rob.scala 693:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48111) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:696 assert (!(io.empty && r_xcpt_val),\n"
            ); // @[rob.scala 696:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_48111) begin
          $fatal; // @[rob.scala 696:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48120) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:699 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n"
            ); // @[rob.scala 699:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_48120) begin
          $fatal; // @[rob.scala 699:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"  RobXcpt[%c%x r:%d b:%x bva:0x%x]\n",T_48223,io_debug_xcpt_uop_exc_cause,
            io_debug_xcpt_uop_rob_idx,io_debug_xcpt_uop_br_mask,io_debug_xcpt_badvaddr); // @[rob.scala 945:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h0,T_48242); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48247_data,row_metadata_has_brorjalr_T_48249_data,T_48252,T_48255,T_48258,T_48261,
            T_48262,T_48263,8'h20,T_26182_0_inst,T_38110_0_inst,T_48274,T_48277); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48292,T_26182_0_pdst,T_26182_0_br_mask,T_26182_0_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48307,T_38110_0_pdst,T_38110_0_br_mask,T_38110_0_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h1,T_48328); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48333_data,row_metadata_has_brorjalr_T_48335_data,T_48338,T_48341,T_48344,T_48347,
            T_48348,T_48349,8'h20,T_26182_1_inst,T_38110_1_inst,T_48360,T_48363); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48378,T_26182_1_pdst,T_26182_1_br_mask,T_26182_1_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48393,T_38110_1_pdst,T_38110_1_br_mask,T_38110_1_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h2,T_48414); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48419_data,row_metadata_has_brorjalr_T_48421_data,T_48424,T_48427,T_48430,T_48433,
            T_48434,T_48435,8'h20,T_26182_2_inst,T_38110_2_inst,T_48446,T_48449); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48464,T_26182_2_pdst,T_26182_2_br_mask,T_26182_2_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48479,T_38110_2_pdst,T_38110_2_br_mask,T_38110_2_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h3,T_48500); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48505_data,row_metadata_has_brorjalr_T_48507_data,T_48510,T_48513,T_48516,T_48519,
            T_48520,T_48521,8'h20,T_26182_3_inst,T_38110_3_inst,T_48532,T_48535); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48550,T_26182_3_pdst,T_26182_3_br_mask,T_26182_3_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48565,T_38110_3_pdst,T_38110_3_br_mask,T_38110_3_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h4,T_48586); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48591_data,row_metadata_has_brorjalr_T_48593_data,T_48596,T_48599,T_48602,T_48605,
            T_48606,T_48607,8'h20,T_26182_4_inst,T_38110_4_inst,T_48618,T_48621); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48636,T_26182_4_pdst,T_26182_4_br_mask,T_26182_4_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48651,T_38110_4_pdst,T_38110_4_br_mask,T_38110_4_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h5,T_48672); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48677_data,row_metadata_has_brorjalr_T_48679_data,T_48682,T_48685,T_48688,T_48691,
            T_48692,T_48693,8'h20,T_26182_5_inst,T_38110_5_inst,T_48704,T_48707); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48722,T_26182_5_pdst,T_26182_5_br_mask,T_26182_5_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48737,T_38110_5_pdst,T_38110_5_br_mask,T_38110_5_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h6,T_48758); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48763_data,row_metadata_has_brorjalr_T_48765_data,T_48768,T_48771,T_48774,T_48777,
            T_48778,T_48779,8'h20,T_26182_6_inst,T_38110_6_inst,T_48790,T_48793); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48808,T_26182_6_pdst,T_26182_6_br_mask,T_26182_6_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48823,T_38110_6_pdst,T_38110_6_br_mask,T_38110_6_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h7,T_48844); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48849_data,row_metadata_has_brorjalr_T_48851_data,T_48854,T_48857,T_48860,T_48863,
            T_48864,T_48865,8'h20,T_26182_7_inst,T_38110_7_inst,T_48876,T_48879); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48894,T_26182_7_pdst,T_26182_7_br_mask,T_26182_7_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48909,T_38110_7_pdst,T_38110_7_br_mask,T_38110_7_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h8,T_48930); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_48935_data,row_metadata_has_brorjalr_T_48937_data,T_48940,T_48943,T_48946,T_48949,
            T_48950,T_48951,8'h20,T_26182_8_inst,T_38110_8_inst,T_48962,T_48965); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48980,T_26182_8_pdst,T_26182_8_br_mask,T_26182_8_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_48995,T_38110_8_pdst,T_38110_8_br_mask,T_38110_8_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h9,T_49016); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49021_data,row_metadata_has_brorjalr_T_49023_data,T_49026,T_49029,T_49032,T_49035,
            T_49036,T_49037,8'h20,T_26182_9_inst,T_38110_9_inst,T_49048,T_49051); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49066,T_26182_9_pdst,T_26182_9_br_mask,T_26182_9_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49081,T_38110_9_pdst,T_38110_9_br_mask,T_38110_9_stale_pdst
            ); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'ha,T_49102); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49107_data,row_metadata_has_brorjalr_T_49109_data,T_49112,T_49115,T_49118,T_49121,
            T_49122,T_49123,8'h20,T_26182_10_inst,T_38110_10_inst,T_49134,T_49137); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49152,T_26182_10_pdst,T_26182_10_br_mask,
            T_26182_10_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49167,T_38110_10_pdst,T_38110_10_br_mask,
            T_38110_10_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'hb,T_49188); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49193_data,row_metadata_has_brorjalr_T_49195_data,T_49198,T_49201,T_49204,T_49207,
            T_49208,T_49209,8'h20,T_26182_11_inst,T_38110_11_inst,T_49220,T_49223); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49238,T_26182_11_pdst,T_26182_11_br_mask,
            T_26182_11_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49253,T_38110_11_pdst,T_38110_11_br_mask,
            T_38110_11_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'hc,T_49274); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49279_data,row_metadata_has_brorjalr_T_49281_data,T_49284,T_49287,T_49290,T_49293,
            T_49294,T_49295,8'h20,T_26182_12_inst,T_38110_12_inst,T_49306,T_49309); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49324,T_26182_12_pdst,T_26182_12_br_mask,
            T_26182_12_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49339,T_38110_12_pdst,T_38110_12_br_mask,
            T_38110_12_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'hd,T_49360); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49365_data,row_metadata_has_brorjalr_T_49367_data,T_49370,T_49373,T_49376,T_49379,
            T_49380,T_49381,8'h20,T_26182_13_inst,T_38110_13_inst,T_49392,T_49395); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49410,T_26182_13_pdst,T_26182_13_br_mask,
            T_26182_13_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49425,T_38110_13_pdst,T_38110_13_br_mask,
            T_38110_13_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'he,T_49446); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49451_data,row_metadata_has_brorjalr_T_49453_data,T_49456,T_49459,T_49462,T_49465,
            T_49466,T_49467,8'h20,T_26182_14_inst,T_38110_14_inst,T_49478,T_49481); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49496,T_26182_14_pdst,T_26182_14_br_mask,
            T_26182_14_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49511,T_38110_14_pdst,T_38110_14_br_mask,
            T_38110_14_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'hf,T_49532); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49537_data,row_metadata_has_brorjalr_T_49539_data,T_49542,T_49545,T_49548,T_49551,
            T_49552,T_49553,8'h20,T_26182_15_inst,T_38110_15_inst,T_49564,T_49567); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49582,T_26182_15_pdst,T_26182_15_br_mask,
            T_26182_15_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49597,T_38110_15_pdst,T_38110_15_br_mask,
            T_38110_15_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h10,T_49618); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49623_data,row_metadata_has_brorjalr_T_49625_data,T_49628,T_49631,T_49634,T_49637,
            T_49638,T_49639,8'h20,T_26182_16_inst,T_38110_16_inst,T_49650,T_49653); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49668,T_26182_16_pdst,T_26182_16_br_mask,
            T_26182_16_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49683,T_38110_16_pdst,T_38110_16_br_mask,
            T_38110_16_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h11,T_49704); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49709_data,row_metadata_has_brorjalr_T_49711_data,T_49714,T_49717,T_49720,T_49723,
            T_49724,T_49725,8'h20,T_26182_17_inst,T_38110_17_inst,T_49736,T_49739); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49754,T_26182_17_pdst,T_26182_17_br_mask,
            T_26182_17_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49769,T_38110_17_pdst,T_38110_17_br_mask,
            T_38110_17_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h12,T_49790); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49795_data,row_metadata_has_brorjalr_T_49797_data,T_49800,T_49803,T_49806,T_49809,
            T_49810,T_49811,8'h20,T_26182_18_inst,T_38110_18_inst,T_49822,T_49825); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49840,T_26182_18_pdst,T_26182_18_br_mask,
            T_26182_18_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49855,T_38110_18_pdst,T_38110_18_br_mask,
            T_38110_18_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h13,T_49876); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49881_data,row_metadata_has_brorjalr_T_49883_data,T_49886,T_49889,T_49892,T_49895,
            T_49896,T_49897,8'h20,T_26182_19_inst,T_38110_19_inst,T_49908,T_49911); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49926,T_26182_19_pdst,T_26182_19_br_mask,
            T_26182_19_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_49941,T_38110_19_pdst,T_38110_19_br_mask,
            T_38110_19_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h14,T_49962); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_49967_data,row_metadata_has_brorjalr_T_49969_data,T_49972,T_49975,T_49978,T_49981,
            T_49982,T_49983,8'h20,T_26182_20_inst,T_38110_20_inst,T_49994,T_49997); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50012,T_26182_20_pdst,T_26182_20_br_mask,
            T_26182_20_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50027,T_38110_20_pdst,T_38110_20_br_mask,
            T_38110_20_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h15,T_50048); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_50053_data,row_metadata_has_brorjalr_T_50055_data,T_50058,T_50061,T_50064,T_50067,
            T_50068,T_50069,8'h20,T_26182_21_inst,T_38110_21_inst,T_50080,T_50083); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50098,T_26182_21_pdst,T_26182_21_br_mask,
            T_26182_21_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50113,T_38110_21_pdst,T_38110_21_br_mask,
            T_38110_21_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h16,T_50134); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_50139_data,row_metadata_has_brorjalr_T_50141_data,T_50144,T_50147,T_50150,T_50153,
            T_50154,T_50155,8'h20,T_26182_22_inst,T_38110_22_inst,T_50166,T_50169); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50184,T_26182_22_pdst,T_26182_22_br_mask,
            T_26182_22_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50199,T_38110_22_pdst,T_38110_22_br_mask,
            T_38110_22_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"    rob[%d] %c (",6'h17,T_50220); // @[rob.scala 967:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ",
            row_metadata_brob_idx_T_50225_data,row_metadata_has_brorjalr_T_50227_data,T_50230,T_50233,T_50236,T_50239,
            T_50240,T_50241,8'h20,T_26182_23_inst,T_38110_23_inst,T_50252,T_50255); // @[rob.scala 993:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50270,T_26182_23_pdst,T_26182_23_br_mask,
            T_26182_23_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"(d:%c p%d, bm:%x sdt:%d) ",T_50285,T_38110_23_pdst,T_38110_23_br_mask,
            T_38110_23_stale_pdst); // @[rob.scala 1047:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_48225) begin
          $fwrite(32'h80000002,"\n"); // @[rob.scala 1061:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  _RAND_3 = {2{`RANDOM}};
  _RAND_4 = {2{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_6 = {2{`RANDOM}};
  _RAND_7 = {2{`RANDOM}};
  _RAND_8 = {2{`RANDOM}};
  _RAND_9 = {2{`RANDOM}};
  _RAND_10 = {2{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
  _RAND_12 = {2{`RANDOM}};
  _RAND_13 = {2{`RANDOM}};
  _RAND_14 = {2{`RANDOM}};
  _RAND_15 = {2{`RANDOM}};
  _RAND_16 = {2{`RANDOM}};
  _RAND_17 = {2{`RANDOM}};
  _RAND_18 = {2{`RANDOM}};
  _RAND_19 = {2{`RANDOM}};
  _RAND_20 = {2{`RANDOM}};
  _RAND_21 = {2{`RANDOM}};
  _RAND_22 = {2{`RANDOM}};
  _RAND_23 = {2{`RANDOM}};
  _RAND_24 = {2{`RANDOM}};
  _RAND_25 = {2{`RANDOM}};
  _RAND_26 = {2{`RANDOM}};
  _RAND_27 = {2{`RANDOM}};
  _RAND_28 = {2{`RANDOM}};
  _RAND_29 = {2{`RANDOM}};
  _RAND_30 = {2{`RANDOM}};
  _RAND_31 = {2{`RANDOM}};
  _RAND_32 = {2{`RANDOM}};
  _RAND_33 = {2{`RANDOM}};
  _RAND_34 = {2{`RANDOM}};
  _RAND_35 = {2{`RANDOM}};
  _RAND_36 = {2{`RANDOM}};
  _RAND_37 = {2{`RANDOM}};
  _RAND_38 = {2{`RANDOM}};
  _RAND_39 = {2{`RANDOM}};
  _RAND_40 = {2{`RANDOM}};
  _RAND_41 = {2{`RANDOM}};
  _RAND_42 = {2{`RANDOM}};
  _RAND_43 = {2{`RANDOM}};
  _RAND_44 = {2{`RANDOM}};
  _RAND_45 = {2{`RANDOM}};
  _RAND_46 = {2{`RANDOM}};
  _RAND_47 = {2{`RANDOM}};
  _RAND_48 = {2{`RANDOM}};
  _RAND_49 = {2{`RANDOM}};
  _RAND_50 = {2{`RANDOM}};
  _RAND_52 = {2{`RANDOM}};
  _RAND_53 = {2{`RANDOM}};
  _RAND_54 = {2{`RANDOM}};
  _RAND_55 = {2{`RANDOM}};
  _RAND_56 = {2{`RANDOM}};
  _RAND_57 = {2{`RANDOM}};
  _RAND_58 = {2{`RANDOM}};
  _RAND_59 = {2{`RANDOM}};
  _RAND_60 = {2{`RANDOM}};
  _RAND_61 = {2{`RANDOM}};
  _RAND_62 = {2{`RANDOM}};
  _RAND_63 = {2{`RANDOM}};
  _RAND_64 = {2{`RANDOM}};
  _RAND_65 = {2{`RANDOM}};
  _RAND_66 = {2{`RANDOM}};
  _RAND_67 = {2{`RANDOM}};
  _RAND_68 = {2{`RANDOM}};
  _RAND_69 = {2{`RANDOM}};
  _RAND_70 = {2{`RANDOM}};
  _RAND_71 = {2{`RANDOM}};
  _RAND_72 = {2{`RANDOM}};
  _RAND_73 = {2{`RANDOM}};
  _RAND_74 = {2{`RANDOM}};
  _RAND_75 = {2{`RANDOM}};
  _RAND_76 = {2{`RANDOM}};
  _RAND_77 = {2{`RANDOM}};
  _RAND_78 = {2{`RANDOM}};
  _RAND_79 = {2{`RANDOM}};
  _RAND_80 = {2{`RANDOM}};
  _RAND_81 = {2{`RANDOM}};
  _RAND_82 = {2{`RANDOM}};
  _RAND_83 = {2{`RANDOM}};
  _RAND_84 = {2{`RANDOM}};
  _RAND_85 = {2{`RANDOM}};
  _RAND_86 = {2{`RANDOM}};
  _RAND_87 = {2{`RANDOM}};
  _RAND_88 = {2{`RANDOM}};
  _RAND_89 = {2{`RANDOM}};
  _RAND_90 = {2{`RANDOM}};
  _RAND_91 = {2{`RANDOM}};
  _RAND_92 = {2{`RANDOM}};
  _RAND_93 = {2{`RANDOM}};
  _RAND_94 = {2{`RANDOM}};
  _RAND_95 = {2{`RANDOM}};
  _RAND_96 = {2{`RANDOM}};
  _RAND_97 = {2{`RANDOM}};
  _RAND_98 = {2{`RANDOM}};
  _RAND_99 = {2{`RANDOM}};
  _RAND_100 = {2{`RANDOM}};
  _RAND_101 = {2{`RANDOM}};
  _RAND_103 = {1{`RANDOM}};
  _RAND_104 = {1{`RANDOM}};
  _RAND_105 = {1{`RANDOM}};
  _RAND_106 = {1{`RANDOM}};
  _RAND_107 = {1{`RANDOM}};
  _RAND_108 = {1{`RANDOM}};
  _RAND_109 = {1{`RANDOM}};
  _RAND_110 = {1{`RANDOM}};
  _RAND_111 = {1{`RANDOM}};
  _RAND_112 = {1{`RANDOM}};
  _RAND_113 = {1{`RANDOM}};
  _RAND_114 = {1{`RANDOM}};
  _RAND_115 = {1{`RANDOM}};
  _RAND_116 = {1{`RANDOM}};
  _RAND_117 = {1{`RANDOM}};
  _RAND_118 = {1{`RANDOM}};
  _RAND_119 = {1{`RANDOM}};
  _RAND_120 = {1{`RANDOM}};
  _RAND_121 = {1{`RANDOM}};
  _RAND_122 = {1{`RANDOM}};
  _RAND_123 = {1{`RANDOM}};
  _RAND_124 = {1{`RANDOM}};
  _RAND_125 = {1{`RANDOM}};
  _RAND_126 = {1{`RANDOM}};
  _RAND_127 = {1{`RANDOM}};
  _RAND_128 = {1{`RANDOM}};
  _RAND_130 = {1{`RANDOM}};
  _RAND_131 = {1{`RANDOM}};
  _RAND_132 = {1{`RANDOM}};
  _RAND_133 = {1{`RANDOM}};
  _RAND_134 = {1{`RANDOM}};
  _RAND_135 = {1{`RANDOM}};
  _RAND_136 = {1{`RANDOM}};
  _RAND_137 = {1{`RANDOM}};
  _RAND_138 = {1{`RANDOM}};
  _RAND_139 = {1{`RANDOM}};
  _RAND_140 = {1{`RANDOM}};
  _RAND_141 = {1{`RANDOM}};
  _RAND_142 = {1{`RANDOM}};
  _RAND_143 = {1{`RANDOM}};
  _RAND_144 = {1{`RANDOM}};
  _RAND_145 = {1{`RANDOM}};
  _RAND_146 = {1{`RANDOM}};
  _RAND_147 = {1{`RANDOM}};
  _RAND_148 = {1{`RANDOM}};
  _RAND_149 = {1{`RANDOM}};
  _RAND_150 = {1{`RANDOM}};
  _RAND_151 = {1{`RANDOM}};
  _RAND_152 = {1{`RANDOM}};
  _RAND_153 = {1{`RANDOM}};
  _RAND_154 = {1{`RANDOM}};
  _RAND_156 = {1{`RANDOM}};
  _RAND_157 = {1{`RANDOM}};
  _RAND_158 = {1{`RANDOM}};
  _RAND_159 = {1{`RANDOM}};
  _RAND_160 = {1{`RANDOM}};
  _RAND_161 = {1{`RANDOM}};
  _RAND_162 = {1{`RANDOM}};
  _RAND_163 = {1{`RANDOM}};
  _RAND_164 = {1{`RANDOM}};
  _RAND_165 = {1{`RANDOM}};
  _RAND_166 = {1{`RANDOM}};
  _RAND_167 = {1{`RANDOM}};
  _RAND_168 = {1{`RANDOM}};
  _RAND_169 = {1{`RANDOM}};
  _RAND_170 = {1{`RANDOM}};
  _RAND_171 = {1{`RANDOM}};
  _RAND_172 = {1{`RANDOM}};
  _RAND_173 = {1{`RANDOM}};
  _RAND_174 = {1{`RANDOM}};
  _RAND_175 = {1{`RANDOM}};
  _RAND_176 = {1{`RANDOM}};
  _RAND_177 = {1{`RANDOM}};
  _RAND_178 = {1{`RANDOM}};
  _RAND_179 = {1{`RANDOM}};
  _RAND_180 = {1{`RANDOM}};
  _RAND_182 = {1{`RANDOM}};
  _RAND_183 = {1{`RANDOM}};
  _RAND_184 = {1{`RANDOM}};
  _RAND_185 = {1{`RANDOM}};
  _RAND_186 = {1{`RANDOM}};
  _RAND_187 = {1{`RANDOM}};
  _RAND_188 = {1{`RANDOM}};
  _RAND_189 = {1{`RANDOM}};
  _RAND_190 = {1{`RANDOM}};
  _RAND_191 = {1{`RANDOM}};
  _RAND_192 = {1{`RANDOM}};
  _RAND_193 = {1{`RANDOM}};
  _RAND_194 = {1{`RANDOM}};
  _RAND_195 = {1{`RANDOM}};
  _RAND_196 = {1{`RANDOM}};
  _RAND_197 = {1{`RANDOM}};
  _RAND_198 = {1{`RANDOM}};
  _RAND_199 = {1{`RANDOM}};
  _RAND_200 = {1{`RANDOM}};
  _RAND_201 = {1{`RANDOM}};
  _RAND_202 = {1{`RANDOM}};
  _RAND_203 = {1{`RANDOM}};
  _RAND_204 = {1{`RANDOM}};
  _RAND_205 = {1{`RANDOM}};
  _RAND_206 = {1{`RANDOM}};
  _RAND_208 = {1{`RANDOM}};
  _RAND_210 = {1{`RANDOM}};
  _RAND_211 = {1{`RANDOM}};
  _RAND_212 = {1{`RANDOM}};
  _RAND_213 = {1{`RANDOM}};
  _RAND_214 = {1{`RANDOM}};
  _RAND_215 = {1{`RANDOM}};
  _RAND_216 = {1{`RANDOM}};
  _RAND_217 = {1{`RANDOM}};
  _RAND_218 = {1{`RANDOM}};
  _RAND_219 = {1{`RANDOM}};
  _RAND_220 = {1{`RANDOM}};
  _RAND_221 = {1{`RANDOM}};
  _RAND_222 = {1{`RANDOM}};
  _RAND_223 = {1{`RANDOM}};
  _RAND_224 = {1{`RANDOM}};
  _RAND_225 = {1{`RANDOM}};
  _RAND_226 = {1{`RANDOM}};
  _RAND_227 = {1{`RANDOM}};
  _RAND_228 = {1{`RANDOM}};
  _RAND_229 = {1{`RANDOM}};
  _RAND_230 = {1{`RANDOM}};
  _RAND_231 = {1{`RANDOM}};
  _RAND_232 = {1{`RANDOM}};
  _RAND_233 = {1{`RANDOM}};
  _RAND_234 = {1{`RANDOM}};
  _RAND_236 = {1{`RANDOM}};
  _RAND_237 = {1{`RANDOM}};
  _RAND_238 = {1{`RANDOM}};
  _RAND_239 = {1{`RANDOM}};
  _RAND_240 = {1{`RANDOM}};
  _RAND_241 = {1{`RANDOM}};
  _RAND_242 = {1{`RANDOM}};
  _RAND_243 = {1{`RANDOM}};
  _RAND_244 = {1{`RANDOM}};
  _RAND_245 = {1{`RANDOM}};
  _RAND_246 = {1{`RANDOM}};
  _RAND_247 = {1{`RANDOM}};
  _RAND_248 = {1{`RANDOM}};
  _RAND_249 = {1{`RANDOM}};
  _RAND_250 = {1{`RANDOM}};
  _RAND_251 = {1{`RANDOM}};
  _RAND_252 = {1{`RANDOM}};
  _RAND_253 = {1{`RANDOM}};
  _RAND_254 = {1{`RANDOM}};
  _RAND_255 = {1{`RANDOM}};
  _RAND_256 = {1{`RANDOM}};
  _RAND_257 = {1{`RANDOM}};
  _RAND_258 = {1{`RANDOM}};
  _RAND_259 = {1{`RANDOM}};
  _RAND_260 = {1{`RANDOM}};
  _RAND_262 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    T_23555[initvar] = _RAND_0[36:0];
  _RAND_51 = {2{`RANDOM}};
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    T_23558[initvar] = _RAND_51[36:0];
  _RAND_102 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    row_metadata_brob_idx[initvar] = _RAND_102[4:0];
  _RAND_129 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    row_metadata_has_brorjalr[initvar] = _RAND_129[0:0];
  _RAND_155 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    T_23710[initvar] = _RAND_155[0:0];
  _RAND_181 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    T_28311[initvar] = _RAND_181[0:0];
  _RAND_207 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    T_28314[initvar] = _RAND_207[4:0];
  _RAND_209 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    T_35638[initvar] = _RAND_209[0:0];
  _RAND_235 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    T_40239[initvar] = _RAND_235[0:0];
  _RAND_261 = {1{`RANDOM}};
  for (initvar = 0; initvar < 24; initvar = initvar+1)
    T_40242[initvar] = _RAND_261[4:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  rob_state = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  rob_head = _RAND_264[4:0];
  _RAND_265 = {1{`RANDOM}};
  rob_tail = _RAND_265[4:0];
  _RAND_266 = {1{`RANDOM}};
  r_xcpt_val = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_xcpt_uop_valid = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_xcpt_uop_iw_state = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  r_xcpt_uop_uopc = _RAND_269[8:0];
  _RAND_270 = {1{`RANDOM}};
  r_xcpt_uop_inst = _RAND_270[31:0];
  _RAND_271 = {2{`RANDOM}};
  r_xcpt_uop_pc = _RAND_271[39:0];
  _RAND_272 = {1{`RANDOM}};
  r_xcpt_uop_fu_code = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_br_type = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_op1_sel = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_op2_sel = _RAND_275[2:0];
  _RAND_276 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_imm_sel = _RAND_276[2:0];
  _RAND_277 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_op_fcn = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_fcn_dw = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_rf_wen = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_csr_cmd = _RAND_280[2:0];
  _RAND_281 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_is_load = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_is_sta = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_xcpt_uop_ctrl_is_std = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_xcpt_uop_wakeup_delay = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  r_xcpt_uop_allocate_brtag = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_xcpt_uop_is_br_or_jmp = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_xcpt_uop_is_jump = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_xcpt_uop_is_jal = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_xcpt_uop_is_ret = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_xcpt_uop_is_call = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_xcpt_uop_br_mask = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  r_xcpt_uop_br_tag = _RAND_292[2:0];
  _RAND_293 = {1{`RANDOM}};
  r_xcpt_uop_br_prediction_bpd_predict_val = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_xcpt_uop_br_prediction_bpd_predict_taken = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_xcpt_uop_br_prediction_btb_hit = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_xcpt_uop_br_prediction_btb_predicted = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_xcpt_uop_br_prediction_is_br_or_jalr = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_xcpt_uop_stat_brjmp_mispredicted = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_xcpt_uop_stat_btb_made_pred = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_xcpt_uop_stat_btb_mispredicted = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_xcpt_uop_stat_bpd_made_pred = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_xcpt_uop_stat_bpd_mispredicted = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_xcpt_uop_fetch_pc_lob = _RAND_303[2:0];
  _RAND_304 = {1{`RANDOM}};
  r_xcpt_uop_imm_packed = _RAND_304[19:0];
  _RAND_305 = {1{`RANDOM}};
  r_xcpt_uop_csr_addr = _RAND_305[11:0];
  _RAND_306 = {1{`RANDOM}};
  r_xcpt_uop_rob_idx = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  r_xcpt_uop_ldq_idx = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  r_xcpt_uop_stq_idx = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  r_xcpt_uop_brob_idx = _RAND_309[4:0];
  _RAND_310 = {1{`RANDOM}};
  r_xcpt_uop_pdst = _RAND_310[6:0];
  _RAND_311 = {1{`RANDOM}};
  r_xcpt_uop_pop1 = _RAND_311[6:0];
  _RAND_312 = {1{`RANDOM}};
  r_xcpt_uop_pop2 = _RAND_312[6:0];
  _RAND_313 = {1{`RANDOM}};
  r_xcpt_uop_pop3 = _RAND_313[6:0];
  _RAND_314 = {1{`RANDOM}};
  r_xcpt_uop_prs1_busy = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_xcpt_uop_prs2_busy = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_xcpt_uop_prs3_busy = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_xcpt_uop_stale_pdst = _RAND_317[6:0];
  _RAND_318 = {1{`RANDOM}};
  r_xcpt_uop_exception = _RAND_318[0:0];
  _RAND_319 = {2{`RANDOM}};
  r_xcpt_uop_exc_cause = _RAND_319[63:0];
  _RAND_320 = {1{`RANDOM}};
  r_xcpt_uop_bypassable = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_xcpt_uop_mem_cmd = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  r_xcpt_uop_mem_typ = _RAND_322[2:0];
  _RAND_323 = {1{`RANDOM}};
  r_xcpt_uop_is_fence = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_xcpt_uop_is_fencei = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_xcpt_uop_is_store = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_xcpt_uop_is_amo = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_xcpt_uop_is_load = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_xcpt_uop_is_unique = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_xcpt_uop_flush_on_commit = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_xcpt_uop_ldst = _RAND_330[5:0];
  _RAND_331 = {1{`RANDOM}};
  r_xcpt_uop_lrs1 = _RAND_331[5:0];
  _RAND_332 = {1{`RANDOM}};
  r_xcpt_uop_lrs2 = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  r_xcpt_uop_lrs3 = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  r_xcpt_uop_ldst_val = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_xcpt_uop_dst_rtype = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  r_xcpt_uop_lrs1_rtype = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  r_xcpt_uop_lrs2_rtype = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  r_xcpt_uop_frs3_en = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_xcpt_uop_fp_val = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_xcpt_uop_fp_single = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_xcpt_uop_xcpt_if = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_xcpt_uop_replay_if = _RAND_342[0:0];
  _RAND_343 = {2{`RANDOM}};
  r_xcpt_uop_debug_wdata = _RAND_343[63:0];
  _RAND_344 = {1{`RANDOM}};
  r_xcpt_uop_debug_events_fetch_seq = _RAND_344[31:0];
  _RAND_345 = {2{`RANDOM}};
  r_xcpt_badvaddr = _RAND_345[39:0];
  _RAND_346 = {1{`RANDOM}};
  T_35634_23 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  T_35634_22 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  T_35634_21 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  T_35634_20 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  T_35634_19 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  T_35634_18 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  T_35634_17 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  T_35634_16 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  T_35634_15 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  T_35634_14 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  T_35634_13 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  T_35634_12 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  T_35634_11 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  T_35634_10 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  T_35634_9 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  T_35634_8 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  T_35634_7 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  T_35634_6 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  T_35634_5 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  T_35634_4 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  T_35634_3 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  T_35634_2 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  T_35634_1 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  T_35634_0 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  T_23706_23 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  T_23706_22 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  T_23706_21 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  T_23706_20 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  T_23706_19 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  T_23706_18 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  T_23706_17 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  T_23706_16 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  T_23706_15 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  T_23706_14 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  T_23706_13 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  T_23706_12 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  T_23706_11 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  T_23706_10 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  T_23706_9 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  T_23706_8 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  T_23706_7 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  T_23706_6 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  T_23706_5 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  T_23706_4 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  T_23706_3 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  T_23706_2 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  T_23706_1 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  T_23706_0 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_partial_row = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  T_26182_0_valid = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  T_26182_0_iw_state = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  T_26182_0_uopc = _RAND_397[8:0];
  _RAND_398 = {1{`RANDOM}};
  T_26182_0_inst = _RAND_398[31:0];
  _RAND_399 = {2{`RANDOM}};
  T_26182_0_pc = _RAND_399[39:0];
  _RAND_400 = {1{`RANDOM}};
  T_26182_0_fu_code = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  T_26182_0_ctrl_br_type = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  T_26182_0_ctrl_op1_sel = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  T_26182_0_ctrl_op2_sel = _RAND_403[2:0];
  _RAND_404 = {1{`RANDOM}};
  T_26182_0_ctrl_imm_sel = _RAND_404[2:0];
  _RAND_405 = {1{`RANDOM}};
  T_26182_0_ctrl_op_fcn = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  T_26182_0_ctrl_fcn_dw = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  T_26182_0_ctrl_rf_wen = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  T_26182_0_ctrl_csr_cmd = _RAND_408[2:0];
  _RAND_409 = {1{`RANDOM}};
  T_26182_0_ctrl_is_load = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  T_26182_0_ctrl_is_sta = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  T_26182_0_ctrl_is_std = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  T_26182_0_wakeup_delay = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  T_26182_0_allocate_brtag = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  T_26182_0_is_br_or_jmp = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  T_26182_0_is_jump = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  T_26182_0_is_jal = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  T_26182_0_is_ret = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  T_26182_0_is_call = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  T_26182_0_br_mask = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  T_26182_0_br_tag = _RAND_420[2:0];
  _RAND_421 = {1{`RANDOM}};
  T_26182_0_br_prediction_bpd_predict_val = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  T_26182_0_br_prediction_bpd_predict_taken = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  T_26182_0_br_prediction_btb_hit = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  T_26182_0_br_prediction_btb_predicted = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  T_26182_0_br_prediction_is_br_or_jalr = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  T_26182_0_stat_brjmp_mispredicted = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  T_26182_0_stat_btb_made_pred = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  T_26182_0_stat_btb_mispredicted = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  T_26182_0_stat_bpd_made_pred = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  T_26182_0_stat_bpd_mispredicted = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  T_26182_0_fetch_pc_lob = _RAND_431[2:0];
  _RAND_432 = {1{`RANDOM}};
  T_26182_0_imm_packed = _RAND_432[19:0];
  _RAND_433 = {1{`RANDOM}};
  T_26182_0_csr_addr = _RAND_433[11:0];
  _RAND_434 = {1{`RANDOM}};
  T_26182_0_rob_idx = _RAND_434[5:0];
  _RAND_435 = {1{`RANDOM}};
  T_26182_0_ldq_idx = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  T_26182_0_stq_idx = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  T_26182_0_brob_idx = _RAND_437[4:0];
  _RAND_438 = {1{`RANDOM}};
  T_26182_0_pdst = _RAND_438[6:0];
  _RAND_439 = {1{`RANDOM}};
  T_26182_0_pop1 = _RAND_439[6:0];
  _RAND_440 = {1{`RANDOM}};
  T_26182_0_pop2 = _RAND_440[6:0];
  _RAND_441 = {1{`RANDOM}};
  T_26182_0_pop3 = _RAND_441[6:0];
  _RAND_442 = {1{`RANDOM}};
  T_26182_0_prs1_busy = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  T_26182_0_prs2_busy = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  T_26182_0_prs3_busy = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  T_26182_0_stale_pdst = _RAND_445[6:0];
  _RAND_446 = {1{`RANDOM}};
  T_26182_0_exception = _RAND_446[0:0];
  _RAND_447 = {2{`RANDOM}};
  T_26182_0_exc_cause = _RAND_447[63:0];
  _RAND_448 = {1{`RANDOM}};
  T_26182_0_bypassable = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  T_26182_0_mem_cmd = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  T_26182_0_mem_typ = _RAND_450[2:0];
  _RAND_451 = {1{`RANDOM}};
  T_26182_0_is_fence = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  T_26182_0_is_fencei = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  T_26182_0_is_store = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  T_26182_0_is_amo = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  T_26182_0_is_load = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  T_26182_0_is_unique = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  T_26182_0_flush_on_commit = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  T_26182_0_ldst = _RAND_458[5:0];
  _RAND_459 = {1{`RANDOM}};
  T_26182_0_lrs1 = _RAND_459[5:0];
  _RAND_460 = {1{`RANDOM}};
  T_26182_0_lrs2 = _RAND_460[5:0];
  _RAND_461 = {1{`RANDOM}};
  T_26182_0_lrs3 = _RAND_461[5:0];
  _RAND_462 = {1{`RANDOM}};
  T_26182_0_ldst_val = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  T_26182_0_dst_rtype = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  T_26182_0_lrs1_rtype = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  T_26182_0_lrs2_rtype = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  T_26182_0_frs3_en = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  T_26182_0_fp_val = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  T_26182_0_fp_single = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  T_26182_0_xcpt_if = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  T_26182_0_replay_if = _RAND_470[0:0];
  _RAND_471 = {2{`RANDOM}};
  T_26182_0_debug_wdata = _RAND_471[63:0];
  _RAND_472 = {1{`RANDOM}};
  T_26182_0_debug_events_fetch_seq = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  T_26182_1_valid = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  T_26182_1_iw_state = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  T_26182_1_uopc = _RAND_475[8:0];
  _RAND_476 = {1{`RANDOM}};
  T_26182_1_inst = _RAND_476[31:0];
  _RAND_477 = {2{`RANDOM}};
  T_26182_1_pc = _RAND_477[39:0];
  _RAND_478 = {1{`RANDOM}};
  T_26182_1_fu_code = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  T_26182_1_ctrl_br_type = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  T_26182_1_ctrl_op1_sel = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  T_26182_1_ctrl_op2_sel = _RAND_481[2:0];
  _RAND_482 = {1{`RANDOM}};
  T_26182_1_ctrl_imm_sel = _RAND_482[2:0];
  _RAND_483 = {1{`RANDOM}};
  T_26182_1_ctrl_op_fcn = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  T_26182_1_ctrl_fcn_dw = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  T_26182_1_ctrl_rf_wen = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  T_26182_1_ctrl_csr_cmd = _RAND_486[2:0];
  _RAND_487 = {1{`RANDOM}};
  T_26182_1_ctrl_is_load = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  T_26182_1_ctrl_is_sta = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  T_26182_1_ctrl_is_std = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  T_26182_1_wakeup_delay = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  T_26182_1_allocate_brtag = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  T_26182_1_is_br_or_jmp = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  T_26182_1_is_jump = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  T_26182_1_is_jal = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  T_26182_1_is_ret = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  T_26182_1_is_call = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  T_26182_1_br_mask = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  T_26182_1_br_tag = _RAND_498[2:0];
  _RAND_499 = {1{`RANDOM}};
  T_26182_1_br_prediction_bpd_predict_val = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  T_26182_1_br_prediction_bpd_predict_taken = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  T_26182_1_br_prediction_btb_hit = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  T_26182_1_br_prediction_btb_predicted = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  T_26182_1_br_prediction_is_br_or_jalr = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  T_26182_1_stat_brjmp_mispredicted = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  T_26182_1_stat_btb_made_pred = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  T_26182_1_stat_btb_mispredicted = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  T_26182_1_stat_bpd_made_pred = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  T_26182_1_stat_bpd_mispredicted = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  T_26182_1_fetch_pc_lob = _RAND_509[2:0];
  _RAND_510 = {1{`RANDOM}};
  T_26182_1_imm_packed = _RAND_510[19:0];
  _RAND_511 = {1{`RANDOM}};
  T_26182_1_csr_addr = _RAND_511[11:0];
  _RAND_512 = {1{`RANDOM}};
  T_26182_1_rob_idx = _RAND_512[5:0];
  _RAND_513 = {1{`RANDOM}};
  T_26182_1_ldq_idx = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  T_26182_1_stq_idx = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  T_26182_1_brob_idx = _RAND_515[4:0];
  _RAND_516 = {1{`RANDOM}};
  T_26182_1_pdst = _RAND_516[6:0];
  _RAND_517 = {1{`RANDOM}};
  T_26182_1_pop1 = _RAND_517[6:0];
  _RAND_518 = {1{`RANDOM}};
  T_26182_1_pop2 = _RAND_518[6:0];
  _RAND_519 = {1{`RANDOM}};
  T_26182_1_pop3 = _RAND_519[6:0];
  _RAND_520 = {1{`RANDOM}};
  T_26182_1_prs1_busy = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  T_26182_1_prs2_busy = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  T_26182_1_prs3_busy = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  T_26182_1_stale_pdst = _RAND_523[6:0];
  _RAND_524 = {1{`RANDOM}};
  T_26182_1_exception = _RAND_524[0:0];
  _RAND_525 = {2{`RANDOM}};
  T_26182_1_exc_cause = _RAND_525[63:0];
  _RAND_526 = {1{`RANDOM}};
  T_26182_1_bypassable = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  T_26182_1_mem_cmd = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  T_26182_1_mem_typ = _RAND_528[2:0];
  _RAND_529 = {1{`RANDOM}};
  T_26182_1_is_fence = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  T_26182_1_is_fencei = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  T_26182_1_is_store = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  T_26182_1_is_amo = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  T_26182_1_is_load = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  T_26182_1_is_unique = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  T_26182_1_flush_on_commit = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  T_26182_1_ldst = _RAND_536[5:0];
  _RAND_537 = {1{`RANDOM}};
  T_26182_1_lrs1 = _RAND_537[5:0];
  _RAND_538 = {1{`RANDOM}};
  T_26182_1_lrs2 = _RAND_538[5:0];
  _RAND_539 = {1{`RANDOM}};
  T_26182_1_lrs3 = _RAND_539[5:0];
  _RAND_540 = {1{`RANDOM}};
  T_26182_1_ldst_val = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  T_26182_1_dst_rtype = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  T_26182_1_lrs1_rtype = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  T_26182_1_lrs2_rtype = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  T_26182_1_frs3_en = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  T_26182_1_fp_val = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  T_26182_1_fp_single = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  T_26182_1_xcpt_if = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  T_26182_1_replay_if = _RAND_548[0:0];
  _RAND_549 = {2{`RANDOM}};
  T_26182_1_debug_wdata = _RAND_549[63:0];
  _RAND_550 = {1{`RANDOM}};
  T_26182_1_debug_events_fetch_seq = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  T_26182_2_valid = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  T_26182_2_iw_state = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  T_26182_2_uopc = _RAND_553[8:0];
  _RAND_554 = {1{`RANDOM}};
  T_26182_2_inst = _RAND_554[31:0];
  _RAND_555 = {2{`RANDOM}};
  T_26182_2_pc = _RAND_555[39:0];
  _RAND_556 = {1{`RANDOM}};
  T_26182_2_fu_code = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  T_26182_2_ctrl_br_type = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  T_26182_2_ctrl_op1_sel = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  T_26182_2_ctrl_op2_sel = _RAND_559[2:0];
  _RAND_560 = {1{`RANDOM}};
  T_26182_2_ctrl_imm_sel = _RAND_560[2:0];
  _RAND_561 = {1{`RANDOM}};
  T_26182_2_ctrl_op_fcn = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  T_26182_2_ctrl_fcn_dw = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  T_26182_2_ctrl_rf_wen = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  T_26182_2_ctrl_csr_cmd = _RAND_564[2:0];
  _RAND_565 = {1{`RANDOM}};
  T_26182_2_ctrl_is_load = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  T_26182_2_ctrl_is_sta = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  T_26182_2_ctrl_is_std = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  T_26182_2_wakeup_delay = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  T_26182_2_allocate_brtag = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  T_26182_2_is_br_or_jmp = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  T_26182_2_is_jump = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  T_26182_2_is_jal = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  T_26182_2_is_ret = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  T_26182_2_is_call = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  T_26182_2_br_mask = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  T_26182_2_br_tag = _RAND_576[2:0];
  _RAND_577 = {1{`RANDOM}};
  T_26182_2_br_prediction_bpd_predict_val = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  T_26182_2_br_prediction_bpd_predict_taken = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  T_26182_2_br_prediction_btb_hit = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  T_26182_2_br_prediction_btb_predicted = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  T_26182_2_br_prediction_is_br_or_jalr = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  T_26182_2_stat_brjmp_mispredicted = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  T_26182_2_stat_btb_made_pred = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  T_26182_2_stat_btb_mispredicted = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  T_26182_2_stat_bpd_made_pred = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  T_26182_2_stat_bpd_mispredicted = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  T_26182_2_fetch_pc_lob = _RAND_587[2:0];
  _RAND_588 = {1{`RANDOM}};
  T_26182_2_imm_packed = _RAND_588[19:0];
  _RAND_589 = {1{`RANDOM}};
  T_26182_2_csr_addr = _RAND_589[11:0];
  _RAND_590 = {1{`RANDOM}};
  T_26182_2_rob_idx = _RAND_590[5:0];
  _RAND_591 = {1{`RANDOM}};
  T_26182_2_ldq_idx = _RAND_591[3:0];
  _RAND_592 = {1{`RANDOM}};
  T_26182_2_stq_idx = _RAND_592[3:0];
  _RAND_593 = {1{`RANDOM}};
  T_26182_2_brob_idx = _RAND_593[4:0];
  _RAND_594 = {1{`RANDOM}};
  T_26182_2_pdst = _RAND_594[6:0];
  _RAND_595 = {1{`RANDOM}};
  T_26182_2_pop1 = _RAND_595[6:0];
  _RAND_596 = {1{`RANDOM}};
  T_26182_2_pop2 = _RAND_596[6:0];
  _RAND_597 = {1{`RANDOM}};
  T_26182_2_pop3 = _RAND_597[6:0];
  _RAND_598 = {1{`RANDOM}};
  T_26182_2_prs1_busy = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  T_26182_2_prs2_busy = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  T_26182_2_prs3_busy = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  T_26182_2_stale_pdst = _RAND_601[6:0];
  _RAND_602 = {1{`RANDOM}};
  T_26182_2_exception = _RAND_602[0:0];
  _RAND_603 = {2{`RANDOM}};
  T_26182_2_exc_cause = _RAND_603[63:0];
  _RAND_604 = {1{`RANDOM}};
  T_26182_2_bypassable = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  T_26182_2_mem_cmd = _RAND_605[3:0];
  _RAND_606 = {1{`RANDOM}};
  T_26182_2_mem_typ = _RAND_606[2:0];
  _RAND_607 = {1{`RANDOM}};
  T_26182_2_is_fence = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  T_26182_2_is_fencei = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  T_26182_2_is_store = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  T_26182_2_is_amo = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  T_26182_2_is_load = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  T_26182_2_is_unique = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  T_26182_2_flush_on_commit = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  T_26182_2_ldst = _RAND_614[5:0];
  _RAND_615 = {1{`RANDOM}};
  T_26182_2_lrs1 = _RAND_615[5:0];
  _RAND_616 = {1{`RANDOM}};
  T_26182_2_lrs2 = _RAND_616[5:0];
  _RAND_617 = {1{`RANDOM}};
  T_26182_2_lrs3 = _RAND_617[5:0];
  _RAND_618 = {1{`RANDOM}};
  T_26182_2_ldst_val = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  T_26182_2_dst_rtype = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  T_26182_2_lrs1_rtype = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  T_26182_2_lrs2_rtype = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  T_26182_2_frs3_en = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  T_26182_2_fp_val = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  T_26182_2_fp_single = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  T_26182_2_xcpt_if = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  T_26182_2_replay_if = _RAND_626[0:0];
  _RAND_627 = {2{`RANDOM}};
  T_26182_2_debug_wdata = _RAND_627[63:0];
  _RAND_628 = {1{`RANDOM}};
  T_26182_2_debug_events_fetch_seq = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  T_26182_3_valid = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  T_26182_3_iw_state = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  T_26182_3_uopc = _RAND_631[8:0];
  _RAND_632 = {1{`RANDOM}};
  T_26182_3_inst = _RAND_632[31:0];
  _RAND_633 = {2{`RANDOM}};
  T_26182_3_pc = _RAND_633[39:0];
  _RAND_634 = {1{`RANDOM}};
  T_26182_3_fu_code = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  T_26182_3_ctrl_br_type = _RAND_635[3:0];
  _RAND_636 = {1{`RANDOM}};
  T_26182_3_ctrl_op1_sel = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  T_26182_3_ctrl_op2_sel = _RAND_637[2:0];
  _RAND_638 = {1{`RANDOM}};
  T_26182_3_ctrl_imm_sel = _RAND_638[2:0];
  _RAND_639 = {1{`RANDOM}};
  T_26182_3_ctrl_op_fcn = _RAND_639[3:0];
  _RAND_640 = {1{`RANDOM}};
  T_26182_3_ctrl_fcn_dw = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  T_26182_3_ctrl_rf_wen = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  T_26182_3_ctrl_csr_cmd = _RAND_642[2:0];
  _RAND_643 = {1{`RANDOM}};
  T_26182_3_ctrl_is_load = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  T_26182_3_ctrl_is_sta = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  T_26182_3_ctrl_is_std = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  T_26182_3_wakeup_delay = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  T_26182_3_allocate_brtag = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  T_26182_3_is_br_or_jmp = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  T_26182_3_is_jump = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  T_26182_3_is_jal = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  T_26182_3_is_ret = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  T_26182_3_is_call = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  T_26182_3_br_mask = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  T_26182_3_br_tag = _RAND_654[2:0];
  _RAND_655 = {1{`RANDOM}};
  T_26182_3_br_prediction_bpd_predict_val = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  T_26182_3_br_prediction_bpd_predict_taken = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  T_26182_3_br_prediction_btb_hit = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  T_26182_3_br_prediction_btb_predicted = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  T_26182_3_br_prediction_is_br_or_jalr = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  T_26182_3_stat_brjmp_mispredicted = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  T_26182_3_stat_btb_made_pred = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  T_26182_3_stat_btb_mispredicted = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  T_26182_3_stat_bpd_made_pred = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  T_26182_3_stat_bpd_mispredicted = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  T_26182_3_fetch_pc_lob = _RAND_665[2:0];
  _RAND_666 = {1{`RANDOM}};
  T_26182_3_imm_packed = _RAND_666[19:0];
  _RAND_667 = {1{`RANDOM}};
  T_26182_3_csr_addr = _RAND_667[11:0];
  _RAND_668 = {1{`RANDOM}};
  T_26182_3_rob_idx = _RAND_668[5:0];
  _RAND_669 = {1{`RANDOM}};
  T_26182_3_ldq_idx = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  T_26182_3_stq_idx = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  T_26182_3_brob_idx = _RAND_671[4:0];
  _RAND_672 = {1{`RANDOM}};
  T_26182_3_pdst = _RAND_672[6:0];
  _RAND_673 = {1{`RANDOM}};
  T_26182_3_pop1 = _RAND_673[6:0];
  _RAND_674 = {1{`RANDOM}};
  T_26182_3_pop2 = _RAND_674[6:0];
  _RAND_675 = {1{`RANDOM}};
  T_26182_3_pop3 = _RAND_675[6:0];
  _RAND_676 = {1{`RANDOM}};
  T_26182_3_prs1_busy = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  T_26182_3_prs2_busy = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  T_26182_3_prs3_busy = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  T_26182_3_stale_pdst = _RAND_679[6:0];
  _RAND_680 = {1{`RANDOM}};
  T_26182_3_exception = _RAND_680[0:0];
  _RAND_681 = {2{`RANDOM}};
  T_26182_3_exc_cause = _RAND_681[63:0];
  _RAND_682 = {1{`RANDOM}};
  T_26182_3_bypassable = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  T_26182_3_mem_cmd = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  T_26182_3_mem_typ = _RAND_684[2:0];
  _RAND_685 = {1{`RANDOM}};
  T_26182_3_is_fence = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  T_26182_3_is_fencei = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  T_26182_3_is_store = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  T_26182_3_is_amo = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  T_26182_3_is_load = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  T_26182_3_is_unique = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  T_26182_3_flush_on_commit = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  T_26182_3_ldst = _RAND_692[5:0];
  _RAND_693 = {1{`RANDOM}};
  T_26182_3_lrs1 = _RAND_693[5:0];
  _RAND_694 = {1{`RANDOM}};
  T_26182_3_lrs2 = _RAND_694[5:0];
  _RAND_695 = {1{`RANDOM}};
  T_26182_3_lrs3 = _RAND_695[5:0];
  _RAND_696 = {1{`RANDOM}};
  T_26182_3_ldst_val = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  T_26182_3_dst_rtype = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  T_26182_3_lrs1_rtype = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  T_26182_3_lrs2_rtype = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  T_26182_3_frs3_en = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  T_26182_3_fp_val = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  T_26182_3_fp_single = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  T_26182_3_xcpt_if = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  T_26182_3_replay_if = _RAND_704[0:0];
  _RAND_705 = {2{`RANDOM}};
  T_26182_3_debug_wdata = _RAND_705[63:0];
  _RAND_706 = {1{`RANDOM}};
  T_26182_3_debug_events_fetch_seq = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  T_26182_4_valid = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  T_26182_4_iw_state = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  T_26182_4_uopc = _RAND_709[8:0];
  _RAND_710 = {1{`RANDOM}};
  T_26182_4_inst = _RAND_710[31:0];
  _RAND_711 = {2{`RANDOM}};
  T_26182_4_pc = _RAND_711[39:0];
  _RAND_712 = {1{`RANDOM}};
  T_26182_4_fu_code = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  T_26182_4_ctrl_br_type = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  T_26182_4_ctrl_op1_sel = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  T_26182_4_ctrl_op2_sel = _RAND_715[2:0];
  _RAND_716 = {1{`RANDOM}};
  T_26182_4_ctrl_imm_sel = _RAND_716[2:0];
  _RAND_717 = {1{`RANDOM}};
  T_26182_4_ctrl_op_fcn = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  T_26182_4_ctrl_fcn_dw = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  T_26182_4_ctrl_rf_wen = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  T_26182_4_ctrl_csr_cmd = _RAND_720[2:0];
  _RAND_721 = {1{`RANDOM}};
  T_26182_4_ctrl_is_load = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  T_26182_4_ctrl_is_sta = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  T_26182_4_ctrl_is_std = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  T_26182_4_wakeup_delay = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  T_26182_4_allocate_brtag = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  T_26182_4_is_br_or_jmp = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  T_26182_4_is_jump = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  T_26182_4_is_jal = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  T_26182_4_is_ret = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  T_26182_4_is_call = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  T_26182_4_br_mask = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  T_26182_4_br_tag = _RAND_732[2:0];
  _RAND_733 = {1{`RANDOM}};
  T_26182_4_br_prediction_bpd_predict_val = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  T_26182_4_br_prediction_bpd_predict_taken = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  T_26182_4_br_prediction_btb_hit = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  T_26182_4_br_prediction_btb_predicted = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  T_26182_4_br_prediction_is_br_or_jalr = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  T_26182_4_stat_brjmp_mispredicted = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  T_26182_4_stat_btb_made_pred = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  T_26182_4_stat_btb_mispredicted = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  T_26182_4_stat_bpd_made_pred = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  T_26182_4_stat_bpd_mispredicted = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  T_26182_4_fetch_pc_lob = _RAND_743[2:0];
  _RAND_744 = {1{`RANDOM}};
  T_26182_4_imm_packed = _RAND_744[19:0];
  _RAND_745 = {1{`RANDOM}};
  T_26182_4_csr_addr = _RAND_745[11:0];
  _RAND_746 = {1{`RANDOM}};
  T_26182_4_rob_idx = _RAND_746[5:0];
  _RAND_747 = {1{`RANDOM}};
  T_26182_4_ldq_idx = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  T_26182_4_stq_idx = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  T_26182_4_brob_idx = _RAND_749[4:0];
  _RAND_750 = {1{`RANDOM}};
  T_26182_4_pdst = _RAND_750[6:0];
  _RAND_751 = {1{`RANDOM}};
  T_26182_4_pop1 = _RAND_751[6:0];
  _RAND_752 = {1{`RANDOM}};
  T_26182_4_pop2 = _RAND_752[6:0];
  _RAND_753 = {1{`RANDOM}};
  T_26182_4_pop3 = _RAND_753[6:0];
  _RAND_754 = {1{`RANDOM}};
  T_26182_4_prs1_busy = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  T_26182_4_prs2_busy = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  T_26182_4_prs3_busy = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  T_26182_4_stale_pdst = _RAND_757[6:0];
  _RAND_758 = {1{`RANDOM}};
  T_26182_4_exception = _RAND_758[0:0];
  _RAND_759 = {2{`RANDOM}};
  T_26182_4_exc_cause = _RAND_759[63:0];
  _RAND_760 = {1{`RANDOM}};
  T_26182_4_bypassable = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  T_26182_4_mem_cmd = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  T_26182_4_mem_typ = _RAND_762[2:0];
  _RAND_763 = {1{`RANDOM}};
  T_26182_4_is_fence = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  T_26182_4_is_fencei = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  T_26182_4_is_store = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  T_26182_4_is_amo = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  T_26182_4_is_load = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  T_26182_4_is_unique = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  T_26182_4_flush_on_commit = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  T_26182_4_ldst = _RAND_770[5:0];
  _RAND_771 = {1{`RANDOM}};
  T_26182_4_lrs1 = _RAND_771[5:0];
  _RAND_772 = {1{`RANDOM}};
  T_26182_4_lrs2 = _RAND_772[5:0];
  _RAND_773 = {1{`RANDOM}};
  T_26182_4_lrs3 = _RAND_773[5:0];
  _RAND_774 = {1{`RANDOM}};
  T_26182_4_ldst_val = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  T_26182_4_dst_rtype = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  T_26182_4_lrs1_rtype = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  T_26182_4_lrs2_rtype = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  T_26182_4_frs3_en = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  T_26182_4_fp_val = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  T_26182_4_fp_single = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  T_26182_4_xcpt_if = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  T_26182_4_replay_if = _RAND_782[0:0];
  _RAND_783 = {2{`RANDOM}};
  T_26182_4_debug_wdata = _RAND_783[63:0];
  _RAND_784 = {1{`RANDOM}};
  T_26182_4_debug_events_fetch_seq = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  T_26182_5_valid = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  T_26182_5_iw_state = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  T_26182_5_uopc = _RAND_787[8:0];
  _RAND_788 = {1{`RANDOM}};
  T_26182_5_inst = _RAND_788[31:0];
  _RAND_789 = {2{`RANDOM}};
  T_26182_5_pc = _RAND_789[39:0];
  _RAND_790 = {1{`RANDOM}};
  T_26182_5_fu_code = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  T_26182_5_ctrl_br_type = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  T_26182_5_ctrl_op1_sel = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  T_26182_5_ctrl_op2_sel = _RAND_793[2:0];
  _RAND_794 = {1{`RANDOM}};
  T_26182_5_ctrl_imm_sel = _RAND_794[2:0];
  _RAND_795 = {1{`RANDOM}};
  T_26182_5_ctrl_op_fcn = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  T_26182_5_ctrl_fcn_dw = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  T_26182_5_ctrl_rf_wen = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  T_26182_5_ctrl_csr_cmd = _RAND_798[2:0];
  _RAND_799 = {1{`RANDOM}};
  T_26182_5_ctrl_is_load = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  T_26182_5_ctrl_is_sta = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  T_26182_5_ctrl_is_std = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  T_26182_5_wakeup_delay = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  T_26182_5_allocate_brtag = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  T_26182_5_is_br_or_jmp = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  T_26182_5_is_jump = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  T_26182_5_is_jal = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  T_26182_5_is_ret = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  T_26182_5_is_call = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  T_26182_5_br_mask = _RAND_809[7:0];
  _RAND_810 = {1{`RANDOM}};
  T_26182_5_br_tag = _RAND_810[2:0];
  _RAND_811 = {1{`RANDOM}};
  T_26182_5_br_prediction_bpd_predict_val = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  T_26182_5_br_prediction_bpd_predict_taken = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  T_26182_5_br_prediction_btb_hit = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  T_26182_5_br_prediction_btb_predicted = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  T_26182_5_br_prediction_is_br_or_jalr = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  T_26182_5_stat_brjmp_mispredicted = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  T_26182_5_stat_btb_made_pred = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  T_26182_5_stat_btb_mispredicted = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  T_26182_5_stat_bpd_made_pred = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  T_26182_5_stat_bpd_mispredicted = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  T_26182_5_fetch_pc_lob = _RAND_821[2:0];
  _RAND_822 = {1{`RANDOM}};
  T_26182_5_imm_packed = _RAND_822[19:0];
  _RAND_823 = {1{`RANDOM}};
  T_26182_5_csr_addr = _RAND_823[11:0];
  _RAND_824 = {1{`RANDOM}};
  T_26182_5_rob_idx = _RAND_824[5:0];
  _RAND_825 = {1{`RANDOM}};
  T_26182_5_ldq_idx = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  T_26182_5_stq_idx = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  T_26182_5_brob_idx = _RAND_827[4:0];
  _RAND_828 = {1{`RANDOM}};
  T_26182_5_pdst = _RAND_828[6:0];
  _RAND_829 = {1{`RANDOM}};
  T_26182_5_pop1 = _RAND_829[6:0];
  _RAND_830 = {1{`RANDOM}};
  T_26182_5_pop2 = _RAND_830[6:0];
  _RAND_831 = {1{`RANDOM}};
  T_26182_5_pop3 = _RAND_831[6:0];
  _RAND_832 = {1{`RANDOM}};
  T_26182_5_prs1_busy = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  T_26182_5_prs2_busy = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  T_26182_5_prs3_busy = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  T_26182_5_stale_pdst = _RAND_835[6:0];
  _RAND_836 = {1{`RANDOM}};
  T_26182_5_exception = _RAND_836[0:0];
  _RAND_837 = {2{`RANDOM}};
  T_26182_5_exc_cause = _RAND_837[63:0];
  _RAND_838 = {1{`RANDOM}};
  T_26182_5_bypassable = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  T_26182_5_mem_cmd = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  T_26182_5_mem_typ = _RAND_840[2:0];
  _RAND_841 = {1{`RANDOM}};
  T_26182_5_is_fence = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  T_26182_5_is_fencei = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  T_26182_5_is_store = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  T_26182_5_is_amo = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  T_26182_5_is_load = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  T_26182_5_is_unique = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  T_26182_5_flush_on_commit = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  T_26182_5_ldst = _RAND_848[5:0];
  _RAND_849 = {1{`RANDOM}};
  T_26182_5_lrs1 = _RAND_849[5:0];
  _RAND_850 = {1{`RANDOM}};
  T_26182_5_lrs2 = _RAND_850[5:0];
  _RAND_851 = {1{`RANDOM}};
  T_26182_5_lrs3 = _RAND_851[5:0];
  _RAND_852 = {1{`RANDOM}};
  T_26182_5_ldst_val = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  T_26182_5_dst_rtype = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  T_26182_5_lrs1_rtype = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  T_26182_5_lrs2_rtype = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  T_26182_5_frs3_en = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  T_26182_5_fp_val = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  T_26182_5_fp_single = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  T_26182_5_xcpt_if = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  T_26182_5_replay_if = _RAND_860[0:0];
  _RAND_861 = {2{`RANDOM}};
  T_26182_5_debug_wdata = _RAND_861[63:0];
  _RAND_862 = {1{`RANDOM}};
  T_26182_5_debug_events_fetch_seq = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  T_26182_6_valid = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  T_26182_6_iw_state = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  T_26182_6_uopc = _RAND_865[8:0];
  _RAND_866 = {1{`RANDOM}};
  T_26182_6_inst = _RAND_866[31:0];
  _RAND_867 = {2{`RANDOM}};
  T_26182_6_pc = _RAND_867[39:0];
  _RAND_868 = {1{`RANDOM}};
  T_26182_6_fu_code = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  T_26182_6_ctrl_br_type = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  T_26182_6_ctrl_op1_sel = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  T_26182_6_ctrl_op2_sel = _RAND_871[2:0];
  _RAND_872 = {1{`RANDOM}};
  T_26182_6_ctrl_imm_sel = _RAND_872[2:0];
  _RAND_873 = {1{`RANDOM}};
  T_26182_6_ctrl_op_fcn = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  T_26182_6_ctrl_fcn_dw = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  T_26182_6_ctrl_rf_wen = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  T_26182_6_ctrl_csr_cmd = _RAND_876[2:0];
  _RAND_877 = {1{`RANDOM}};
  T_26182_6_ctrl_is_load = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  T_26182_6_ctrl_is_sta = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  T_26182_6_ctrl_is_std = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  T_26182_6_wakeup_delay = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  T_26182_6_allocate_brtag = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  T_26182_6_is_br_or_jmp = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  T_26182_6_is_jump = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  T_26182_6_is_jal = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  T_26182_6_is_ret = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  T_26182_6_is_call = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  T_26182_6_br_mask = _RAND_887[7:0];
  _RAND_888 = {1{`RANDOM}};
  T_26182_6_br_tag = _RAND_888[2:0];
  _RAND_889 = {1{`RANDOM}};
  T_26182_6_br_prediction_bpd_predict_val = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  T_26182_6_br_prediction_bpd_predict_taken = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  T_26182_6_br_prediction_btb_hit = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  T_26182_6_br_prediction_btb_predicted = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  T_26182_6_br_prediction_is_br_or_jalr = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  T_26182_6_stat_brjmp_mispredicted = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  T_26182_6_stat_btb_made_pred = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  T_26182_6_stat_btb_mispredicted = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  T_26182_6_stat_bpd_made_pred = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  T_26182_6_stat_bpd_mispredicted = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  T_26182_6_fetch_pc_lob = _RAND_899[2:0];
  _RAND_900 = {1{`RANDOM}};
  T_26182_6_imm_packed = _RAND_900[19:0];
  _RAND_901 = {1{`RANDOM}};
  T_26182_6_csr_addr = _RAND_901[11:0];
  _RAND_902 = {1{`RANDOM}};
  T_26182_6_rob_idx = _RAND_902[5:0];
  _RAND_903 = {1{`RANDOM}};
  T_26182_6_ldq_idx = _RAND_903[3:0];
  _RAND_904 = {1{`RANDOM}};
  T_26182_6_stq_idx = _RAND_904[3:0];
  _RAND_905 = {1{`RANDOM}};
  T_26182_6_brob_idx = _RAND_905[4:0];
  _RAND_906 = {1{`RANDOM}};
  T_26182_6_pdst = _RAND_906[6:0];
  _RAND_907 = {1{`RANDOM}};
  T_26182_6_pop1 = _RAND_907[6:0];
  _RAND_908 = {1{`RANDOM}};
  T_26182_6_pop2 = _RAND_908[6:0];
  _RAND_909 = {1{`RANDOM}};
  T_26182_6_pop3 = _RAND_909[6:0];
  _RAND_910 = {1{`RANDOM}};
  T_26182_6_prs1_busy = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  T_26182_6_prs2_busy = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  T_26182_6_prs3_busy = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  T_26182_6_stale_pdst = _RAND_913[6:0];
  _RAND_914 = {1{`RANDOM}};
  T_26182_6_exception = _RAND_914[0:0];
  _RAND_915 = {2{`RANDOM}};
  T_26182_6_exc_cause = _RAND_915[63:0];
  _RAND_916 = {1{`RANDOM}};
  T_26182_6_bypassable = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  T_26182_6_mem_cmd = _RAND_917[3:0];
  _RAND_918 = {1{`RANDOM}};
  T_26182_6_mem_typ = _RAND_918[2:0];
  _RAND_919 = {1{`RANDOM}};
  T_26182_6_is_fence = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  T_26182_6_is_fencei = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  T_26182_6_is_store = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  T_26182_6_is_amo = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  T_26182_6_is_load = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  T_26182_6_is_unique = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  T_26182_6_flush_on_commit = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  T_26182_6_ldst = _RAND_926[5:0];
  _RAND_927 = {1{`RANDOM}};
  T_26182_6_lrs1 = _RAND_927[5:0];
  _RAND_928 = {1{`RANDOM}};
  T_26182_6_lrs2 = _RAND_928[5:0];
  _RAND_929 = {1{`RANDOM}};
  T_26182_6_lrs3 = _RAND_929[5:0];
  _RAND_930 = {1{`RANDOM}};
  T_26182_6_ldst_val = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  T_26182_6_dst_rtype = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  T_26182_6_lrs1_rtype = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  T_26182_6_lrs2_rtype = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  T_26182_6_frs3_en = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  T_26182_6_fp_val = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  T_26182_6_fp_single = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  T_26182_6_xcpt_if = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  T_26182_6_replay_if = _RAND_938[0:0];
  _RAND_939 = {2{`RANDOM}};
  T_26182_6_debug_wdata = _RAND_939[63:0];
  _RAND_940 = {1{`RANDOM}};
  T_26182_6_debug_events_fetch_seq = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  T_26182_7_valid = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  T_26182_7_iw_state = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  T_26182_7_uopc = _RAND_943[8:0];
  _RAND_944 = {1{`RANDOM}};
  T_26182_7_inst = _RAND_944[31:0];
  _RAND_945 = {2{`RANDOM}};
  T_26182_7_pc = _RAND_945[39:0];
  _RAND_946 = {1{`RANDOM}};
  T_26182_7_fu_code = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  T_26182_7_ctrl_br_type = _RAND_947[3:0];
  _RAND_948 = {1{`RANDOM}};
  T_26182_7_ctrl_op1_sel = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  T_26182_7_ctrl_op2_sel = _RAND_949[2:0];
  _RAND_950 = {1{`RANDOM}};
  T_26182_7_ctrl_imm_sel = _RAND_950[2:0];
  _RAND_951 = {1{`RANDOM}};
  T_26182_7_ctrl_op_fcn = _RAND_951[3:0];
  _RAND_952 = {1{`RANDOM}};
  T_26182_7_ctrl_fcn_dw = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  T_26182_7_ctrl_rf_wen = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  T_26182_7_ctrl_csr_cmd = _RAND_954[2:0];
  _RAND_955 = {1{`RANDOM}};
  T_26182_7_ctrl_is_load = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  T_26182_7_ctrl_is_sta = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  T_26182_7_ctrl_is_std = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  T_26182_7_wakeup_delay = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  T_26182_7_allocate_brtag = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  T_26182_7_is_br_or_jmp = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  T_26182_7_is_jump = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  T_26182_7_is_jal = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  T_26182_7_is_ret = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  T_26182_7_is_call = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  T_26182_7_br_mask = _RAND_965[7:0];
  _RAND_966 = {1{`RANDOM}};
  T_26182_7_br_tag = _RAND_966[2:0];
  _RAND_967 = {1{`RANDOM}};
  T_26182_7_br_prediction_bpd_predict_val = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  T_26182_7_br_prediction_bpd_predict_taken = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  T_26182_7_br_prediction_btb_hit = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  T_26182_7_br_prediction_btb_predicted = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  T_26182_7_br_prediction_is_br_or_jalr = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  T_26182_7_stat_brjmp_mispredicted = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  T_26182_7_stat_btb_made_pred = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  T_26182_7_stat_btb_mispredicted = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  T_26182_7_stat_bpd_made_pred = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  T_26182_7_stat_bpd_mispredicted = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  T_26182_7_fetch_pc_lob = _RAND_977[2:0];
  _RAND_978 = {1{`RANDOM}};
  T_26182_7_imm_packed = _RAND_978[19:0];
  _RAND_979 = {1{`RANDOM}};
  T_26182_7_csr_addr = _RAND_979[11:0];
  _RAND_980 = {1{`RANDOM}};
  T_26182_7_rob_idx = _RAND_980[5:0];
  _RAND_981 = {1{`RANDOM}};
  T_26182_7_ldq_idx = _RAND_981[3:0];
  _RAND_982 = {1{`RANDOM}};
  T_26182_7_stq_idx = _RAND_982[3:0];
  _RAND_983 = {1{`RANDOM}};
  T_26182_7_brob_idx = _RAND_983[4:0];
  _RAND_984 = {1{`RANDOM}};
  T_26182_7_pdst = _RAND_984[6:0];
  _RAND_985 = {1{`RANDOM}};
  T_26182_7_pop1 = _RAND_985[6:0];
  _RAND_986 = {1{`RANDOM}};
  T_26182_7_pop2 = _RAND_986[6:0];
  _RAND_987 = {1{`RANDOM}};
  T_26182_7_pop3 = _RAND_987[6:0];
  _RAND_988 = {1{`RANDOM}};
  T_26182_7_prs1_busy = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  T_26182_7_prs2_busy = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  T_26182_7_prs3_busy = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  T_26182_7_stale_pdst = _RAND_991[6:0];
  _RAND_992 = {1{`RANDOM}};
  T_26182_7_exception = _RAND_992[0:0];
  _RAND_993 = {2{`RANDOM}};
  T_26182_7_exc_cause = _RAND_993[63:0];
  _RAND_994 = {1{`RANDOM}};
  T_26182_7_bypassable = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  T_26182_7_mem_cmd = _RAND_995[3:0];
  _RAND_996 = {1{`RANDOM}};
  T_26182_7_mem_typ = _RAND_996[2:0];
  _RAND_997 = {1{`RANDOM}};
  T_26182_7_is_fence = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  T_26182_7_is_fencei = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  T_26182_7_is_store = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  T_26182_7_is_amo = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  T_26182_7_is_load = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  T_26182_7_is_unique = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  T_26182_7_flush_on_commit = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  T_26182_7_ldst = _RAND_1004[5:0];
  _RAND_1005 = {1{`RANDOM}};
  T_26182_7_lrs1 = _RAND_1005[5:0];
  _RAND_1006 = {1{`RANDOM}};
  T_26182_7_lrs2 = _RAND_1006[5:0];
  _RAND_1007 = {1{`RANDOM}};
  T_26182_7_lrs3 = _RAND_1007[5:0];
  _RAND_1008 = {1{`RANDOM}};
  T_26182_7_ldst_val = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  T_26182_7_dst_rtype = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  T_26182_7_lrs1_rtype = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  T_26182_7_lrs2_rtype = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  T_26182_7_frs3_en = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  T_26182_7_fp_val = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  T_26182_7_fp_single = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  T_26182_7_xcpt_if = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  T_26182_7_replay_if = _RAND_1016[0:0];
  _RAND_1017 = {2{`RANDOM}};
  T_26182_7_debug_wdata = _RAND_1017[63:0];
  _RAND_1018 = {1{`RANDOM}};
  T_26182_7_debug_events_fetch_seq = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  T_26182_8_valid = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  T_26182_8_iw_state = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  T_26182_8_uopc = _RAND_1021[8:0];
  _RAND_1022 = {1{`RANDOM}};
  T_26182_8_inst = _RAND_1022[31:0];
  _RAND_1023 = {2{`RANDOM}};
  T_26182_8_pc = _RAND_1023[39:0];
  _RAND_1024 = {1{`RANDOM}};
  T_26182_8_fu_code = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  T_26182_8_ctrl_br_type = _RAND_1025[3:0];
  _RAND_1026 = {1{`RANDOM}};
  T_26182_8_ctrl_op1_sel = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  T_26182_8_ctrl_op2_sel = _RAND_1027[2:0];
  _RAND_1028 = {1{`RANDOM}};
  T_26182_8_ctrl_imm_sel = _RAND_1028[2:0];
  _RAND_1029 = {1{`RANDOM}};
  T_26182_8_ctrl_op_fcn = _RAND_1029[3:0];
  _RAND_1030 = {1{`RANDOM}};
  T_26182_8_ctrl_fcn_dw = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  T_26182_8_ctrl_rf_wen = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  T_26182_8_ctrl_csr_cmd = _RAND_1032[2:0];
  _RAND_1033 = {1{`RANDOM}};
  T_26182_8_ctrl_is_load = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  T_26182_8_ctrl_is_sta = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  T_26182_8_ctrl_is_std = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  T_26182_8_wakeup_delay = _RAND_1036[1:0];
  _RAND_1037 = {1{`RANDOM}};
  T_26182_8_allocate_brtag = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  T_26182_8_is_br_or_jmp = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  T_26182_8_is_jump = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  T_26182_8_is_jal = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  T_26182_8_is_ret = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  T_26182_8_is_call = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  T_26182_8_br_mask = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  T_26182_8_br_tag = _RAND_1044[2:0];
  _RAND_1045 = {1{`RANDOM}};
  T_26182_8_br_prediction_bpd_predict_val = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  T_26182_8_br_prediction_bpd_predict_taken = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  T_26182_8_br_prediction_btb_hit = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  T_26182_8_br_prediction_btb_predicted = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  T_26182_8_br_prediction_is_br_or_jalr = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  T_26182_8_stat_brjmp_mispredicted = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  T_26182_8_stat_btb_made_pred = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  T_26182_8_stat_btb_mispredicted = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  T_26182_8_stat_bpd_made_pred = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  T_26182_8_stat_bpd_mispredicted = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  T_26182_8_fetch_pc_lob = _RAND_1055[2:0];
  _RAND_1056 = {1{`RANDOM}};
  T_26182_8_imm_packed = _RAND_1056[19:0];
  _RAND_1057 = {1{`RANDOM}};
  T_26182_8_csr_addr = _RAND_1057[11:0];
  _RAND_1058 = {1{`RANDOM}};
  T_26182_8_rob_idx = _RAND_1058[5:0];
  _RAND_1059 = {1{`RANDOM}};
  T_26182_8_ldq_idx = _RAND_1059[3:0];
  _RAND_1060 = {1{`RANDOM}};
  T_26182_8_stq_idx = _RAND_1060[3:0];
  _RAND_1061 = {1{`RANDOM}};
  T_26182_8_brob_idx = _RAND_1061[4:0];
  _RAND_1062 = {1{`RANDOM}};
  T_26182_8_pdst = _RAND_1062[6:0];
  _RAND_1063 = {1{`RANDOM}};
  T_26182_8_pop1 = _RAND_1063[6:0];
  _RAND_1064 = {1{`RANDOM}};
  T_26182_8_pop2 = _RAND_1064[6:0];
  _RAND_1065 = {1{`RANDOM}};
  T_26182_8_pop3 = _RAND_1065[6:0];
  _RAND_1066 = {1{`RANDOM}};
  T_26182_8_prs1_busy = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  T_26182_8_prs2_busy = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  T_26182_8_prs3_busy = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  T_26182_8_stale_pdst = _RAND_1069[6:0];
  _RAND_1070 = {1{`RANDOM}};
  T_26182_8_exception = _RAND_1070[0:0];
  _RAND_1071 = {2{`RANDOM}};
  T_26182_8_exc_cause = _RAND_1071[63:0];
  _RAND_1072 = {1{`RANDOM}};
  T_26182_8_bypassable = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  T_26182_8_mem_cmd = _RAND_1073[3:0];
  _RAND_1074 = {1{`RANDOM}};
  T_26182_8_mem_typ = _RAND_1074[2:0];
  _RAND_1075 = {1{`RANDOM}};
  T_26182_8_is_fence = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  T_26182_8_is_fencei = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  T_26182_8_is_store = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  T_26182_8_is_amo = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  T_26182_8_is_load = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  T_26182_8_is_unique = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  T_26182_8_flush_on_commit = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  T_26182_8_ldst = _RAND_1082[5:0];
  _RAND_1083 = {1{`RANDOM}};
  T_26182_8_lrs1 = _RAND_1083[5:0];
  _RAND_1084 = {1{`RANDOM}};
  T_26182_8_lrs2 = _RAND_1084[5:0];
  _RAND_1085 = {1{`RANDOM}};
  T_26182_8_lrs3 = _RAND_1085[5:0];
  _RAND_1086 = {1{`RANDOM}};
  T_26182_8_ldst_val = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  T_26182_8_dst_rtype = _RAND_1087[1:0];
  _RAND_1088 = {1{`RANDOM}};
  T_26182_8_lrs1_rtype = _RAND_1088[1:0];
  _RAND_1089 = {1{`RANDOM}};
  T_26182_8_lrs2_rtype = _RAND_1089[1:0];
  _RAND_1090 = {1{`RANDOM}};
  T_26182_8_frs3_en = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  T_26182_8_fp_val = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  T_26182_8_fp_single = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  T_26182_8_xcpt_if = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  T_26182_8_replay_if = _RAND_1094[0:0];
  _RAND_1095 = {2{`RANDOM}};
  T_26182_8_debug_wdata = _RAND_1095[63:0];
  _RAND_1096 = {1{`RANDOM}};
  T_26182_8_debug_events_fetch_seq = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  T_26182_9_valid = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  T_26182_9_iw_state = _RAND_1098[1:0];
  _RAND_1099 = {1{`RANDOM}};
  T_26182_9_uopc = _RAND_1099[8:0];
  _RAND_1100 = {1{`RANDOM}};
  T_26182_9_inst = _RAND_1100[31:0];
  _RAND_1101 = {2{`RANDOM}};
  T_26182_9_pc = _RAND_1101[39:0];
  _RAND_1102 = {1{`RANDOM}};
  T_26182_9_fu_code = _RAND_1102[7:0];
  _RAND_1103 = {1{`RANDOM}};
  T_26182_9_ctrl_br_type = _RAND_1103[3:0];
  _RAND_1104 = {1{`RANDOM}};
  T_26182_9_ctrl_op1_sel = _RAND_1104[1:0];
  _RAND_1105 = {1{`RANDOM}};
  T_26182_9_ctrl_op2_sel = _RAND_1105[2:0];
  _RAND_1106 = {1{`RANDOM}};
  T_26182_9_ctrl_imm_sel = _RAND_1106[2:0];
  _RAND_1107 = {1{`RANDOM}};
  T_26182_9_ctrl_op_fcn = _RAND_1107[3:0];
  _RAND_1108 = {1{`RANDOM}};
  T_26182_9_ctrl_fcn_dw = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  T_26182_9_ctrl_rf_wen = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  T_26182_9_ctrl_csr_cmd = _RAND_1110[2:0];
  _RAND_1111 = {1{`RANDOM}};
  T_26182_9_ctrl_is_load = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  T_26182_9_ctrl_is_sta = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  T_26182_9_ctrl_is_std = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  T_26182_9_wakeup_delay = _RAND_1114[1:0];
  _RAND_1115 = {1{`RANDOM}};
  T_26182_9_allocate_brtag = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  T_26182_9_is_br_or_jmp = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  T_26182_9_is_jump = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  T_26182_9_is_jal = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  T_26182_9_is_ret = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  T_26182_9_is_call = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  T_26182_9_br_mask = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  T_26182_9_br_tag = _RAND_1122[2:0];
  _RAND_1123 = {1{`RANDOM}};
  T_26182_9_br_prediction_bpd_predict_val = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  T_26182_9_br_prediction_bpd_predict_taken = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  T_26182_9_br_prediction_btb_hit = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  T_26182_9_br_prediction_btb_predicted = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  T_26182_9_br_prediction_is_br_or_jalr = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  T_26182_9_stat_brjmp_mispredicted = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  T_26182_9_stat_btb_made_pred = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  T_26182_9_stat_btb_mispredicted = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  T_26182_9_stat_bpd_made_pred = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  T_26182_9_stat_bpd_mispredicted = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  T_26182_9_fetch_pc_lob = _RAND_1133[2:0];
  _RAND_1134 = {1{`RANDOM}};
  T_26182_9_imm_packed = _RAND_1134[19:0];
  _RAND_1135 = {1{`RANDOM}};
  T_26182_9_csr_addr = _RAND_1135[11:0];
  _RAND_1136 = {1{`RANDOM}};
  T_26182_9_rob_idx = _RAND_1136[5:0];
  _RAND_1137 = {1{`RANDOM}};
  T_26182_9_ldq_idx = _RAND_1137[3:0];
  _RAND_1138 = {1{`RANDOM}};
  T_26182_9_stq_idx = _RAND_1138[3:0];
  _RAND_1139 = {1{`RANDOM}};
  T_26182_9_brob_idx = _RAND_1139[4:0];
  _RAND_1140 = {1{`RANDOM}};
  T_26182_9_pdst = _RAND_1140[6:0];
  _RAND_1141 = {1{`RANDOM}};
  T_26182_9_pop1 = _RAND_1141[6:0];
  _RAND_1142 = {1{`RANDOM}};
  T_26182_9_pop2 = _RAND_1142[6:0];
  _RAND_1143 = {1{`RANDOM}};
  T_26182_9_pop3 = _RAND_1143[6:0];
  _RAND_1144 = {1{`RANDOM}};
  T_26182_9_prs1_busy = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  T_26182_9_prs2_busy = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  T_26182_9_prs3_busy = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  T_26182_9_stale_pdst = _RAND_1147[6:0];
  _RAND_1148 = {1{`RANDOM}};
  T_26182_9_exception = _RAND_1148[0:0];
  _RAND_1149 = {2{`RANDOM}};
  T_26182_9_exc_cause = _RAND_1149[63:0];
  _RAND_1150 = {1{`RANDOM}};
  T_26182_9_bypassable = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  T_26182_9_mem_cmd = _RAND_1151[3:0];
  _RAND_1152 = {1{`RANDOM}};
  T_26182_9_mem_typ = _RAND_1152[2:0];
  _RAND_1153 = {1{`RANDOM}};
  T_26182_9_is_fence = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  T_26182_9_is_fencei = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  T_26182_9_is_store = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  T_26182_9_is_amo = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  T_26182_9_is_load = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  T_26182_9_is_unique = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  T_26182_9_flush_on_commit = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  T_26182_9_ldst = _RAND_1160[5:0];
  _RAND_1161 = {1{`RANDOM}};
  T_26182_9_lrs1 = _RAND_1161[5:0];
  _RAND_1162 = {1{`RANDOM}};
  T_26182_9_lrs2 = _RAND_1162[5:0];
  _RAND_1163 = {1{`RANDOM}};
  T_26182_9_lrs3 = _RAND_1163[5:0];
  _RAND_1164 = {1{`RANDOM}};
  T_26182_9_ldst_val = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  T_26182_9_dst_rtype = _RAND_1165[1:0];
  _RAND_1166 = {1{`RANDOM}};
  T_26182_9_lrs1_rtype = _RAND_1166[1:0];
  _RAND_1167 = {1{`RANDOM}};
  T_26182_9_lrs2_rtype = _RAND_1167[1:0];
  _RAND_1168 = {1{`RANDOM}};
  T_26182_9_frs3_en = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  T_26182_9_fp_val = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  T_26182_9_fp_single = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  T_26182_9_xcpt_if = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  T_26182_9_replay_if = _RAND_1172[0:0];
  _RAND_1173 = {2{`RANDOM}};
  T_26182_9_debug_wdata = _RAND_1173[63:0];
  _RAND_1174 = {1{`RANDOM}};
  T_26182_9_debug_events_fetch_seq = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  T_26182_10_valid = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  T_26182_10_iw_state = _RAND_1176[1:0];
  _RAND_1177 = {1{`RANDOM}};
  T_26182_10_uopc = _RAND_1177[8:0];
  _RAND_1178 = {1{`RANDOM}};
  T_26182_10_inst = _RAND_1178[31:0];
  _RAND_1179 = {2{`RANDOM}};
  T_26182_10_pc = _RAND_1179[39:0];
  _RAND_1180 = {1{`RANDOM}};
  T_26182_10_fu_code = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  T_26182_10_ctrl_br_type = _RAND_1181[3:0];
  _RAND_1182 = {1{`RANDOM}};
  T_26182_10_ctrl_op1_sel = _RAND_1182[1:0];
  _RAND_1183 = {1{`RANDOM}};
  T_26182_10_ctrl_op2_sel = _RAND_1183[2:0];
  _RAND_1184 = {1{`RANDOM}};
  T_26182_10_ctrl_imm_sel = _RAND_1184[2:0];
  _RAND_1185 = {1{`RANDOM}};
  T_26182_10_ctrl_op_fcn = _RAND_1185[3:0];
  _RAND_1186 = {1{`RANDOM}};
  T_26182_10_ctrl_fcn_dw = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  T_26182_10_ctrl_rf_wen = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  T_26182_10_ctrl_csr_cmd = _RAND_1188[2:0];
  _RAND_1189 = {1{`RANDOM}};
  T_26182_10_ctrl_is_load = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  T_26182_10_ctrl_is_sta = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  T_26182_10_ctrl_is_std = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  T_26182_10_wakeup_delay = _RAND_1192[1:0];
  _RAND_1193 = {1{`RANDOM}};
  T_26182_10_allocate_brtag = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  T_26182_10_is_br_or_jmp = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  T_26182_10_is_jump = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  T_26182_10_is_jal = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  T_26182_10_is_ret = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  T_26182_10_is_call = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  T_26182_10_br_mask = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  T_26182_10_br_tag = _RAND_1200[2:0];
  _RAND_1201 = {1{`RANDOM}};
  T_26182_10_br_prediction_bpd_predict_val = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  T_26182_10_br_prediction_bpd_predict_taken = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  T_26182_10_br_prediction_btb_hit = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  T_26182_10_br_prediction_btb_predicted = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  T_26182_10_br_prediction_is_br_or_jalr = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  T_26182_10_stat_brjmp_mispredicted = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  T_26182_10_stat_btb_made_pred = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  T_26182_10_stat_btb_mispredicted = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  T_26182_10_stat_bpd_made_pred = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  T_26182_10_stat_bpd_mispredicted = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  T_26182_10_fetch_pc_lob = _RAND_1211[2:0];
  _RAND_1212 = {1{`RANDOM}};
  T_26182_10_imm_packed = _RAND_1212[19:0];
  _RAND_1213 = {1{`RANDOM}};
  T_26182_10_csr_addr = _RAND_1213[11:0];
  _RAND_1214 = {1{`RANDOM}};
  T_26182_10_rob_idx = _RAND_1214[5:0];
  _RAND_1215 = {1{`RANDOM}};
  T_26182_10_ldq_idx = _RAND_1215[3:0];
  _RAND_1216 = {1{`RANDOM}};
  T_26182_10_stq_idx = _RAND_1216[3:0];
  _RAND_1217 = {1{`RANDOM}};
  T_26182_10_brob_idx = _RAND_1217[4:0];
  _RAND_1218 = {1{`RANDOM}};
  T_26182_10_pdst = _RAND_1218[6:0];
  _RAND_1219 = {1{`RANDOM}};
  T_26182_10_pop1 = _RAND_1219[6:0];
  _RAND_1220 = {1{`RANDOM}};
  T_26182_10_pop2 = _RAND_1220[6:0];
  _RAND_1221 = {1{`RANDOM}};
  T_26182_10_pop3 = _RAND_1221[6:0];
  _RAND_1222 = {1{`RANDOM}};
  T_26182_10_prs1_busy = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  T_26182_10_prs2_busy = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  T_26182_10_prs3_busy = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  T_26182_10_stale_pdst = _RAND_1225[6:0];
  _RAND_1226 = {1{`RANDOM}};
  T_26182_10_exception = _RAND_1226[0:0];
  _RAND_1227 = {2{`RANDOM}};
  T_26182_10_exc_cause = _RAND_1227[63:0];
  _RAND_1228 = {1{`RANDOM}};
  T_26182_10_bypassable = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  T_26182_10_mem_cmd = _RAND_1229[3:0];
  _RAND_1230 = {1{`RANDOM}};
  T_26182_10_mem_typ = _RAND_1230[2:0];
  _RAND_1231 = {1{`RANDOM}};
  T_26182_10_is_fence = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  T_26182_10_is_fencei = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  T_26182_10_is_store = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  T_26182_10_is_amo = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  T_26182_10_is_load = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  T_26182_10_is_unique = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  T_26182_10_flush_on_commit = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  T_26182_10_ldst = _RAND_1238[5:0];
  _RAND_1239 = {1{`RANDOM}};
  T_26182_10_lrs1 = _RAND_1239[5:0];
  _RAND_1240 = {1{`RANDOM}};
  T_26182_10_lrs2 = _RAND_1240[5:0];
  _RAND_1241 = {1{`RANDOM}};
  T_26182_10_lrs3 = _RAND_1241[5:0];
  _RAND_1242 = {1{`RANDOM}};
  T_26182_10_ldst_val = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  T_26182_10_dst_rtype = _RAND_1243[1:0];
  _RAND_1244 = {1{`RANDOM}};
  T_26182_10_lrs1_rtype = _RAND_1244[1:0];
  _RAND_1245 = {1{`RANDOM}};
  T_26182_10_lrs2_rtype = _RAND_1245[1:0];
  _RAND_1246 = {1{`RANDOM}};
  T_26182_10_frs3_en = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  T_26182_10_fp_val = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  T_26182_10_fp_single = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  T_26182_10_xcpt_if = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  T_26182_10_replay_if = _RAND_1250[0:0];
  _RAND_1251 = {2{`RANDOM}};
  T_26182_10_debug_wdata = _RAND_1251[63:0];
  _RAND_1252 = {1{`RANDOM}};
  T_26182_10_debug_events_fetch_seq = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  T_26182_11_valid = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  T_26182_11_iw_state = _RAND_1254[1:0];
  _RAND_1255 = {1{`RANDOM}};
  T_26182_11_uopc = _RAND_1255[8:0];
  _RAND_1256 = {1{`RANDOM}};
  T_26182_11_inst = _RAND_1256[31:0];
  _RAND_1257 = {2{`RANDOM}};
  T_26182_11_pc = _RAND_1257[39:0];
  _RAND_1258 = {1{`RANDOM}};
  T_26182_11_fu_code = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  T_26182_11_ctrl_br_type = _RAND_1259[3:0];
  _RAND_1260 = {1{`RANDOM}};
  T_26182_11_ctrl_op1_sel = _RAND_1260[1:0];
  _RAND_1261 = {1{`RANDOM}};
  T_26182_11_ctrl_op2_sel = _RAND_1261[2:0];
  _RAND_1262 = {1{`RANDOM}};
  T_26182_11_ctrl_imm_sel = _RAND_1262[2:0];
  _RAND_1263 = {1{`RANDOM}};
  T_26182_11_ctrl_op_fcn = _RAND_1263[3:0];
  _RAND_1264 = {1{`RANDOM}};
  T_26182_11_ctrl_fcn_dw = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  T_26182_11_ctrl_rf_wen = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  T_26182_11_ctrl_csr_cmd = _RAND_1266[2:0];
  _RAND_1267 = {1{`RANDOM}};
  T_26182_11_ctrl_is_load = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  T_26182_11_ctrl_is_sta = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  T_26182_11_ctrl_is_std = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  T_26182_11_wakeup_delay = _RAND_1270[1:0];
  _RAND_1271 = {1{`RANDOM}};
  T_26182_11_allocate_brtag = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  T_26182_11_is_br_or_jmp = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  T_26182_11_is_jump = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  T_26182_11_is_jal = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  T_26182_11_is_ret = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  T_26182_11_is_call = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  T_26182_11_br_mask = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  T_26182_11_br_tag = _RAND_1278[2:0];
  _RAND_1279 = {1{`RANDOM}};
  T_26182_11_br_prediction_bpd_predict_val = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  T_26182_11_br_prediction_bpd_predict_taken = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  T_26182_11_br_prediction_btb_hit = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  T_26182_11_br_prediction_btb_predicted = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  T_26182_11_br_prediction_is_br_or_jalr = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  T_26182_11_stat_brjmp_mispredicted = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  T_26182_11_stat_btb_made_pred = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  T_26182_11_stat_btb_mispredicted = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  T_26182_11_stat_bpd_made_pred = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  T_26182_11_stat_bpd_mispredicted = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  T_26182_11_fetch_pc_lob = _RAND_1289[2:0];
  _RAND_1290 = {1{`RANDOM}};
  T_26182_11_imm_packed = _RAND_1290[19:0];
  _RAND_1291 = {1{`RANDOM}};
  T_26182_11_csr_addr = _RAND_1291[11:0];
  _RAND_1292 = {1{`RANDOM}};
  T_26182_11_rob_idx = _RAND_1292[5:0];
  _RAND_1293 = {1{`RANDOM}};
  T_26182_11_ldq_idx = _RAND_1293[3:0];
  _RAND_1294 = {1{`RANDOM}};
  T_26182_11_stq_idx = _RAND_1294[3:0];
  _RAND_1295 = {1{`RANDOM}};
  T_26182_11_brob_idx = _RAND_1295[4:0];
  _RAND_1296 = {1{`RANDOM}};
  T_26182_11_pdst = _RAND_1296[6:0];
  _RAND_1297 = {1{`RANDOM}};
  T_26182_11_pop1 = _RAND_1297[6:0];
  _RAND_1298 = {1{`RANDOM}};
  T_26182_11_pop2 = _RAND_1298[6:0];
  _RAND_1299 = {1{`RANDOM}};
  T_26182_11_pop3 = _RAND_1299[6:0];
  _RAND_1300 = {1{`RANDOM}};
  T_26182_11_prs1_busy = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  T_26182_11_prs2_busy = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  T_26182_11_prs3_busy = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  T_26182_11_stale_pdst = _RAND_1303[6:0];
  _RAND_1304 = {1{`RANDOM}};
  T_26182_11_exception = _RAND_1304[0:0];
  _RAND_1305 = {2{`RANDOM}};
  T_26182_11_exc_cause = _RAND_1305[63:0];
  _RAND_1306 = {1{`RANDOM}};
  T_26182_11_bypassable = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  T_26182_11_mem_cmd = _RAND_1307[3:0];
  _RAND_1308 = {1{`RANDOM}};
  T_26182_11_mem_typ = _RAND_1308[2:0];
  _RAND_1309 = {1{`RANDOM}};
  T_26182_11_is_fence = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  T_26182_11_is_fencei = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  T_26182_11_is_store = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  T_26182_11_is_amo = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  T_26182_11_is_load = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  T_26182_11_is_unique = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  T_26182_11_flush_on_commit = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  T_26182_11_ldst = _RAND_1316[5:0];
  _RAND_1317 = {1{`RANDOM}};
  T_26182_11_lrs1 = _RAND_1317[5:0];
  _RAND_1318 = {1{`RANDOM}};
  T_26182_11_lrs2 = _RAND_1318[5:0];
  _RAND_1319 = {1{`RANDOM}};
  T_26182_11_lrs3 = _RAND_1319[5:0];
  _RAND_1320 = {1{`RANDOM}};
  T_26182_11_ldst_val = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  T_26182_11_dst_rtype = _RAND_1321[1:0];
  _RAND_1322 = {1{`RANDOM}};
  T_26182_11_lrs1_rtype = _RAND_1322[1:0];
  _RAND_1323 = {1{`RANDOM}};
  T_26182_11_lrs2_rtype = _RAND_1323[1:0];
  _RAND_1324 = {1{`RANDOM}};
  T_26182_11_frs3_en = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  T_26182_11_fp_val = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  T_26182_11_fp_single = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  T_26182_11_xcpt_if = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  T_26182_11_replay_if = _RAND_1328[0:0];
  _RAND_1329 = {2{`RANDOM}};
  T_26182_11_debug_wdata = _RAND_1329[63:0];
  _RAND_1330 = {1{`RANDOM}};
  T_26182_11_debug_events_fetch_seq = _RAND_1330[31:0];
  _RAND_1331 = {1{`RANDOM}};
  T_26182_12_valid = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  T_26182_12_iw_state = _RAND_1332[1:0];
  _RAND_1333 = {1{`RANDOM}};
  T_26182_12_uopc = _RAND_1333[8:0];
  _RAND_1334 = {1{`RANDOM}};
  T_26182_12_inst = _RAND_1334[31:0];
  _RAND_1335 = {2{`RANDOM}};
  T_26182_12_pc = _RAND_1335[39:0];
  _RAND_1336 = {1{`RANDOM}};
  T_26182_12_fu_code = _RAND_1336[7:0];
  _RAND_1337 = {1{`RANDOM}};
  T_26182_12_ctrl_br_type = _RAND_1337[3:0];
  _RAND_1338 = {1{`RANDOM}};
  T_26182_12_ctrl_op1_sel = _RAND_1338[1:0];
  _RAND_1339 = {1{`RANDOM}};
  T_26182_12_ctrl_op2_sel = _RAND_1339[2:0];
  _RAND_1340 = {1{`RANDOM}};
  T_26182_12_ctrl_imm_sel = _RAND_1340[2:0];
  _RAND_1341 = {1{`RANDOM}};
  T_26182_12_ctrl_op_fcn = _RAND_1341[3:0];
  _RAND_1342 = {1{`RANDOM}};
  T_26182_12_ctrl_fcn_dw = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  T_26182_12_ctrl_rf_wen = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  T_26182_12_ctrl_csr_cmd = _RAND_1344[2:0];
  _RAND_1345 = {1{`RANDOM}};
  T_26182_12_ctrl_is_load = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  T_26182_12_ctrl_is_sta = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  T_26182_12_ctrl_is_std = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  T_26182_12_wakeup_delay = _RAND_1348[1:0];
  _RAND_1349 = {1{`RANDOM}};
  T_26182_12_allocate_brtag = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  T_26182_12_is_br_or_jmp = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  T_26182_12_is_jump = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  T_26182_12_is_jal = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  T_26182_12_is_ret = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  T_26182_12_is_call = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  T_26182_12_br_mask = _RAND_1355[7:0];
  _RAND_1356 = {1{`RANDOM}};
  T_26182_12_br_tag = _RAND_1356[2:0];
  _RAND_1357 = {1{`RANDOM}};
  T_26182_12_br_prediction_bpd_predict_val = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  T_26182_12_br_prediction_bpd_predict_taken = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  T_26182_12_br_prediction_btb_hit = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  T_26182_12_br_prediction_btb_predicted = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  T_26182_12_br_prediction_is_br_or_jalr = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  T_26182_12_stat_brjmp_mispredicted = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  T_26182_12_stat_btb_made_pred = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  T_26182_12_stat_btb_mispredicted = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  T_26182_12_stat_bpd_made_pred = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  T_26182_12_stat_bpd_mispredicted = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  T_26182_12_fetch_pc_lob = _RAND_1367[2:0];
  _RAND_1368 = {1{`RANDOM}};
  T_26182_12_imm_packed = _RAND_1368[19:0];
  _RAND_1369 = {1{`RANDOM}};
  T_26182_12_csr_addr = _RAND_1369[11:0];
  _RAND_1370 = {1{`RANDOM}};
  T_26182_12_rob_idx = _RAND_1370[5:0];
  _RAND_1371 = {1{`RANDOM}};
  T_26182_12_ldq_idx = _RAND_1371[3:0];
  _RAND_1372 = {1{`RANDOM}};
  T_26182_12_stq_idx = _RAND_1372[3:0];
  _RAND_1373 = {1{`RANDOM}};
  T_26182_12_brob_idx = _RAND_1373[4:0];
  _RAND_1374 = {1{`RANDOM}};
  T_26182_12_pdst = _RAND_1374[6:0];
  _RAND_1375 = {1{`RANDOM}};
  T_26182_12_pop1 = _RAND_1375[6:0];
  _RAND_1376 = {1{`RANDOM}};
  T_26182_12_pop2 = _RAND_1376[6:0];
  _RAND_1377 = {1{`RANDOM}};
  T_26182_12_pop3 = _RAND_1377[6:0];
  _RAND_1378 = {1{`RANDOM}};
  T_26182_12_prs1_busy = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  T_26182_12_prs2_busy = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  T_26182_12_prs3_busy = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  T_26182_12_stale_pdst = _RAND_1381[6:0];
  _RAND_1382 = {1{`RANDOM}};
  T_26182_12_exception = _RAND_1382[0:0];
  _RAND_1383 = {2{`RANDOM}};
  T_26182_12_exc_cause = _RAND_1383[63:0];
  _RAND_1384 = {1{`RANDOM}};
  T_26182_12_bypassable = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  T_26182_12_mem_cmd = _RAND_1385[3:0];
  _RAND_1386 = {1{`RANDOM}};
  T_26182_12_mem_typ = _RAND_1386[2:0];
  _RAND_1387 = {1{`RANDOM}};
  T_26182_12_is_fence = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  T_26182_12_is_fencei = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  T_26182_12_is_store = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  T_26182_12_is_amo = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  T_26182_12_is_load = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  T_26182_12_is_unique = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  T_26182_12_flush_on_commit = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  T_26182_12_ldst = _RAND_1394[5:0];
  _RAND_1395 = {1{`RANDOM}};
  T_26182_12_lrs1 = _RAND_1395[5:0];
  _RAND_1396 = {1{`RANDOM}};
  T_26182_12_lrs2 = _RAND_1396[5:0];
  _RAND_1397 = {1{`RANDOM}};
  T_26182_12_lrs3 = _RAND_1397[5:0];
  _RAND_1398 = {1{`RANDOM}};
  T_26182_12_ldst_val = _RAND_1398[0:0];
  _RAND_1399 = {1{`RANDOM}};
  T_26182_12_dst_rtype = _RAND_1399[1:0];
  _RAND_1400 = {1{`RANDOM}};
  T_26182_12_lrs1_rtype = _RAND_1400[1:0];
  _RAND_1401 = {1{`RANDOM}};
  T_26182_12_lrs2_rtype = _RAND_1401[1:0];
  _RAND_1402 = {1{`RANDOM}};
  T_26182_12_frs3_en = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  T_26182_12_fp_val = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  T_26182_12_fp_single = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  T_26182_12_xcpt_if = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  T_26182_12_replay_if = _RAND_1406[0:0];
  _RAND_1407 = {2{`RANDOM}};
  T_26182_12_debug_wdata = _RAND_1407[63:0];
  _RAND_1408 = {1{`RANDOM}};
  T_26182_12_debug_events_fetch_seq = _RAND_1408[31:0];
  _RAND_1409 = {1{`RANDOM}};
  T_26182_13_valid = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  T_26182_13_iw_state = _RAND_1410[1:0];
  _RAND_1411 = {1{`RANDOM}};
  T_26182_13_uopc = _RAND_1411[8:0];
  _RAND_1412 = {1{`RANDOM}};
  T_26182_13_inst = _RAND_1412[31:0];
  _RAND_1413 = {2{`RANDOM}};
  T_26182_13_pc = _RAND_1413[39:0];
  _RAND_1414 = {1{`RANDOM}};
  T_26182_13_fu_code = _RAND_1414[7:0];
  _RAND_1415 = {1{`RANDOM}};
  T_26182_13_ctrl_br_type = _RAND_1415[3:0];
  _RAND_1416 = {1{`RANDOM}};
  T_26182_13_ctrl_op1_sel = _RAND_1416[1:0];
  _RAND_1417 = {1{`RANDOM}};
  T_26182_13_ctrl_op2_sel = _RAND_1417[2:0];
  _RAND_1418 = {1{`RANDOM}};
  T_26182_13_ctrl_imm_sel = _RAND_1418[2:0];
  _RAND_1419 = {1{`RANDOM}};
  T_26182_13_ctrl_op_fcn = _RAND_1419[3:0];
  _RAND_1420 = {1{`RANDOM}};
  T_26182_13_ctrl_fcn_dw = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  T_26182_13_ctrl_rf_wen = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  T_26182_13_ctrl_csr_cmd = _RAND_1422[2:0];
  _RAND_1423 = {1{`RANDOM}};
  T_26182_13_ctrl_is_load = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  T_26182_13_ctrl_is_sta = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  T_26182_13_ctrl_is_std = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  T_26182_13_wakeup_delay = _RAND_1426[1:0];
  _RAND_1427 = {1{`RANDOM}};
  T_26182_13_allocate_brtag = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  T_26182_13_is_br_or_jmp = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  T_26182_13_is_jump = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  T_26182_13_is_jal = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  T_26182_13_is_ret = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  T_26182_13_is_call = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  T_26182_13_br_mask = _RAND_1433[7:0];
  _RAND_1434 = {1{`RANDOM}};
  T_26182_13_br_tag = _RAND_1434[2:0];
  _RAND_1435 = {1{`RANDOM}};
  T_26182_13_br_prediction_bpd_predict_val = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  T_26182_13_br_prediction_bpd_predict_taken = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  T_26182_13_br_prediction_btb_hit = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  T_26182_13_br_prediction_btb_predicted = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  T_26182_13_br_prediction_is_br_or_jalr = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  T_26182_13_stat_brjmp_mispredicted = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  T_26182_13_stat_btb_made_pred = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  T_26182_13_stat_btb_mispredicted = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  T_26182_13_stat_bpd_made_pred = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  T_26182_13_stat_bpd_mispredicted = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  T_26182_13_fetch_pc_lob = _RAND_1445[2:0];
  _RAND_1446 = {1{`RANDOM}};
  T_26182_13_imm_packed = _RAND_1446[19:0];
  _RAND_1447 = {1{`RANDOM}};
  T_26182_13_csr_addr = _RAND_1447[11:0];
  _RAND_1448 = {1{`RANDOM}};
  T_26182_13_rob_idx = _RAND_1448[5:0];
  _RAND_1449 = {1{`RANDOM}};
  T_26182_13_ldq_idx = _RAND_1449[3:0];
  _RAND_1450 = {1{`RANDOM}};
  T_26182_13_stq_idx = _RAND_1450[3:0];
  _RAND_1451 = {1{`RANDOM}};
  T_26182_13_brob_idx = _RAND_1451[4:0];
  _RAND_1452 = {1{`RANDOM}};
  T_26182_13_pdst = _RAND_1452[6:0];
  _RAND_1453 = {1{`RANDOM}};
  T_26182_13_pop1 = _RAND_1453[6:0];
  _RAND_1454 = {1{`RANDOM}};
  T_26182_13_pop2 = _RAND_1454[6:0];
  _RAND_1455 = {1{`RANDOM}};
  T_26182_13_pop3 = _RAND_1455[6:0];
  _RAND_1456 = {1{`RANDOM}};
  T_26182_13_prs1_busy = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  T_26182_13_prs2_busy = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  T_26182_13_prs3_busy = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  T_26182_13_stale_pdst = _RAND_1459[6:0];
  _RAND_1460 = {1{`RANDOM}};
  T_26182_13_exception = _RAND_1460[0:0];
  _RAND_1461 = {2{`RANDOM}};
  T_26182_13_exc_cause = _RAND_1461[63:0];
  _RAND_1462 = {1{`RANDOM}};
  T_26182_13_bypassable = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  T_26182_13_mem_cmd = _RAND_1463[3:0];
  _RAND_1464 = {1{`RANDOM}};
  T_26182_13_mem_typ = _RAND_1464[2:0];
  _RAND_1465 = {1{`RANDOM}};
  T_26182_13_is_fence = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  T_26182_13_is_fencei = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  T_26182_13_is_store = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  T_26182_13_is_amo = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  T_26182_13_is_load = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  T_26182_13_is_unique = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  T_26182_13_flush_on_commit = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  T_26182_13_ldst = _RAND_1472[5:0];
  _RAND_1473 = {1{`RANDOM}};
  T_26182_13_lrs1 = _RAND_1473[5:0];
  _RAND_1474 = {1{`RANDOM}};
  T_26182_13_lrs2 = _RAND_1474[5:0];
  _RAND_1475 = {1{`RANDOM}};
  T_26182_13_lrs3 = _RAND_1475[5:0];
  _RAND_1476 = {1{`RANDOM}};
  T_26182_13_ldst_val = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  T_26182_13_dst_rtype = _RAND_1477[1:0];
  _RAND_1478 = {1{`RANDOM}};
  T_26182_13_lrs1_rtype = _RAND_1478[1:0];
  _RAND_1479 = {1{`RANDOM}};
  T_26182_13_lrs2_rtype = _RAND_1479[1:0];
  _RAND_1480 = {1{`RANDOM}};
  T_26182_13_frs3_en = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  T_26182_13_fp_val = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  T_26182_13_fp_single = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  T_26182_13_xcpt_if = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  T_26182_13_replay_if = _RAND_1484[0:0];
  _RAND_1485 = {2{`RANDOM}};
  T_26182_13_debug_wdata = _RAND_1485[63:0];
  _RAND_1486 = {1{`RANDOM}};
  T_26182_13_debug_events_fetch_seq = _RAND_1486[31:0];
  _RAND_1487 = {1{`RANDOM}};
  T_26182_14_valid = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  T_26182_14_iw_state = _RAND_1488[1:0];
  _RAND_1489 = {1{`RANDOM}};
  T_26182_14_uopc = _RAND_1489[8:0];
  _RAND_1490 = {1{`RANDOM}};
  T_26182_14_inst = _RAND_1490[31:0];
  _RAND_1491 = {2{`RANDOM}};
  T_26182_14_pc = _RAND_1491[39:0];
  _RAND_1492 = {1{`RANDOM}};
  T_26182_14_fu_code = _RAND_1492[7:0];
  _RAND_1493 = {1{`RANDOM}};
  T_26182_14_ctrl_br_type = _RAND_1493[3:0];
  _RAND_1494 = {1{`RANDOM}};
  T_26182_14_ctrl_op1_sel = _RAND_1494[1:0];
  _RAND_1495 = {1{`RANDOM}};
  T_26182_14_ctrl_op2_sel = _RAND_1495[2:0];
  _RAND_1496 = {1{`RANDOM}};
  T_26182_14_ctrl_imm_sel = _RAND_1496[2:0];
  _RAND_1497 = {1{`RANDOM}};
  T_26182_14_ctrl_op_fcn = _RAND_1497[3:0];
  _RAND_1498 = {1{`RANDOM}};
  T_26182_14_ctrl_fcn_dw = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  T_26182_14_ctrl_rf_wen = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  T_26182_14_ctrl_csr_cmd = _RAND_1500[2:0];
  _RAND_1501 = {1{`RANDOM}};
  T_26182_14_ctrl_is_load = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  T_26182_14_ctrl_is_sta = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  T_26182_14_ctrl_is_std = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  T_26182_14_wakeup_delay = _RAND_1504[1:0];
  _RAND_1505 = {1{`RANDOM}};
  T_26182_14_allocate_brtag = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  T_26182_14_is_br_or_jmp = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  T_26182_14_is_jump = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  T_26182_14_is_jal = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  T_26182_14_is_ret = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  T_26182_14_is_call = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  T_26182_14_br_mask = _RAND_1511[7:0];
  _RAND_1512 = {1{`RANDOM}};
  T_26182_14_br_tag = _RAND_1512[2:0];
  _RAND_1513 = {1{`RANDOM}};
  T_26182_14_br_prediction_bpd_predict_val = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  T_26182_14_br_prediction_bpd_predict_taken = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  T_26182_14_br_prediction_btb_hit = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  T_26182_14_br_prediction_btb_predicted = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  T_26182_14_br_prediction_is_br_or_jalr = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  T_26182_14_stat_brjmp_mispredicted = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  T_26182_14_stat_btb_made_pred = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  T_26182_14_stat_btb_mispredicted = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  T_26182_14_stat_bpd_made_pred = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  T_26182_14_stat_bpd_mispredicted = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  T_26182_14_fetch_pc_lob = _RAND_1523[2:0];
  _RAND_1524 = {1{`RANDOM}};
  T_26182_14_imm_packed = _RAND_1524[19:0];
  _RAND_1525 = {1{`RANDOM}};
  T_26182_14_csr_addr = _RAND_1525[11:0];
  _RAND_1526 = {1{`RANDOM}};
  T_26182_14_rob_idx = _RAND_1526[5:0];
  _RAND_1527 = {1{`RANDOM}};
  T_26182_14_ldq_idx = _RAND_1527[3:0];
  _RAND_1528 = {1{`RANDOM}};
  T_26182_14_stq_idx = _RAND_1528[3:0];
  _RAND_1529 = {1{`RANDOM}};
  T_26182_14_brob_idx = _RAND_1529[4:0];
  _RAND_1530 = {1{`RANDOM}};
  T_26182_14_pdst = _RAND_1530[6:0];
  _RAND_1531 = {1{`RANDOM}};
  T_26182_14_pop1 = _RAND_1531[6:0];
  _RAND_1532 = {1{`RANDOM}};
  T_26182_14_pop2 = _RAND_1532[6:0];
  _RAND_1533 = {1{`RANDOM}};
  T_26182_14_pop3 = _RAND_1533[6:0];
  _RAND_1534 = {1{`RANDOM}};
  T_26182_14_prs1_busy = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  T_26182_14_prs2_busy = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  T_26182_14_prs3_busy = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  T_26182_14_stale_pdst = _RAND_1537[6:0];
  _RAND_1538 = {1{`RANDOM}};
  T_26182_14_exception = _RAND_1538[0:0];
  _RAND_1539 = {2{`RANDOM}};
  T_26182_14_exc_cause = _RAND_1539[63:0];
  _RAND_1540 = {1{`RANDOM}};
  T_26182_14_bypassable = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  T_26182_14_mem_cmd = _RAND_1541[3:0];
  _RAND_1542 = {1{`RANDOM}};
  T_26182_14_mem_typ = _RAND_1542[2:0];
  _RAND_1543 = {1{`RANDOM}};
  T_26182_14_is_fence = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  T_26182_14_is_fencei = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  T_26182_14_is_store = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  T_26182_14_is_amo = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  T_26182_14_is_load = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  T_26182_14_is_unique = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  T_26182_14_flush_on_commit = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  T_26182_14_ldst = _RAND_1550[5:0];
  _RAND_1551 = {1{`RANDOM}};
  T_26182_14_lrs1 = _RAND_1551[5:0];
  _RAND_1552 = {1{`RANDOM}};
  T_26182_14_lrs2 = _RAND_1552[5:0];
  _RAND_1553 = {1{`RANDOM}};
  T_26182_14_lrs3 = _RAND_1553[5:0];
  _RAND_1554 = {1{`RANDOM}};
  T_26182_14_ldst_val = _RAND_1554[0:0];
  _RAND_1555 = {1{`RANDOM}};
  T_26182_14_dst_rtype = _RAND_1555[1:0];
  _RAND_1556 = {1{`RANDOM}};
  T_26182_14_lrs1_rtype = _RAND_1556[1:0];
  _RAND_1557 = {1{`RANDOM}};
  T_26182_14_lrs2_rtype = _RAND_1557[1:0];
  _RAND_1558 = {1{`RANDOM}};
  T_26182_14_frs3_en = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  T_26182_14_fp_val = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  T_26182_14_fp_single = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  T_26182_14_xcpt_if = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  T_26182_14_replay_if = _RAND_1562[0:0];
  _RAND_1563 = {2{`RANDOM}};
  T_26182_14_debug_wdata = _RAND_1563[63:0];
  _RAND_1564 = {1{`RANDOM}};
  T_26182_14_debug_events_fetch_seq = _RAND_1564[31:0];
  _RAND_1565 = {1{`RANDOM}};
  T_26182_15_valid = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  T_26182_15_iw_state = _RAND_1566[1:0];
  _RAND_1567 = {1{`RANDOM}};
  T_26182_15_uopc = _RAND_1567[8:0];
  _RAND_1568 = {1{`RANDOM}};
  T_26182_15_inst = _RAND_1568[31:0];
  _RAND_1569 = {2{`RANDOM}};
  T_26182_15_pc = _RAND_1569[39:0];
  _RAND_1570 = {1{`RANDOM}};
  T_26182_15_fu_code = _RAND_1570[7:0];
  _RAND_1571 = {1{`RANDOM}};
  T_26182_15_ctrl_br_type = _RAND_1571[3:0];
  _RAND_1572 = {1{`RANDOM}};
  T_26182_15_ctrl_op1_sel = _RAND_1572[1:0];
  _RAND_1573 = {1{`RANDOM}};
  T_26182_15_ctrl_op2_sel = _RAND_1573[2:0];
  _RAND_1574 = {1{`RANDOM}};
  T_26182_15_ctrl_imm_sel = _RAND_1574[2:0];
  _RAND_1575 = {1{`RANDOM}};
  T_26182_15_ctrl_op_fcn = _RAND_1575[3:0];
  _RAND_1576 = {1{`RANDOM}};
  T_26182_15_ctrl_fcn_dw = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  T_26182_15_ctrl_rf_wen = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  T_26182_15_ctrl_csr_cmd = _RAND_1578[2:0];
  _RAND_1579 = {1{`RANDOM}};
  T_26182_15_ctrl_is_load = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  T_26182_15_ctrl_is_sta = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  T_26182_15_ctrl_is_std = _RAND_1581[0:0];
  _RAND_1582 = {1{`RANDOM}};
  T_26182_15_wakeup_delay = _RAND_1582[1:0];
  _RAND_1583 = {1{`RANDOM}};
  T_26182_15_allocate_brtag = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  T_26182_15_is_br_or_jmp = _RAND_1584[0:0];
  _RAND_1585 = {1{`RANDOM}};
  T_26182_15_is_jump = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  T_26182_15_is_jal = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  T_26182_15_is_ret = _RAND_1587[0:0];
  _RAND_1588 = {1{`RANDOM}};
  T_26182_15_is_call = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  T_26182_15_br_mask = _RAND_1589[7:0];
  _RAND_1590 = {1{`RANDOM}};
  T_26182_15_br_tag = _RAND_1590[2:0];
  _RAND_1591 = {1{`RANDOM}};
  T_26182_15_br_prediction_bpd_predict_val = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  T_26182_15_br_prediction_bpd_predict_taken = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  T_26182_15_br_prediction_btb_hit = _RAND_1593[0:0];
  _RAND_1594 = {1{`RANDOM}};
  T_26182_15_br_prediction_btb_predicted = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  T_26182_15_br_prediction_is_br_or_jalr = _RAND_1595[0:0];
  _RAND_1596 = {1{`RANDOM}};
  T_26182_15_stat_brjmp_mispredicted = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  T_26182_15_stat_btb_made_pred = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  T_26182_15_stat_btb_mispredicted = _RAND_1598[0:0];
  _RAND_1599 = {1{`RANDOM}};
  T_26182_15_stat_bpd_made_pred = _RAND_1599[0:0];
  _RAND_1600 = {1{`RANDOM}};
  T_26182_15_stat_bpd_mispredicted = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  T_26182_15_fetch_pc_lob = _RAND_1601[2:0];
  _RAND_1602 = {1{`RANDOM}};
  T_26182_15_imm_packed = _RAND_1602[19:0];
  _RAND_1603 = {1{`RANDOM}};
  T_26182_15_csr_addr = _RAND_1603[11:0];
  _RAND_1604 = {1{`RANDOM}};
  T_26182_15_rob_idx = _RAND_1604[5:0];
  _RAND_1605 = {1{`RANDOM}};
  T_26182_15_ldq_idx = _RAND_1605[3:0];
  _RAND_1606 = {1{`RANDOM}};
  T_26182_15_stq_idx = _RAND_1606[3:0];
  _RAND_1607 = {1{`RANDOM}};
  T_26182_15_brob_idx = _RAND_1607[4:0];
  _RAND_1608 = {1{`RANDOM}};
  T_26182_15_pdst = _RAND_1608[6:0];
  _RAND_1609 = {1{`RANDOM}};
  T_26182_15_pop1 = _RAND_1609[6:0];
  _RAND_1610 = {1{`RANDOM}};
  T_26182_15_pop2 = _RAND_1610[6:0];
  _RAND_1611 = {1{`RANDOM}};
  T_26182_15_pop3 = _RAND_1611[6:0];
  _RAND_1612 = {1{`RANDOM}};
  T_26182_15_prs1_busy = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  T_26182_15_prs2_busy = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  T_26182_15_prs3_busy = _RAND_1614[0:0];
  _RAND_1615 = {1{`RANDOM}};
  T_26182_15_stale_pdst = _RAND_1615[6:0];
  _RAND_1616 = {1{`RANDOM}};
  T_26182_15_exception = _RAND_1616[0:0];
  _RAND_1617 = {2{`RANDOM}};
  T_26182_15_exc_cause = _RAND_1617[63:0];
  _RAND_1618 = {1{`RANDOM}};
  T_26182_15_bypassable = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  T_26182_15_mem_cmd = _RAND_1619[3:0];
  _RAND_1620 = {1{`RANDOM}};
  T_26182_15_mem_typ = _RAND_1620[2:0];
  _RAND_1621 = {1{`RANDOM}};
  T_26182_15_is_fence = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  T_26182_15_is_fencei = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  T_26182_15_is_store = _RAND_1623[0:0];
  _RAND_1624 = {1{`RANDOM}};
  T_26182_15_is_amo = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  T_26182_15_is_load = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  T_26182_15_is_unique = _RAND_1626[0:0];
  _RAND_1627 = {1{`RANDOM}};
  T_26182_15_flush_on_commit = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  T_26182_15_ldst = _RAND_1628[5:0];
  _RAND_1629 = {1{`RANDOM}};
  T_26182_15_lrs1 = _RAND_1629[5:0];
  _RAND_1630 = {1{`RANDOM}};
  T_26182_15_lrs2 = _RAND_1630[5:0];
  _RAND_1631 = {1{`RANDOM}};
  T_26182_15_lrs3 = _RAND_1631[5:0];
  _RAND_1632 = {1{`RANDOM}};
  T_26182_15_ldst_val = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  T_26182_15_dst_rtype = _RAND_1633[1:0];
  _RAND_1634 = {1{`RANDOM}};
  T_26182_15_lrs1_rtype = _RAND_1634[1:0];
  _RAND_1635 = {1{`RANDOM}};
  T_26182_15_lrs2_rtype = _RAND_1635[1:0];
  _RAND_1636 = {1{`RANDOM}};
  T_26182_15_frs3_en = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  T_26182_15_fp_val = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  T_26182_15_fp_single = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  T_26182_15_xcpt_if = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  T_26182_15_replay_if = _RAND_1640[0:0];
  _RAND_1641 = {2{`RANDOM}};
  T_26182_15_debug_wdata = _RAND_1641[63:0];
  _RAND_1642 = {1{`RANDOM}};
  T_26182_15_debug_events_fetch_seq = _RAND_1642[31:0];
  _RAND_1643 = {1{`RANDOM}};
  T_26182_16_valid = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  T_26182_16_iw_state = _RAND_1644[1:0];
  _RAND_1645 = {1{`RANDOM}};
  T_26182_16_uopc = _RAND_1645[8:0];
  _RAND_1646 = {1{`RANDOM}};
  T_26182_16_inst = _RAND_1646[31:0];
  _RAND_1647 = {2{`RANDOM}};
  T_26182_16_pc = _RAND_1647[39:0];
  _RAND_1648 = {1{`RANDOM}};
  T_26182_16_fu_code = _RAND_1648[7:0];
  _RAND_1649 = {1{`RANDOM}};
  T_26182_16_ctrl_br_type = _RAND_1649[3:0];
  _RAND_1650 = {1{`RANDOM}};
  T_26182_16_ctrl_op1_sel = _RAND_1650[1:0];
  _RAND_1651 = {1{`RANDOM}};
  T_26182_16_ctrl_op2_sel = _RAND_1651[2:0];
  _RAND_1652 = {1{`RANDOM}};
  T_26182_16_ctrl_imm_sel = _RAND_1652[2:0];
  _RAND_1653 = {1{`RANDOM}};
  T_26182_16_ctrl_op_fcn = _RAND_1653[3:0];
  _RAND_1654 = {1{`RANDOM}};
  T_26182_16_ctrl_fcn_dw = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  T_26182_16_ctrl_rf_wen = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  T_26182_16_ctrl_csr_cmd = _RAND_1656[2:0];
  _RAND_1657 = {1{`RANDOM}};
  T_26182_16_ctrl_is_load = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  T_26182_16_ctrl_is_sta = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  T_26182_16_ctrl_is_std = _RAND_1659[0:0];
  _RAND_1660 = {1{`RANDOM}};
  T_26182_16_wakeup_delay = _RAND_1660[1:0];
  _RAND_1661 = {1{`RANDOM}};
  T_26182_16_allocate_brtag = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  T_26182_16_is_br_or_jmp = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  T_26182_16_is_jump = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  T_26182_16_is_jal = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  T_26182_16_is_ret = _RAND_1665[0:0];
  _RAND_1666 = {1{`RANDOM}};
  T_26182_16_is_call = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  T_26182_16_br_mask = _RAND_1667[7:0];
  _RAND_1668 = {1{`RANDOM}};
  T_26182_16_br_tag = _RAND_1668[2:0];
  _RAND_1669 = {1{`RANDOM}};
  T_26182_16_br_prediction_bpd_predict_val = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  T_26182_16_br_prediction_bpd_predict_taken = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  T_26182_16_br_prediction_btb_hit = _RAND_1671[0:0];
  _RAND_1672 = {1{`RANDOM}};
  T_26182_16_br_prediction_btb_predicted = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  T_26182_16_br_prediction_is_br_or_jalr = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  T_26182_16_stat_brjmp_mispredicted = _RAND_1674[0:0];
  _RAND_1675 = {1{`RANDOM}};
  T_26182_16_stat_btb_made_pred = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  T_26182_16_stat_btb_mispredicted = _RAND_1676[0:0];
  _RAND_1677 = {1{`RANDOM}};
  T_26182_16_stat_bpd_made_pred = _RAND_1677[0:0];
  _RAND_1678 = {1{`RANDOM}};
  T_26182_16_stat_bpd_mispredicted = _RAND_1678[0:0];
  _RAND_1679 = {1{`RANDOM}};
  T_26182_16_fetch_pc_lob = _RAND_1679[2:0];
  _RAND_1680 = {1{`RANDOM}};
  T_26182_16_imm_packed = _RAND_1680[19:0];
  _RAND_1681 = {1{`RANDOM}};
  T_26182_16_csr_addr = _RAND_1681[11:0];
  _RAND_1682 = {1{`RANDOM}};
  T_26182_16_rob_idx = _RAND_1682[5:0];
  _RAND_1683 = {1{`RANDOM}};
  T_26182_16_ldq_idx = _RAND_1683[3:0];
  _RAND_1684 = {1{`RANDOM}};
  T_26182_16_stq_idx = _RAND_1684[3:0];
  _RAND_1685 = {1{`RANDOM}};
  T_26182_16_brob_idx = _RAND_1685[4:0];
  _RAND_1686 = {1{`RANDOM}};
  T_26182_16_pdst = _RAND_1686[6:0];
  _RAND_1687 = {1{`RANDOM}};
  T_26182_16_pop1 = _RAND_1687[6:0];
  _RAND_1688 = {1{`RANDOM}};
  T_26182_16_pop2 = _RAND_1688[6:0];
  _RAND_1689 = {1{`RANDOM}};
  T_26182_16_pop3 = _RAND_1689[6:0];
  _RAND_1690 = {1{`RANDOM}};
  T_26182_16_prs1_busy = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  T_26182_16_prs2_busy = _RAND_1691[0:0];
  _RAND_1692 = {1{`RANDOM}};
  T_26182_16_prs3_busy = _RAND_1692[0:0];
  _RAND_1693 = {1{`RANDOM}};
  T_26182_16_stale_pdst = _RAND_1693[6:0];
  _RAND_1694 = {1{`RANDOM}};
  T_26182_16_exception = _RAND_1694[0:0];
  _RAND_1695 = {2{`RANDOM}};
  T_26182_16_exc_cause = _RAND_1695[63:0];
  _RAND_1696 = {1{`RANDOM}};
  T_26182_16_bypassable = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  T_26182_16_mem_cmd = _RAND_1697[3:0];
  _RAND_1698 = {1{`RANDOM}};
  T_26182_16_mem_typ = _RAND_1698[2:0];
  _RAND_1699 = {1{`RANDOM}};
  T_26182_16_is_fence = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  T_26182_16_is_fencei = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  T_26182_16_is_store = _RAND_1701[0:0];
  _RAND_1702 = {1{`RANDOM}};
  T_26182_16_is_amo = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  T_26182_16_is_load = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  T_26182_16_is_unique = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  T_26182_16_flush_on_commit = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  T_26182_16_ldst = _RAND_1706[5:0];
  _RAND_1707 = {1{`RANDOM}};
  T_26182_16_lrs1 = _RAND_1707[5:0];
  _RAND_1708 = {1{`RANDOM}};
  T_26182_16_lrs2 = _RAND_1708[5:0];
  _RAND_1709 = {1{`RANDOM}};
  T_26182_16_lrs3 = _RAND_1709[5:0];
  _RAND_1710 = {1{`RANDOM}};
  T_26182_16_ldst_val = _RAND_1710[0:0];
  _RAND_1711 = {1{`RANDOM}};
  T_26182_16_dst_rtype = _RAND_1711[1:0];
  _RAND_1712 = {1{`RANDOM}};
  T_26182_16_lrs1_rtype = _RAND_1712[1:0];
  _RAND_1713 = {1{`RANDOM}};
  T_26182_16_lrs2_rtype = _RAND_1713[1:0];
  _RAND_1714 = {1{`RANDOM}};
  T_26182_16_frs3_en = _RAND_1714[0:0];
  _RAND_1715 = {1{`RANDOM}};
  T_26182_16_fp_val = _RAND_1715[0:0];
  _RAND_1716 = {1{`RANDOM}};
  T_26182_16_fp_single = _RAND_1716[0:0];
  _RAND_1717 = {1{`RANDOM}};
  T_26182_16_xcpt_if = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  T_26182_16_replay_if = _RAND_1718[0:0];
  _RAND_1719 = {2{`RANDOM}};
  T_26182_16_debug_wdata = _RAND_1719[63:0];
  _RAND_1720 = {1{`RANDOM}};
  T_26182_16_debug_events_fetch_seq = _RAND_1720[31:0];
  _RAND_1721 = {1{`RANDOM}};
  T_26182_17_valid = _RAND_1721[0:0];
  _RAND_1722 = {1{`RANDOM}};
  T_26182_17_iw_state = _RAND_1722[1:0];
  _RAND_1723 = {1{`RANDOM}};
  T_26182_17_uopc = _RAND_1723[8:0];
  _RAND_1724 = {1{`RANDOM}};
  T_26182_17_inst = _RAND_1724[31:0];
  _RAND_1725 = {2{`RANDOM}};
  T_26182_17_pc = _RAND_1725[39:0];
  _RAND_1726 = {1{`RANDOM}};
  T_26182_17_fu_code = _RAND_1726[7:0];
  _RAND_1727 = {1{`RANDOM}};
  T_26182_17_ctrl_br_type = _RAND_1727[3:0];
  _RAND_1728 = {1{`RANDOM}};
  T_26182_17_ctrl_op1_sel = _RAND_1728[1:0];
  _RAND_1729 = {1{`RANDOM}};
  T_26182_17_ctrl_op2_sel = _RAND_1729[2:0];
  _RAND_1730 = {1{`RANDOM}};
  T_26182_17_ctrl_imm_sel = _RAND_1730[2:0];
  _RAND_1731 = {1{`RANDOM}};
  T_26182_17_ctrl_op_fcn = _RAND_1731[3:0];
  _RAND_1732 = {1{`RANDOM}};
  T_26182_17_ctrl_fcn_dw = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  T_26182_17_ctrl_rf_wen = _RAND_1733[0:0];
  _RAND_1734 = {1{`RANDOM}};
  T_26182_17_ctrl_csr_cmd = _RAND_1734[2:0];
  _RAND_1735 = {1{`RANDOM}};
  T_26182_17_ctrl_is_load = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  T_26182_17_ctrl_is_sta = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  T_26182_17_ctrl_is_std = _RAND_1737[0:0];
  _RAND_1738 = {1{`RANDOM}};
  T_26182_17_wakeup_delay = _RAND_1738[1:0];
  _RAND_1739 = {1{`RANDOM}};
  T_26182_17_allocate_brtag = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  T_26182_17_is_br_or_jmp = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  T_26182_17_is_jump = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  T_26182_17_is_jal = _RAND_1742[0:0];
  _RAND_1743 = {1{`RANDOM}};
  T_26182_17_is_ret = _RAND_1743[0:0];
  _RAND_1744 = {1{`RANDOM}};
  T_26182_17_is_call = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  T_26182_17_br_mask = _RAND_1745[7:0];
  _RAND_1746 = {1{`RANDOM}};
  T_26182_17_br_tag = _RAND_1746[2:0];
  _RAND_1747 = {1{`RANDOM}};
  T_26182_17_br_prediction_bpd_predict_val = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  T_26182_17_br_prediction_bpd_predict_taken = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  T_26182_17_br_prediction_btb_hit = _RAND_1749[0:0];
  _RAND_1750 = {1{`RANDOM}};
  T_26182_17_br_prediction_btb_predicted = _RAND_1750[0:0];
  _RAND_1751 = {1{`RANDOM}};
  T_26182_17_br_prediction_is_br_or_jalr = _RAND_1751[0:0];
  _RAND_1752 = {1{`RANDOM}};
  T_26182_17_stat_brjmp_mispredicted = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  T_26182_17_stat_btb_made_pred = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  T_26182_17_stat_btb_mispredicted = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  T_26182_17_stat_bpd_made_pred = _RAND_1755[0:0];
  _RAND_1756 = {1{`RANDOM}};
  T_26182_17_stat_bpd_mispredicted = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  T_26182_17_fetch_pc_lob = _RAND_1757[2:0];
  _RAND_1758 = {1{`RANDOM}};
  T_26182_17_imm_packed = _RAND_1758[19:0];
  _RAND_1759 = {1{`RANDOM}};
  T_26182_17_csr_addr = _RAND_1759[11:0];
  _RAND_1760 = {1{`RANDOM}};
  T_26182_17_rob_idx = _RAND_1760[5:0];
  _RAND_1761 = {1{`RANDOM}};
  T_26182_17_ldq_idx = _RAND_1761[3:0];
  _RAND_1762 = {1{`RANDOM}};
  T_26182_17_stq_idx = _RAND_1762[3:0];
  _RAND_1763 = {1{`RANDOM}};
  T_26182_17_brob_idx = _RAND_1763[4:0];
  _RAND_1764 = {1{`RANDOM}};
  T_26182_17_pdst = _RAND_1764[6:0];
  _RAND_1765 = {1{`RANDOM}};
  T_26182_17_pop1 = _RAND_1765[6:0];
  _RAND_1766 = {1{`RANDOM}};
  T_26182_17_pop2 = _RAND_1766[6:0];
  _RAND_1767 = {1{`RANDOM}};
  T_26182_17_pop3 = _RAND_1767[6:0];
  _RAND_1768 = {1{`RANDOM}};
  T_26182_17_prs1_busy = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  T_26182_17_prs2_busy = _RAND_1769[0:0];
  _RAND_1770 = {1{`RANDOM}};
  T_26182_17_prs3_busy = _RAND_1770[0:0];
  _RAND_1771 = {1{`RANDOM}};
  T_26182_17_stale_pdst = _RAND_1771[6:0];
  _RAND_1772 = {1{`RANDOM}};
  T_26182_17_exception = _RAND_1772[0:0];
  _RAND_1773 = {2{`RANDOM}};
  T_26182_17_exc_cause = _RAND_1773[63:0];
  _RAND_1774 = {1{`RANDOM}};
  T_26182_17_bypassable = _RAND_1774[0:0];
  _RAND_1775 = {1{`RANDOM}};
  T_26182_17_mem_cmd = _RAND_1775[3:0];
  _RAND_1776 = {1{`RANDOM}};
  T_26182_17_mem_typ = _RAND_1776[2:0];
  _RAND_1777 = {1{`RANDOM}};
  T_26182_17_is_fence = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  T_26182_17_is_fencei = _RAND_1778[0:0];
  _RAND_1779 = {1{`RANDOM}};
  T_26182_17_is_store = _RAND_1779[0:0];
  _RAND_1780 = {1{`RANDOM}};
  T_26182_17_is_amo = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  T_26182_17_is_load = _RAND_1781[0:0];
  _RAND_1782 = {1{`RANDOM}};
  T_26182_17_is_unique = _RAND_1782[0:0];
  _RAND_1783 = {1{`RANDOM}};
  T_26182_17_flush_on_commit = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  T_26182_17_ldst = _RAND_1784[5:0];
  _RAND_1785 = {1{`RANDOM}};
  T_26182_17_lrs1 = _RAND_1785[5:0];
  _RAND_1786 = {1{`RANDOM}};
  T_26182_17_lrs2 = _RAND_1786[5:0];
  _RAND_1787 = {1{`RANDOM}};
  T_26182_17_lrs3 = _RAND_1787[5:0];
  _RAND_1788 = {1{`RANDOM}};
  T_26182_17_ldst_val = _RAND_1788[0:0];
  _RAND_1789 = {1{`RANDOM}};
  T_26182_17_dst_rtype = _RAND_1789[1:0];
  _RAND_1790 = {1{`RANDOM}};
  T_26182_17_lrs1_rtype = _RAND_1790[1:0];
  _RAND_1791 = {1{`RANDOM}};
  T_26182_17_lrs2_rtype = _RAND_1791[1:0];
  _RAND_1792 = {1{`RANDOM}};
  T_26182_17_frs3_en = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  T_26182_17_fp_val = _RAND_1793[0:0];
  _RAND_1794 = {1{`RANDOM}};
  T_26182_17_fp_single = _RAND_1794[0:0];
  _RAND_1795 = {1{`RANDOM}};
  T_26182_17_xcpt_if = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  T_26182_17_replay_if = _RAND_1796[0:0];
  _RAND_1797 = {2{`RANDOM}};
  T_26182_17_debug_wdata = _RAND_1797[63:0];
  _RAND_1798 = {1{`RANDOM}};
  T_26182_17_debug_events_fetch_seq = _RAND_1798[31:0];
  _RAND_1799 = {1{`RANDOM}};
  T_26182_18_valid = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  T_26182_18_iw_state = _RAND_1800[1:0];
  _RAND_1801 = {1{`RANDOM}};
  T_26182_18_uopc = _RAND_1801[8:0];
  _RAND_1802 = {1{`RANDOM}};
  T_26182_18_inst = _RAND_1802[31:0];
  _RAND_1803 = {2{`RANDOM}};
  T_26182_18_pc = _RAND_1803[39:0];
  _RAND_1804 = {1{`RANDOM}};
  T_26182_18_fu_code = _RAND_1804[7:0];
  _RAND_1805 = {1{`RANDOM}};
  T_26182_18_ctrl_br_type = _RAND_1805[3:0];
  _RAND_1806 = {1{`RANDOM}};
  T_26182_18_ctrl_op1_sel = _RAND_1806[1:0];
  _RAND_1807 = {1{`RANDOM}};
  T_26182_18_ctrl_op2_sel = _RAND_1807[2:0];
  _RAND_1808 = {1{`RANDOM}};
  T_26182_18_ctrl_imm_sel = _RAND_1808[2:0];
  _RAND_1809 = {1{`RANDOM}};
  T_26182_18_ctrl_op_fcn = _RAND_1809[3:0];
  _RAND_1810 = {1{`RANDOM}};
  T_26182_18_ctrl_fcn_dw = _RAND_1810[0:0];
  _RAND_1811 = {1{`RANDOM}};
  T_26182_18_ctrl_rf_wen = _RAND_1811[0:0];
  _RAND_1812 = {1{`RANDOM}};
  T_26182_18_ctrl_csr_cmd = _RAND_1812[2:0];
  _RAND_1813 = {1{`RANDOM}};
  T_26182_18_ctrl_is_load = _RAND_1813[0:0];
  _RAND_1814 = {1{`RANDOM}};
  T_26182_18_ctrl_is_sta = _RAND_1814[0:0];
  _RAND_1815 = {1{`RANDOM}};
  T_26182_18_ctrl_is_std = _RAND_1815[0:0];
  _RAND_1816 = {1{`RANDOM}};
  T_26182_18_wakeup_delay = _RAND_1816[1:0];
  _RAND_1817 = {1{`RANDOM}};
  T_26182_18_allocate_brtag = _RAND_1817[0:0];
  _RAND_1818 = {1{`RANDOM}};
  T_26182_18_is_br_or_jmp = _RAND_1818[0:0];
  _RAND_1819 = {1{`RANDOM}};
  T_26182_18_is_jump = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  T_26182_18_is_jal = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  T_26182_18_is_ret = _RAND_1821[0:0];
  _RAND_1822 = {1{`RANDOM}};
  T_26182_18_is_call = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  T_26182_18_br_mask = _RAND_1823[7:0];
  _RAND_1824 = {1{`RANDOM}};
  T_26182_18_br_tag = _RAND_1824[2:0];
  _RAND_1825 = {1{`RANDOM}};
  T_26182_18_br_prediction_bpd_predict_val = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  T_26182_18_br_prediction_bpd_predict_taken = _RAND_1826[0:0];
  _RAND_1827 = {1{`RANDOM}};
  T_26182_18_br_prediction_btb_hit = _RAND_1827[0:0];
  _RAND_1828 = {1{`RANDOM}};
  T_26182_18_br_prediction_btb_predicted = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  T_26182_18_br_prediction_is_br_or_jalr = _RAND_1829[0:0];
  _RAND_1830 = {1{`RANDOM}};
  T_26182_18_stat_brjmp_mispredicted = _RAND_1830[0:0];
  _RAND_1831 = {1{`RANDOM}};
  T_26182_18_stat_btb_made_pred = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  T_26182_18_stat_btb_mispredicted = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  T_26182_18_stat_bpd_made_pred = _RAND_1833[0:0];
  _RAND_1834 = {1{`RANDOM}};
  T_26182_18_stat_bpd_mispredicted = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  T_26182_18_fetch_pc_lob = _RAND_1835[2:0];
  _RAND_1836 = {1{`RANDOM}};
  T_26182_18_imm_packed = _RAND_1836[19:0];
  _RAND_1837 = {1{`RANDOM}};
  T_26182_18_csr_addr = _RAND_1837[11:0];
  _RAND_1838 = {1{`RANDOM}};
  T_26182_18_rob_idx = _RAND_1838[5:0];
  _RAND_1839 = {1{`RANDOM}};
  T_26182_18_ldq_idx = _RAND_1839[3:0];
  _RAND_1840 = {1{`RANDOM}};
  T_26182_18_stq_idx = _RAND_1840[3:0];
  _RAND_1841 = {1{`RANDOM}};
  T_26182_18_brob_idx = _RAND_1841[4:0];
  _RAND_1842 = {1{`RANDOM}};
  T_26182_18_pdst = _RAND_1842[6:0];
  _RAND_1843 = {1{`RANDOM}};
  T_26182_18_pop1 = _RAND_1843[6:0];
  _RAND_1844 = {1{`RANDOM}};
  T_26182_18_pop2 = _RAND_1844[6:0];
  _RAND_1845 = {1{`RANDOM}};
  T_26182_18_pop3 = _RAND_1845[6:0];
  _RAND_1846 = {1{`RANDOM}};
  T_26182_18_prs1_busy = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  T_26182_18_prs2_busy = _RAND_1847[0:0];
  _RAND_1848 = {1{`RANDOM}};
  T_26182_18_prs3_busy = _RAND_1848[0:0];
  _RAND_1849 = {1{`RANDOM}};
  T_26182_18_stale_pdst = _RAND_1849[6:0];
  _RAND_1850 = {1{`RANDOM}};
  T_26182_18_exception = _RAND_1850[0:0];
  _RAND_1851 = {2{`RANDOM}};
  T_26182_18_exc_cause = _RAND_1851[63:0];
  _RAND_1852 = {1{`RANDOM}};
  T_26182_18_bypassable = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  T_26182_18_mem_cmd = _RAND_1853[3:0];
  _RAND_1854 = {1{`RANDOM}};
  T_26182_18_mem_typ = _RAND_1854[2:0];
  _RAND_1855 = {1{`RANDOM}};
  T_26182_18_is_fence = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  T_26182_18_is_fencei = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  T_26182_18_is_store = _RAND_1857[0:0];
  _RAND_1858 = {1{`RANDOM}};
  T_26182_18_is_amo = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  T_26182_18_is_load = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  T_26182_18_is_unique = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  T_26182_18_flush_on_commit = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  T_26182_18_ldst = _RAND_1862[5:0];
  _RAND_1863 = {1{`RANDOM}};
  T_26182_18_lrs1 = _RAND_1863[5:0];
  _RAND_1864 = {1{`RANDOM}};
  T_26182_18_lrs2 = _RAND_1864[5:0];
  _RAND_1865 = {1{`RANDOM}};
  T_26182_18_lrs3 = _RAND_1865[5:0];
  _RAND_1866 = {1{`RANDOM}};
  T_26182_18_ldst_val = _RAND_1866[0:0];
  _RAND_1867 = {1{`RANDOM}};
  T_26182_18_dst_rtype = _RAND_1867[1:0];
  _RAND_1868 = {1{`RANDOM}};
  T_26182_18_lrs1_rtype = _RAND_1868[1:0];
  _RAND_1869 = {1{`RANDOM}};
  T_26182_18_lrs2_rtype = _RAND_1869[1:0];
  _RAND_1870 = {1{`RANDOM}};
  T_26182_18_frs3_en = _RAND_1870[0:0];
  _RAND_1871 = {1{`RANDOM}};
  T_26182_18_fp_val = _RAND_1871[0:0];
  _RAND_1872 = {1{`RANDOM}};
  T_26182_18_fp_single = _RAND_1872[0:0];
  _RAND_1873 = {1{`RANDOM}};
  T_26182_18_xcpt_if = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  T_26182_18_replay_if = _RAND_1874[0:0];
  _RAND_1875 = {2{`RANDOM}};
  T_26182_18_debug_wdata = _RAND_1875[63:0];
  _RAND_1876 = {1{`RANDOM}};
  T_26182_18_debug_events_fetch_seq = _RAND_1876[31:0];
  _RAND_1877 = {1{`RANDOM}};
  T_26182_19_valid = _RAND_1877[0:0];
  _RAND_1878 = {1{`RANDOM}};
  T_26182_19_iw_state = _RAND_1878[1:0];
  _RAND_1879 = {1{`RANDOM}};
  T_26182_19_uopc = _RAND_1879[8:0];
  _RAND_1880 = {1{`RANDOM}};
  T_26182_19_inst = _RAND_1880[31:0];
  _RAND_1881 = {2{`RANDOM}};
  T_26182_19_pc = _RAND_1881[39:0];
  _RAND_1882 = {1{`RANDOM}};
  T_26182_19_fu_code = _RAND_1882[7:0];
  _RAND_1883 = {1{`RANDOM}};
  T_26182_19_ctrl_br_type = _RAND_1883[3:0];
  _RAND_1884 = {1{`RANDOM}};
  T_26182_19_ctrl_op1_sel = _RAND_1884[1:0];
  _RAND_1885 = {1{`RANDOM}};
  T_26182_19_ctrl_op2_sel = _RAND_1885[2:0];
  _RAND_1886 = {1{`RANDOM}};
  T_26182_19_ctrl_imm_sel = _RAND_1886[2:0];
  _RAND_1887 = {1{`RANDOM}};
  T_26182_19_ctrl_op_fcn = _RAND_1887[3:0];
  _RAND_1888 = {1{`RANDOM}};
  T_26182_19_ctrl_fcn_dw = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  T_26182_19_ctrl_rf_wen = _RAND_1889[0:0];
  _RAND_1890 = {1{`RANDOM}};
  T_26182_19_ctrl_csr_cmd = _RAND_1890[2:0];
  _RAND_1891 = {1{`RANDOM}};
  T_26182_19_ctrl_is_load = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  T_26182_19_ctrl_is_sta = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  T_26182_19_ctrl_is_std = _RAND_1893[0:0];
  _RAND_1894 = {1{`RANDOM}};
  T_26182_19_wakeup_delay = _RAND_1894[1:0];
  _RAND_1895 = {1{`RANDOM}};
  T_26182_19_allocate_brtag = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  T_26182_19_is_br_or_jmp = _RAND_1896[0:0];
  _RAND_1897 = {1{`RANDOM}};
  T_26182_19_is_jump = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  T_26182_19_is_jal = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  T_26182_19_is_ret = _RAND_1899[0:0];
  _RAND_1900 = {1{`RANDOM}};
  T_26182_19_is_call = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  T_26182_19_br_mask = _RAND_1901[7:0];
  _RAND_1902 = {1{`RANDOM}};
  T_26182_19_br_tag = _RAND_1902[2:0];
  _RAND_1903 = {1{`RANDOM}};
  T_26182_19_br_prediction_bpd_predict_val = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  T_26182_19_br_prediction_bpd_predict_taken = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  T_26182_19_br_prediction_btb_hit = _RAND_1905[0:0];
  _RAND_1906 = {1{`RANDOM}};
  T_26182_19_br_prediction_btb_predicted = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  T_26182_19_br_prediction_is_br_or_jalr = _RAND_1907[0:0];
  _RAND_1908 = {1{`RANDOM}};
  T_26182_19_stat_brjmp_mispredicted = _RAND_1908[0:0];
  _RAND_1909 = {1{`RANDOM}};
  T_26182_19_stat_btb_made_pred = _RAND_1909[0:0];
  _RAND_1910 = {1{`RANDOM}};
  T_26182_19_stat_btb_mispredicted = _RAND_1910[0:0];
  _RAND_1911 = {1{`RANDOM}};
  T_26182_19_stat_bpd_made_pred = _RAND_1911[0:0];
  _RAND_1912 = {1{`RANDOM}};
  T_26182_19_stat_bpd_mispredicted = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  T_26182_19_fetch_pc_lob = _RAND_1913[2:0];
  _RAND_1914 = {1{`RANDOM}};
  T_26182_19_imm_packed = _RAND_1914[19:0];
  _RAND_1915 = {1{`RANDOM}};
  T_26182_19_csr_addr = _RAND_1915[11:0];
  _RAND_1916 = {1{`RANDOM}};
  T_26182_19_rob_idx = _RAND_1916[5:0];
  _RAND_1917 = {1{`RANDOM}};
  T_26182_19_ldq_idx = _RAND_1917[3:0];
  _RAND_1918 = {1{`RANDOM}};
  T_26182_19_stq_idx = _RAND_1918[3:0];
  _RAND_1919 = {1{`RANDOM}};
  T_26182_19_brob_idx = _RAND_1919[4:0];
  _RAND_1920 = {1{`RANDOM}};
  T_26182_19_pdst = _RAND_1920[6:0];
  _RAND_1921 = {1{`RANDOM}};
  T_26182_19_pop1 = _RAND_1921[6:0];
  _RAND_1922 = {1{`RANDOM}};
  T_26182_19_pop2 = _RAND_1922[6:0];
  _RAND_1923 = {1{`RANDOM}};
  T_26182_19_pop3 = _RAND_1923[6:0];
  _RAND_1924 = {1{`RANDOM}};
  T_26182_19_prs1_busy = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  T_26182_19_prs2_busy = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  T_26182_19_prs3_busy = _RAND_1926[0:0];
  _RAND_1927 = {1{`RANDOM}};
  T_26182_19_stale_pdst = _RAND_1927[6:0];
  _RAND_1928 = {1{`RANDOM}};
  T_26182_19_exception = _RAND_1928[0:0];
  _RAND_1929 = {2{`RANDOM}};
  T_26182_19_exc_cause = _RAND_1929[63:0];
  _RAND_1930 = {1{`RANDOM}};
  T_26182_19_bypassable = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  T_26182_19_mem_cmd = _RAND_1931[3:0];
  _RAND_1932 = {1{`RANDOM}};
  T_26182_19_mem_typ = _RAND_1932[2:0];
  _RAND_1933 = {1{`RANDOM}};
  T_26182_19_is_fence = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  T_26182_19_is_fencei = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  T_26182_19_is_store = _RAND_1935[0:0];
  _RAND_1936 = {1{`RANDOM}};
  T_26182_19_is_amo = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  T_26182_19_is_load = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  T_26182_19_is_unique = _RAND_1938[0:0];
  _RAND_1939 = {1{`RANDOM}};
  T_26182_19_flush_on_commit = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  T_26182_19_ldst = _RAND_1940[5:0];
  _RAND_1941 = {1{`RANDOM}};
  T_26182_19_lrs1 = _RAND_1941[5:0];
  _RAND_1942 = {1{`RANDOM}};
  T_26182_19_lrs2 = _RAND_1942[5:0];
  _RAND_1943 = {1{`RANDOM}};
  T_26182_19_lrs3 = _RAND_1943[5:0];
  _RAND_1944 = {1{`RANDOM}};
  T_26182_19_ldst_val = _RAND_1944[0:0];
  _RAND_1945 = {1{`RANDOM}};
  T_26182_19_dst_rtype = _RAND_1945[1:0];
  _RAND_1946 = {1{`RANDOM}};
  T_26182_19_lrs1_rtype = _RAND_1946[1:0];
  _RAND_1947 = {1{`RANDOM}};
  T_26182_19_lrs2_rtype = _RAND_1947[1:0];
  _RAND_1948 = {1{`RANDOM}};
  T_26182_19_frs3_en = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  T_26182_19_fp_val = _RAND_1949[0:0];
  _RAND_1950 = {1{`RANDOM}};
  T_26182_19_fp_single = _RAND_1950[0:0];
  _RAND_1951 = {1{`RANDOM}};
  T_26182_19_xcpt_if = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  T_26182_19_replay_if = _RAND_1952[0:0];
  _RAND_1953 = {2{`RANDOM}};
  T_26182_19_debug_wdata = _RAND_1953[63:0];
  _RAND_1954 = {1{`RANDOM}};
  T_26182_19_debug_events_fetch_seq = _RAND_1954[31:0];
  _RAND_1955 = {1{`RANDOM}};
  T_26182_20_valid = _RAND_1955[0:0];
  _RAND_1956 = {1{`RANDOM}};
  T_26182_20_iw_state = _RAND_1956[1:0];
  _RAND_1957 = {1{`RANDOM}};
  T_26182_20_uopc = _RAND_1957[8:0];
  _RAND_1958 = {1{`RANDOM}};
  T_26182_20_inst = _RAND_1958[31:0];
  _RAND_1959 = {2{`RANDOM}};
  T_26182_20_pc = _RAND_1959[39:0];
  _RAND_1960 = {1{`RANDOM}};
  T_26182_20_fu_code = _RAND_1960[7:0];
  _RAND_1961 = {1{`RANDOM}};
  T_26182_20_ctrl_br_type = _RAND_1961[3:0];
  _RAND_1962 = {1{`RANDOM}};
  T_26182_20_ctrl_op1_sel = _RAND_1962[1:0];
  _RAND_1963 = {1{`RANDOM}};
  T_26182_20_ctrl_op2_sel = _RAND_1963[2:0];
  _RAND_1964 = {1{`RANDOM}};
  T_26182_20_ctrl_imm_sel = _RAND_1964[2:0];
  _RAND_1965 = {1{`RANDOM}};
  T_26182_20_ctrl_op_fcn = _RAND_1965[3:0];
  _RAND_1966 = {1{`RANDOM}};
  T_26182_20_ctrl_fcn_dw = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  T_26182_20_ctrl_rf_wen = _RAND_1967[0:0];
  _RAND_1968 = {1{`RANDOM}};
  T_26182_20_ctrl_csr_cmd = _RAND_1968[2:0];
  _RAND_1969 = {1{`RANDOM}};
  T_26182_20_ctrl_is_load = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  T_26182_20_ctrl_is_sta = _RAND_1970[0:0];
  _RAND_1971 = {1{`RANDOM}};
  T_26182_20_ctrl_is_std = _RAND_1971[0:0];
  _RAND_1972 = {1{`RANDOM}};
  T_26182_20_wakeup_delay = _RAND_1972[1:0];
  _RAND_1973 = {1{`RANDOM}};
  T_26182_20_allocate_brtag = _RAND_1973[0:0];
  _RAND_1974 = {1{`RANDOM}};
  T_26182_20_is_br_or_jmp = _RAND_1974[0:0];
  _RAND_1975 = {1{`RANDOM}};
  T_26182_20_is_jump = _RAND_1975[0:0];
  _RAND_1976 = {1{`RANDOM}};
  T_26182_20_is_jal = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  T_26182_20_is_ret = _RAND_1977[0:0];
  _RAND_1978 = {1{`RANDOM}};
  T_26182_20_is_call = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  T_26182_20_br_mask = _RAND_1979[7:0];
  _RAND_1980 = {1{`RANDOM}};
  T_26182_20_br_tag = _RAND_1980[2:0];
  _RAND_1981 = {1{`RANDOM}};
  T_26182_20_br_prediction_bpd_predict_val = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  T_26182_20_br_prediction_bpd_predict_taken = _RAND_1982[0:0];
  _RAND_1983 = {1{`RANDOM}};
  T_26182_20_br_prediction_btb_hit = _RAND_1983[0:0];
  _RAND_1984 = {1{`RANDOM}};
  T_26182_20_br_prediction_btb_predicted = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  T_26182_20_br_prediction_is_br_or_jalr = _RAND_1985[0:0];
  _RAND_1986 = {1{`RANDOM}};
  T_26182_20_stat_brjmp_mispredicted = _RAND_1986[0:0];
  _RAND_1987 = {1{`RANDOM}};
  T_26182_20_stat_btb_made_pred = _RAND_1987[0:0];
  _RAND_1988 = {1{`RANDOM}};
  T_26182_20_stat_btb_mispredicted = _RAND_1988[0:0];
  _RAND_1989 = {1{`RANDOM}};
  T_26182_20_stat_bpd_made_pred = _RAND_1989[0:0];
  _RAND_1990 = {1{`RANDOM}};
  T_26182_20_stat_bpd_mispredicted = _RAND_1990[0:0];
  _RAND_1991 = {1{`RANDOM}};
  T_26182_20_fetch_pc_lob = _RAND_1991[2:0];
  _RAND_1992 = {1{`RANDOM}};
  T_26182_20_imm_packed = _RAND_1992[19:0];
  _RAND_1993 = {1{`RANDOM}};
  T_26182_20_csr_addr = _RAND_1993[11:0];
  _RAND_1994 = {1{`RANDOM}};
  T_26182_20_rob_idx = _RAND_1994[5:0];
  _RAND_1995 = {1{`RANDOM}};
  T_26182_20_ldq_idx = _RAND_1995[3:0];
  _RAND_1996 = {1{`RANDOM}};
  T_26182_20_stq_idx = _RAND_1996[3:0];
  _RAND_1997 = {1{`RANDOM}};
  T_26182_20_brob_idx = _RAND_1997[4:0];
  _RAND_1998 = {1{`RANDOM}};
  T_26182_20_pdst = _RAND_1998[6:0];
  _RAND_1999 = {1{`RANDOM}};
  T_26182_20_pop1 = _RAND_1999[6:0];
  _RAND_2000 = {1{`RANDOM}};
  T_26182_20_pop2 = _RAND_2000[6:0];
  _RAND_2001 = {1{`RANDOM}};
  T_26182_20_pop3 = _RAND_2001[6:0];
  _RAND_2002 = {1{`RANDOM}};
  T_26182_20_prs1_busy = _RAND_2002[0:0];
  _RAND_2003 = {1{`RANDOM}};
  T_26182_20_prs2_busy = _RAND_2003[0:0];
  _RAND_2004 = {1{`RANDOM}};
  T_26182_20_prs3_busy = _RAND_2004[0:0];
  _RAND_2005 = {1{`RANDOM}};
  T_26182_20_stale_pdst = _RAND_2005[6:0];
  _RAND_2006 = {1{`RANDOM}};
  T_26182_20_exception = _RAND_2006[0:0];
  _RAND_2007 = {2{`RANDOM}};
  T_26182_20_exc_cause = _RAND_2007[63:0];
  _RAND_2008 = {1{`RANDOM}};
  T_26182_20_bypassable = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  T_26182_20_mem_cmd = _RAND_2009[3:0];
  _RAND_2010 = {1{`RANDOM}};
  T_26182_20_mem_typ = _RAND_2010[2:0];
  _RAND_2011 = {1{`RANDOM}};
  T_26182_20_is_fence = _RAND_2011[0:0];
  _RAND_2012 = {1{`RANDOM}};
  T_26182_20_is_fencei = _RAND_2012[0:0];
  _RAND_2013 = {1{`RANDOM}};
  T_26182_20_is_store = _RAND_2013[0:0];
  _RAND_2014 = {1{`RANDOM}};
  T_26182_20_is_amo = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  T_26182_20_is_load = _RAND_2015[0:0];
  _RAND_2016 = {1{`RANDOM}};
  T_26182_20_is_unique = _RAND_2016[0:0];
  _RAND_2017 = {1{`RANDOM}};
  T_26182_20_flush_on_commit = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  T_26182_20_ldst = _RAND_2018[5:0];
  _RAND_2019 = {1{`RANDOM}};
  T_26182_20_lrs1 = _RAND_2019[5:0];
  _RAND_2020 = {1{`RANDOM}};
  T_26182_20_lrs2 = _RAND_2020[5:0];
  _RAND_2021 = {1{`RANDOM}};
  T_26182_20_lrs3 = _RAND_2021[5:0];
  _RAND_2022 = {1{`RANDOM}};
  T_26182_20_ldst_val = _RAND_2022[0:0];
  _RAND_2023 = {1{`RANDOM}};
  T_26182_20_dst_rtype = _RAND_2023[1:0];
  _RAND_2024 = {1{`RANDOM}};
  T_26182_20_lrs1_rtype = _RAND_2024[1:0];
  _RAND_2025 = {1{`RANDOM}};
  T_26182_20_lrs2_rtype = _RAND_2025[1:0];
  _RAND_2026 = {1{`RANDOM}};
  T_26182_20_frs3_en = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  T_26182_20_fp_val = _RAND_2027[0:0];
  _RAND_2028 = {1{`RANDOM}};
  T_26182_20_fp_single = _RAND_2028[0:0];
  _RAND_2029 = {1{`RANDOM}};
  T_26182_20_xcpt_if = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  T_26182_20_replay_if = _RAND_2030[0:0];
  _RAND_2031 = {2{`RANDOM}};
  T_26182_20_debug_wdata = _RAND_2031[63:0];
  _RAND_2032 = {1{`RANDOM}};
  T_26182_20_debug_events_fetch_seq = _RAND_2032[31:0];
  _RAND_2033 = {1{`RANDOM}};
  T_26182_21_valid = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  T_26182_21_iw_state = _RAND_2034[1:0];
  _RAND_2035 = {1{`RANDOM}};
  T_26182_21_uopc = _RAND_2035[8:0];
  _RAND_2036 = {1{`RANDOM}};
  T_26182_21_inst = _RAND_2036[31:0];
  _RAND_2037 = {2{`RANDOM}};
  T_26182_21_pc = _RAND_2037[39:0];
  _RAND_2038 = {1{`RANDOM}};
  T_26182_21_fu_code = _RAND_2038[7:0];
  _RAND_2039 = {1{`RANDOM}};
  T_26182_21_ctrl_br_type = _RAND_2039[3:0];
  _RAND_2040 = {1{`RANDOM}};
  T_26182_21_ctrl_op1_sel = _RAND_2040[1:0];
  _RAND_2041 = {1{`RANDOM}};
  T_26182_21_ctrl_op2_sel = _RAND_2041[2:0];
  _RAND_2042 = {1{`RANDOM}};
  T_26182_21_ctrl_imm_sel = _RAND_2042[2:0];
  _RAND_2043 = {1{`RANDOM}};
  T_26182_21_ctrl_op_fcn = _RAND_2043[3:0];
  _RAND_2044 = {1{`RANDOM}};
  T_26182_21_ctrl_fcn_dw = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  T_26182_21_ctrl_rf_wen = _RAND_2045[0:0];
  _RAND_2046 = {1{`RANDOM}};
  T_26182_21_ctrl_csr_cmd = _RAND_2046[2:0];
  _RAND_2047 = {1{`RANDOM}};
  T_26182_21_ctrl_is_load = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  T_26182_21_ctrl_is_sta = _RAND_2048[0:0];
  _RAND_2049 = {1{`RANDOM}};
  T_26182_21_ctrl_is_std = _RAND_2049[0:0];
  _RAND_2050 = {1{`RANDOM}};
  T_26182_21_wakeup_delay = _RAND_2050[1:0];
  _RAND_2051 = {1{`RANDOM}};
  T_26182_21_allocate_brtag = _RAND_2051[0:0];
  _RAND_2052 = {1{`RANDOM}};
  T_26182_21_is_br_or_jmp = _RAND_2052[0:0];
  _RAND_2053 = {1{`RANDOM}};
  T_26182_21_is_jump = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  T_26182_21_is_jal = _RAND_2054[0:0];
  _RAND_2055 = {1{`RANDOM}};
  T_26182_21_is_ret = _RAND_2055[0:0];
  _RAND_2056 = {1{`RANDOM}};
  T_26182_21_is_call = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  T_26182_21_br_mask = _RAND_2057[7:0];
  _RAND_2058 = {1{`RANDOM}};
  T_26182_21_br_tag = _RAND_2058[2:0];
  _RAND_2059 = {1{`RANDOM}};
  T_26182_21_br_prediction_bpd_predict_val = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  T_26182_21_br_prediction_bpd_predict_taken = _RAND_2060[0:0];
  _RAND_2061 = {1{`RANDOM}};
  T_26182_21_br_prediction_btb_hit = _RAND_2061[0:0];
  _RAND_2062 = {1{`RANDOM}};
  T_26182_21_br_prediction_btb_predicted = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  T_26182_21_br_prediction_is_br_or_jalr = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  T_26182_21_stat_brjmp_mispredicted = _RAND_2064[0:0];
  _RAND_2065 = {1{`RANDOM}};
  T_26182_21_stat_btb_made_pred = _RAND_2065[0:0];
  _RAND_2066 = {1{`RANDOM}};
  T_26182_21_stat_btb_mispredicted = _RAND_2066[0:0];
  _RAND_2067 = {1{`RANDOM}};
  T_26182_21_stat_bpd_made_pred = _RAND_2067[0:0];
  _RAND_2068 = {1{`RANDOM}};
  T_26182_21_stat_bpd_mispredicted = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  T_26182_21_fetch_pc_lob = _RAND_2069[2:0];
  _RAND_2070 = {1{`RANDOM}};
  T_26182_21_imm_packed = _RAND_2070[19:0];
  _RAND_2071 = {1{`RANDOM}};
  T_26182_21_csr_addr = _RAND_2071[11:0];
  _RAND_2072 = {1{`RANDOM}};
  T_26182_21_rob_idx = _RAND_2072[5:0];
  _RAND_2073 = {1{`RANDOM}};
  T_26182_21_ldq_idx = _RAND_2073[3:0];
  _RAND_2074 = {1{`RANDOM}};
  T_26182_21_stq_idx = _RAND_2074[3:0];
  _RAND_2075 = {1{`RANDOM}};
  T_26182_21_brob_idx = _RAND_2075[4:0];
  _RAND_2076 = {1{`RANDOM}};
  T_26182_21_pdst = _RAND_2076[6:0];
  _RAND_2077 = {1{`RANDOM}};
  T_26182_21_pop1 = _RAND_2077[6:0];
  _RAND_2078 = {1{`RANDOM}};
  T_26182_21_pop2 = _RAND_2078[6:0];
  _RAND_2079 = {1{`RANDOM}};
  T_26182_21_pop3 = _RAND_2079[6:0];
  _RAND_2080 = {1{`RANDOM}};
  T_26182_21_prs1_busy = _RAND_2080[0:0];
  _RAND_2081 = {1{`RANDOM}};
  T_26182_21_prs2_busy = _RAND_2081[0:0];
  _RAND_2082 = {1{`RANDOM}};
  T_26182_21_prs3_busy = _RAND_2082[0:0];
  _RAND_2083 = {1{`RANDOM}};
  T_26182_21_stale_pdst = _RAND_2083[6:0];
  _RAND_2084 = {1{`RANDOM}};
  T_26182_21_exception = _RAND_2084[0:0];
  _RAND_2085 = {2{`RANDOM}};
  T_26182_21_exc_cause = _RAND_2085[63:0];
  _RAND_2086 = {1{`RANDOM}};
  T_26182_21_bypassable = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  T_26182_21_mem_cmd = _RAND_2087[3:0];
  _RAND_2088 = {1{`RANDOM}};
  T_26182_21_mem_typ = _RAND_2088[2:0];
  _RAND_2089 = {1{`RANDOM}};
  T_26182_21_is_fence = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  T_26182_21_is_fencei = _RAND_2090[0:0];
  _RAND_2091 = {1{`RANDOM}};
  T_26182_21_is_store = _RAND_2091[0:0];
  _RAND_2092 = {1{`RANDOM}};
  T_26182_21_is_amo = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  T_26182_21_is_load = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  T_26182_21_is_unique = _RAND_2094[0:0];
  _RAND_2095 = {1{`RANDOM}};
  T_26182_21_flush_on_commit = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  T_26182_21_ldst = _RAND_2096[5:0];
  _RAND_2097 = {1{`RANDOM}};
  T_26182_21_lrs1 = _RAND_2097[5:0];
  _RAND_2098 = {1{`RANDOM}};
  T_26182_21_lrs2 = _RAND_2098[5:0];
  _RAND_2099 = {1{`RANDOM}};
  T_26182_21_lrs3 = _RAND_2099[5:0];
  _RAND_2100 = {1{`RANDOM}};
  T_26182_21_ldst_val = _RAND_2100[0:0];
  _RAND_2101 = {1{`RANDOM}};
  T_26182_21_dst_rtype = _RAND_2101[1:0];
  _RAND_2102 = {1{`RANDOM}};
  T_26182_21_lrs1_rtype = _RAND_2102[1:0];
  _RAND_2103 = {1{`RANDOM}};
  T_26182_21_lrs2_rtype = _RAND_2103[1:0];
  _RAND_2104 = {1{`RANDOM}};
  T_26182_21_frs3_en = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  T_26182_21_fp_val = _RAND_2105[0:0];
  _RAND_2106 = {1{`RANDOM}};
  T_26182_21_fp_single = _RAND_2106[0:0];
  _RAND_2107 = {1{`RANDOM}};
  T_26182_21_xcpt_if = _RAND_2107[0:0];
  _RAND_2108 = {1{`RANDOM}};
  T_26182_21_replay_if = _RAND_2108[0:0];
  _RAND_2109 = {2{`RANDOM}};
  T_26182_21_debug_wdata = _RAND_2109[63:0];
  _RAND_2110 = {1{`RANDOM}};
  T_26182_21_debug_events_fetch_seq = _RAND_2110[31:0];
  _RAND_2111 = {1{`RANDOM}};
  T_26182_22_valid = _RAND_2111[0:0];
  _RAND_2112 = {1{`RANDOM}};
  T_26182_22_iw_state = _RAND_2112[1:0];
  _RAND_2113 = {1{`RANDOM}};
  T_26182_22_uopc = _RAND_2113[8:0];
  _RAND_2114 = {1{`RANDOM}};
  T_26182_22_inst = _RAND_2114[31:0];
  _RAND_2115 = {2{`RANDOM}};
  T_26182_22_pc = _RAND_2115[39:0];
  _RAND_2116 = {1{`RANDOM}};
  T_26182_22_fu_code = _RAND_2116[7:0];
  _RAND_2117 = {1{`RANDOM}};
  T_26182_22_ctrl_br_type = _RAND_2117[3:0];
  _RAND_2118 = {1{`RANDOM}};
  T_26182_22_ctrl_op1_sel = _RAND_2118[1:0];
  _RAND_2119 = {1{`RANDOM}};
  T_26182_22_ctrl_op2_sel = _RAND_2119[2:0];
  _RAND_2120 = {1{`RANDOM}};
  T_26182_22_ctrl_imm_sel = _RAND_2120[2:0];
  _RAND_2121 = {1{`RANDOM}};
  T_26182_22_ctrl_op_fcn = _RAND_2121[3:0];
  _RAND_2122 = {1{`RANDOM}};
  T_26182_22_ctrl_fcn_dw = _RAND_2122[0:0];
  _RAND_2123 = {1{`RANDOM}};
  T_26182_22_ctrl_rf_wen = _RAND_2123[0:0];
  _RAND_2124 = {1{`RANDOM}};
  T_26182_22_ctrl_csr_cmd = _RAND_2124[2:0];
  _RAND_2125 = {1{`RANDOM}};
  T_26182_22_ctrl_is_load = _RAND_2125[0:0];
  _RAND_2126 = {1{`RANDOM}};
  T_26182_22_ctrl_is_sta = _RAND_2126[0:0];
  _RAND_2127 = {1{`RANDOM}};
  T_26182_22_ctrl_is_std = _RAND_2127[0:0];
  _RAND_2128 = {1{`RANDOM}};
  T_26182_22_wakeup_delay = _RAND_2128[1:0];
  _RAND_2129 = {1{`RANDOM}};
  T_26182_22_allocate_brtag = _RAND_2129[0:0];
  _RAND_2130 = {1{`RANDOM}};
  T_26182_22_is_br_or_jmp = _RAND_2130[0:0];
  _RAND_2131 = {1{`RANDOM}};
  T_26182_22_is_jump = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  T_26182_22_is_jal = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  T_26182_22_is_ret = _RAND_2133[0:0];
  _RAND_2134 = {1{`RANDOM}};
  T_26182_22_is_call = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  T_26182_22_br_mask = _RAND_2135[7:0];
  _RAND_2136 = {1{`RANDOM}};
  T_26182_22_br_tag = _RAND_2136[2:0];
  _RAND_2137 = {1{`RANDOM}};
  T_26182_22_br_prediction_bpd_predict_val = _RAND_2137[0:0];
  _RAND_2138 = {1{`RANDOM}};
  T_26182_22_br_prediction_bpd_predict_taken = _RAND_2138[0:0];
  _RAND_2139 = {1{`RANDOM}};
  T_26182_22_br_prediction_btb_hit = _RAND_2139[0:0];
  _RAND_2140 = {1{`RANDOM}};
  T_26182_22_br_prediction_btb_predicted = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  T_26182_22_br_prediction_is_br_or_jalr = _RAND_2141[0:0];
  _RAND_2142 = {1{`RANDOM}};
  T_26182_22_stat_brjmp_mispredicted = _RAND_2142[0:0];
  _RAND_2143 = {1{`RANDOM}};
  T_26182_22_stat_btb_made_pred = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  T_26182_22_stat_btb_mispredicted = _RAND_2144[0:0];
  _RAND_2145 = {1{`RANDOM}};
  T_26182_22_stat_bpd_made_pred = _RAND_2145[0:0];
  _RAND_2146 = {1{`RANDOM}};
  T_26182_22_stat_bpd_mispredicted = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  T_26182_22_fetch_pc_lob = _RAND_2147[2:0];
  _RAND_2148 = {1{`RANDOM}};
  T_26182_22_imm_packed = _RAND_2148[19:0];
  _RAND_2149 = {1{`RANDOM}};
  T_26182_22_csr_addr = _RAND_2149[11:0];
  _RAND_2150 = {1{`RANDOM}};
  T_26182_22_rob_idx = _RAND_2150[5:0];
  _RAND_2151 = {1{`RANDOM}};
  T_26182_22_ldq_idx = _RAND_2151[3:0];
  _RAND_2152 = {1{`RANDOM}};
  T_26182_22_stq_idx = _RAND_2152[3:0];
  _RAND_2153 = {1{`RANDOM}};
  T_26182_22_brob_idx = _RAND_2153[4:0];
  _RAND_2154 = {1{`RANDOM}};
  T_26182_22_pdst = _RAND_2154[6:0];
  _RAND_2155 = {1{`RANDOM}};
  T_26182_22_pop1 = _RAND_2155[6:0];
  _RAND_2156 = {1{`RANDOM}};
  T_26182_22_pop2 = _RAND_2156[6:0];
  _RAND_2157 = {1{`RANDOM}};
  T_26182_22_pop3 = _RAND_2157[6:0];
  _RAND_2158 = {1{`RANDOM}};
  T_26182_22_prs1_busy = _RAND_2158[0:0];
  _RAND_2159 = {1{`RANDOM}};
  T_26182_22_prs2_busy = _RAND_2159[0:0];
  _RAND_2160 = {1{`RANDOM}};
  T_26182_22_prs3_busy = _RAND_2160[0:0];
  _RAND_2161 = {1{`RANDOM}};
  T_26182_22_stale_pdst = _RAND_2161[6:0];
  _RAND_2162 = {1{`RANDOM}};
  T_26182_22_exception = _RAND_2162[0:0];
  _RAND_2163 = {2{`RANDOM}};
  T_26182_22_exc_cause = _RAND_2163[63:0];
  _RAND_2164 = {1{`RANDOM}};
  T_26182_22_bypassable = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  T_26182_22_mem_cmd = _RAND_2165[3:0];
  _RAND_2166 = {1{`RANDOM}};
  T_26182_22_mem_typ = _RAND_2166[2:0];
  _RAND_2167 = {1{`RANDOM}};
  T_26182_22_is_fence = _RAND_2167[0:0];
  _RAND_2168 = {1{`RANDOM}};
  T_26182_22_is_fencei = _RAND_2168[0:0];
  _RAND_2169 = {1{`RANDOM}};
  T_26182_22_is_store = _RAND_2169[0:0];
  _RAND_2170 = {1{`RANDOM}};
  T_26182_22_is_amo = _RAND_2170[0:0];
  _RAND_2171 = {1{`RANDOM}};
  T_26182_22_is_load = _RAND_2171[0:0];
  _RAND_2172 = {1{`RANDOM}};
  T_26182_22_is_unique = _RAND_2172[0:0];
  _RAND_2173 = {1{`RANDOM}};
  T_26182_22_flush_on_commit = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  T_26182_22_ldst = _RAND_2174[5:0];
  _RAND_2175 = {1{`RANDOM}};
  T_26182_22_lrs1 = _RAND_2175[5:0];
  _RAND_2176 = {1{`RANDOM}};
  T_26182_22_lrs2 = _RAND_2176[5:0];
  _RAND_2177 = {1{`RANDOM}};
  T_26182_22_lrs3 = _RAND_2177[5:0];
  _RAND_2178 = {1{`RANDOM}};
  T_26182_22_ldst_val = _RAND_2178[0:0];
  _RAND_2179 = {1{`RANDOM}};
  T_26182_22_dst_rtype = _RAND_2179[1:0];
  _RAND_2180 = {1{`RANDOM}};
  T_26182_22_lrs1_rtype = _RAND_2180[1:0];
  _RAND_2181 = {1{`RANDOM}};
  T_26182_22_lrs2_rtype = _RAND_2181[1:0];
  _RAND_2182 = {1{`RANDOM}};
  T_26182_22_frs3_en = _RAND_2182[0:0];
  _RAND_2183 = {1{`RANDOM}};
  T_26182_22_fp_val = _RAND_2183[0:0];
  _RAND_2184 = {1{`RANDOM}};
  T_26182_22_fp_single = _RAND_2184[0:0];
  _RAND_2185 = {1{`RANDOM}};
  T_26182_22_xcpt_if = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  T_26182_22_replay_if = _RAND_2186[0:0];
  _RAND_2187 = {2{`RANDOM}};
  T_26182_22_debug_wdata = _RAND_2187[63:0];
  _RAND_2188 = {1{`RANDOM}};
  T_26182_22_debug_events_fetch_seq = _RAND_2188[31:0];
  _RAND_2189 = {1{`RANDOM}};
  T_26182_23_valid = _RAND_2189[0:0];
  _RAND_2190 = {1{`RANDOM}};
  T_26182_23_iw_state = _RAND_2190[1:0];
  _RAND_2191 = {1{`RANDOM}};
  T_26182_23_uopc = _RAND_2191[8:0];
  _RAND_2192 = {1{`RANDOM}};
  T_26182_23_inst = _RAND_2192[31:0];
  _RAND_2193 = {2{`RANDOM}};
  T_26182_23_pc = _RAND_2193[39:0];
  _RAND_2194 = {1{`RANDOM}};
  T_26182_23_fu_code = _RAND_2194[7:0];
  _RAND_2195 = {1{`RANDOM}};
  T_26182_23_ctrl_br_type = _RAND_2195[3:0];
  _RAND_2196 = {1{`RANDOM}};
  T_26182_23_ctrl_op1_sel = _RAND_2196[1:0];
  _RAND_2197 = {1{`RANDOM}};
  T_26182_23_ctrl_op2_sel = _RAND_2197[2:0];
  _RAND_2198 = {1{`RANDOM}};
  T_26182_23_ctrl_imm_sel = _RAND_2198[2:0];
  _RAND_2199 = {1{`RANDOM}};
  T_26182_23_ctrl_op_fcn = _RAND_2199[3:0];
  _RAND_2200 = {1{`RANDOM}};
  T_26182_23_ctrl_fcn_dw = _RAND_2200[0:0];
  _RAND_2201 = {1{`RANDOM}};
  T_26182_23_ctrl_rf_wen = _RAND_2201[0:0];
  _RAND_2202 = {1{`RANDOM}};
  T_26182_23_ctrl_csr_cmd = _RAND_2202[2:0];
  _RAND_2203 = {1{`RANDOM}};
  T_26182_23_ctrl_is_load = _RAND_2203[0:0];
  _RAND_2204 = {1{`RANDOM}};
  T_26182_23_ctrl_is_sta = _RAND_2204[0:0];
  _RAND_2205 = {1{`RANDOM}};
  T_26182_23_ctrl_is_std = _RAND_2205[0:0];
  _RAND_2206 = {1{`RANDOM}};
  T_26182_23_wakeup_delay = _RAND_2206[1:0];
  _RAND_2207 = {1{`RANDOM}};
  T_26182_23_allocate_brtag = _RAND_2207[0:0];
  _RAND_2208 = {1{`RANDOM}};
  T_26182_23_is_br_or_jmp = _RAND_2208[0:0];
  _RAND_2209 = {1{`RANDOM}};
  T_26182_23_is_jump = _RAND_2209[0:0];
  _RAND_2210 = {1{`RANDOM}};
  T_26182_23_is_jal = _RAND_2210[0:0];
  _RAND_2211 = {1{`RANDOM}};
  T_26182_23_is_ret = _RAND_2211[0:0];
  _RAND_2212 = {1{`RANDOM}};
  T_26182_23_is_call = _RAND_2212[0:0];
  _RAND_2213 = {1{`RANDOM}};
  T_26182_23_br_mask = _RAND_2213[7:0];
  _RAND_2214 = {1{`RANDOM}};
  T_26182_23_br_tag = _RAND_2214[2:0];
  _RAND_2215 = {1{`RANDOM}};
  T_26182_23_br_prediction_bpd_predict_val = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  T_26182_23_br_prediction_bpd_predict_taken = _RAND_2216[0:0];
  _RAND_2217 = {1{`RANDOM}};
  T_26182_23_br_prediction_btb_hit = _RAND_2217[0:0];
  _RAND_2218 = {1{`RANDOM}};
  T_26182_23_br_prediction_btb_predicted = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  T_26182_23_br_prediction_is_br_or_jalr = _RAND_2219[0:0];
  _RAND_2220 = {1{`RANDOM}};
  T_26182_23_stat_brjmp_mispredicted = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  T_26182_23_stat_btb_made_pred = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  T_26182_23_stat_btb_mispredicted = _RAND_2222[0:0];
  _RAND_2223 = {1{`RANDOM}};
  T_26182_23_stat_bpd_made_pred = _RAND_2223[0:0];
  _RAND_2224 = {1{`RANDOM}};
  T_26182_23_stat_bpd_mispredicted = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  T_26182_23_fetch_pc_lob = _RAND_2225[2:0];
  _RAND_2226 = {1{`RANDOM}};
  T_26182_23_imm_packed = _RAND_2226[19:0];
  _RAND_2227 = {1{`RANDOM}};
  T_26182_23_csr_addr = _RAND_2227[11:0];
  _RAND_2228 = {1{`RANDOM}};
  T_26182_23_rob_idx = _RAND_2228[5:0];
  _RAND_2229 = {1{`RANDOM}};
  T_26182_23_ldq_idx = _RAND_2229[3:0];
  _RAND_2230 = {1{`RANDOM}};
  T_26182_23_stq_idx = _RAND_2230[3:0];
  _RAND_2231 = {1{`RANDOM}};
  T_26182_23_brob_idx = _RAND_2231[4:0];
  _RAND_2232 = {1{`RANDOM}};
  T_26182_23_pdst = _RAND_2232[6:0];
  _RAND_2233 = {1{`RANDOM}};
  T_26182_23_pop1 = _RAND_2233[6:0];
  _RAND_2234 = {1{`RANDOM}};
  T_26182_23_pop2 = _RAND_2234[6:0];
  _RAND_2235 = {1{`RANDOM}};
  T_26182_23_pop3 = _RAND_2235[6:0];
  _RAND_2236 = {1{`RANDOM}};
  T_26182_23_prs1_busy = _RAND_2236[0:0];
  _RAND_2237 = {1{`RANDOM}};
  T_26182_23_prs2_busy = _RAND_2237[0:0];
  _RAND_2238 = {1{`RANDOM}};
  T_26182_23_prs3_busy = _RAND_2238[0:0];
  _RAND_2239 = {1{`RANDOM}};
  T_26182_23_stale_pdst = _RAND_2239[6:0];
  _RAND_2240 = {1{`RANDOM}};
  T_26182_23_exception = _RAND_2240[0:0];
  _RAND_2241 = {2{`RANDOM}};
  T_26182_23_exc_cause = _RAND_2241[63:0];
  _RAND_2242 = {1{`RANDOM}};
  T_26182_23_bypassable = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  T_26182_23_mem_cmd = _RAND_2243[3:0];
  _RAND_2244 = {1{`RANDOM}};
  T_26182_23_mem_typ = _RAND_2244[2:0];
  _RAND_2245 = {1{`RANDOM}};
  T_26182_23_is_fence = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  T_26182_23_is_fencei = _RAND_2246[0:0];
  _RAND_2247 = {1{`RANDOM}};
  T_26182_23_is_store = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  T_26182_23_is_amo = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  T_26182_23_is_load = _RAND_2249[0:0];
  _RAND_2250 = {1{`RANDOM}};
  T_26182_23_is_unique = _RAND_2250[0:0];
  _RAND_2251 = {1{`RANDOM}};
  T_26182_23_flush_on_commit = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  T_26182_23_ldst = _RAND_2252[5:0];
  _RAND_2253 = {1{`RANDOM}};
  T_26182_23_lrs1 = _RAND_2253[5:0];
  _RAND_2254 = {1{`RANDOM}};
  T_26182_23_lrs2 = _RAND_2254[5:0];
  _RAND_2255 = {1{`RANDOM}};
  T_26182_23_lrs3 = _RAND_2255[5:0];
  _RAND_2256 = {1{`RANDOM}};
  T_26182_23_ldst_val = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  T_26182_23_dst_rtype = _RAND_2257[1:0];
  _RAND_2258 = {1{`RANDOM}};
  T_26182_23_lrs1_rtype = _RAND_2258[1:0];
  _RAND_2259 = {1{`RANDOM}};
  T_26182_23_lrs2_rtype = _RAND_2259[1:0];
  _RAND_2260 = {1{`RANDOM}};
  T_26182_23_frs3_en = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  T_26182_23_fp_val = _RAND_2261[0:0];
  _RAND_2262 = {1{`RANDOM}};
  T_26182_23_fp_single = _RAND_2262[0:0];
  _RAND_2263 = {1{`RANDOM}};
  T_26182_23_xcpt_if = _RAND_2263[0:0];
  _RAND_2264 = {1{`RANDOM}};
  T_26182_23_replay_if = _RAND_2264[0:0];
  _RAND_2265 = {2{`RANDOM}};
  T_26182_23_debug_wdata = _RAND_2265[63:0];
  _RAND_2266 = {1{`RANDOM}};
  T_26182_23_debug_events_fetch_seq = _RAND_2266[31:0];
  _RAND_2267 = {1{`RANDOM}};
  T_38110_0_valid = _RAND_2267[0:0];
  _RAND_2268 = {1{`RANDOM}};
  T_38110_0_iw_state = _RAND_2268[1:0];
  _RAND_2269 = {1{`RANDOM}};
  T_38110_0_uopc = _RAND_2269[8:0];
  _RAND_2270 = {1{`RANDOM}};
  T_38110_0_inst = _RAND_2270[31:0];
  _RAND_2271 = {2{`RANDOM}};
  T_38110_0_pc = _RAND_2271[39:0];
  _RAND_2272 = {1{`RANDOM}};
  T_38110_0_fu_code = _RAND_2272[7:0];
  _RAND_2273 = {1{`RANDOM}};
  T_38110_0_ctrl_br_type = _RAND_2273[3:0];
  _RAND_2274 = {1{`RANDOM}};
  T_38110_0_ctrl_op1_sel = _RAND_2274[1:0];
  _RAND_2275 = {1{`RANDOM}};
  T_38110_0_ctrl_op2_sel = _RAND_2275[2:0];
  _RAND_2276 = {1{`RANDOM}};
  T_38110_0_ctrl_imm_sel = _RAND_2276[2:0];
  _RAND_2277 = {1{`RANDOM}};
  T_38110_0_ctrl_op_fcn = _RAND_2277[3:0];
  _RAND_2278 = {1{`RANDOM}};
  T_38110_0_ctrl_fcn_dw = _RAND_2278[0:0];
  _RAND_2279 = {1{`RANDOM}};
  T_38110_0_ctrl_rf_wen = _RAND_2279[0:0];
  _RAND_2280 = {1{`RANDOM}};
  T_38110_0_ctrl_csr_cmd = _RAND_2280[2:0];
  _RAND_2281 = {1{`RANDOM}};
  T_38110_0_ctrl_is_load = _RAND_2281[0:0];
  _RAND_2282 = {1{`RANDOM}};
  T_38110_0_ctrl_is_sta = _RAND_2282[0:0];
  _RAND_2283 = {1{`RANDOM}};
  T_38110_0_ctrl_is_std = _RAND_2283[0:0];
  _RAND_2284 = {1{`RANDOM}};
  T_38110_0_wakeup_delay = _RAND_2284[1:0];
  _RAND_2285 = {1{`RANDOM}};
  T_38110_0_allocate_brtag = _RAND_2285[0:0];
  _RAND_2286 = {1{`RANDOM}};
  T_38110_0_is_br_or_jmp = _RAND_2286[0:0];
  _RAND_2287 = {1{`RANDOM}};
  T_38110_0_is_jump = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  T_38110_0_is_jal = _RAND_2288[0:0];
  _RAND_2289 = {1{`RANDOM}};
  T_38110_0_is_ret = _RAND_2289[0:0];
  _RAND_2290 = {1{`RANDOM}};
  T_38110_0_is_call = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  T_38110_0_br_mask = _RAND_2291[7:0];
  _RAND_2292 = {1{`RANDOM}};
  T_38110_0_br_tag = _RAND_2292[2:0];
  _RAND_2293 = {1{`RANDOM}};
  T_38110_0_br_prediction_bpd_predict_val = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  T_38110_0_br_prediction_bpd_predict_taken = _RAND_2294[0:0];
  _RAND_2295 = {1{`RANDOM}};
  T_38110_0_br_prediction_btb_hit = _RAND_2295[0:0];
  _RAND_2296 = {1{`RANDOM}};
  T_38110_0_br_prediction_btb_predicted = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  T_38110_0_br_prediction_is_br_or_jalr = _RAND_2297[0:0];
  _RAND_2298 = {1{`RANDOM}};
  T_38110_0_stat_brjmp_mispredicted = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  T_38110_0_stat_btb_made_pred = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  T_38110_0_stat_btb_mispredicted = _RAND_2300[0:0];
  _RAND_2301 = {1{`RANDOM}};
  T_38110_0_stat_bpd_made_pred = _RAND_2301[0:0];
  _RAND_2302 = {1{`RANDOM}};
  T_38110_0_stat_bpd_mispredicted = _RAND_2302[0:0];
  _RAND_2303 = {1{`RANDOM}};
  T_38110_0_fetch_pc_lob = _RAND_2303[2:0];
  _RAND_2304 = {1{`RANDOM}};
  T_38110_0_imm_packed = _RAND_2304[19:0];
  _RAND_2305 = {1{`RANDOM}};
  T_38110_0_csr_addr = _RAND_2305[11:0];
  _RAND_2306 = {1{`RANDOM}};
  T_38110_0_rob_idx = _RAND_2306[5:0];
  _RAND_2307 = {1{`RANDOM}};
  T_38110_0_ldq_idx = _RAND_2307[3:0];
  _RAND_2308 = {1{`RANDOM}};
  T_38110_0_stq_idx = _RAND_2308[3:0];
  _RAND_2309 = {1{`RANDOM}};
  T_38110_0_brob_idx = _RAND_2309[4:0];
  _RAND_2310 = {1{`RANDOM}};
  T_38110_0_pdst = _RAND_2310[6:0];
  _RAND_2311 = {1{`RANDOM}};
  T_38110_0_pop1 = _RAND_2311[6:0];
  _RAND_2312 = {1{`RANDOM}};
  T_38110_0_pop2 = _RAND_2312[6:0];
  _RAND_2313 = {1{`RANDOM}};
  T_38110_0_pop3 = _RAND_2313[6:0];
  _RAND_2314 = {1{`RANDOM}};
  T_38110_0_prs1_busy = _RAND_2314[0:0];
  _RAND_2315 = {1{`RANDOM}};
  T_38110_0_prs2_busy = _RAND_2315[0:0];
  _RAND_2316 = {1{`RANDOM}};
  T_38110_0_prs3_busy = _RAND_2316[0:0];
  _RAND_2317 = {1{`RANDOM}};
  T_38110_0_stale_pdst = _RAND_2317[6:0];
  _RAND_2318 = {1{`RANDOM}};
  T_38110_0_exception = _RAND_2318[0:0];
  _RAND_2319 = {2{`RANDOM}};
  T_38110_0_exc_cause = _RAND_2319[63:0];
  _RAND_2320 = {1{`RANDOM}};
  T_38110_0_bypassable = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  T_38110_0_mem_cmd = _RAND_2321[3:0];
  _RAND_2322 = {1{`RANDOM}};
  T_38110_0_mem_typ = _RAND_2322[2:0];
  _RAND_2323 = {1{`RANDOM}};
  T_38110_0_is_fence = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  T_38110_0_is_fencei = _RAND_2324[0:0];
  _RAND_2325 = {1{`RANDOM}};
  T_38110_0_is_store = _RAND_2325[0:0];
  _RAND_2326 = {1{`RANDOM}};
  T_38110_0_is_amo = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  T_38110_0_is_load = _RAND_2327[0:0];
  _RAND_2328 = {1{`RANDOM}};
  T_38110_0_is_unique = _RAND_2328[0:0];
  _RAND_2329 = {1{`RANDOM}};
  T_38110_0_flush_on_commit = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  T_38110_0_ldst = _RAND_2330[5:0];
  _RAND_2331 = {1{`RANDOM}};
  T_38110_0_lrs1 = _RAND_2331[5:0];
  _RAND_2332 = {1{`RANDOM}};
  T_38110_0_lrs2 = _RAND_2332[5:0];
  _RAND_2333 = {1{`RANDOM}};
  T_38110_0_lrs3 = _RAND_2333[5:0];
  _RAND_2334 = {1{`RANDOM}};
  T_38110_0_ldst_val = _RAND_2334[0:0];
  _RAND_2335 = {1{`RANDOM}};
  T_38110_0_dst_rtype = _RAND_2335[1:0];
  _RAND_2336 = {1{`RANDOM}};
  T_38110_0_lrs1_rtype = _RAND_2336[1:0];
  _RAND_2337 = {1{`RANDOM}};
  T_38110_0_lrs2_rtype = _RAND_2337[1:0];
  _RAND_2338 = {1{`RANDOM}};
  T_38110_0_frs3_en = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  T_38110_0_fp_val = _RAND_2339[0:0];
  _RAND_2340 = {1{`RANDOM}};
  T_38110_0_fp_single = _RAND_2340[0:0];
  _RAND_2341 = {1{`RANDOM}};
  T_38110_0_xcpt_if = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  T_38110_0_replay_if = _RAND_2342[0:0];
  _RAND_2343 = {2{`RANDOM}};
  T_38110_0_debug_wdata = _RAND_2343[63:0];
  _RAND_2344 = {1{`RANDOM}};
  T_38110_0_debug_events_fetch_seq = _RAND_2344[31:0];
  _RAND_2345 = {1{`RANDOM}};
  T_38110_1_valid = _RAND_2345[0:0];
  _RAND_2346 = {1{`RANDOM}};
  T_38110_1_iw_state = _RAND_2346[1:0];
  _RAND_2347 = {1{`RANDOM}};
  T_38110_1_uopc = _RAND_2347[8:0];
  _RAND_2348 = {1{`RANDOM}};
  T_38110_1_inst = _RAND_2348[31:0];
  _RAND_2349 = {2{`RANDOM}};
  T_38110_1_pc = _RAND_2349[39:0];
  _RAND_2350 = {1{`RANDOM}};
  T_38110_1_fu_code = _RAND_2350[7:0];
  _RAND_2351 = {1{`RANDOM}};
  T_38110_1_ctrl_br_type = _RAND_2351[3:0];
  _RAND_2352 = {1{`RANDOM}};
  T_38110_1_ctrl_op1_sel = _RAND_2352[1:0];
  _RAND_2353 = {1{`RANDOM}};
  T_38110_1_ctrl_op2_sel = _RAND_2353[2:0];
  _RAND_2354 = {1{`RANDOM}};
  T_38110_1_ctrl_imm_sel = _RAND_2354[2:0];
  _RAND_2355 = {1{`RANDOM}};
  T_38110_1_ctrl_op_fcn = _RAND_2355[3:0];
  _RAND_2356 = {1{`RANDOM}};
  T_38110_1_ctrl_fcn_dw = _RAND_2356[0:0];
  _RAND_2357 = {1{`RANDOM}};
  T_38110_1_ctrl_rf_wen = _RAND_2357[0:0];
  _RAND_2358 = {1{`RANDOM}};
  T_38110_1_ctrl_csr_cmd = _RAND_2358[2:0];
  _RAND_2359 = {1{`RANDOM}};
  T_38110_1_ctrl_is_load = _RAND_2359[0:0];
  _RAND_2360 = {1{`RANDOM}};
  T_38110_1_ctrl_is_sta = _RAND_2360[0:0];
  _RAND_2361 = {1{`RANDOM}};
  T_38110_1_ctrl_is_std = _RAND_2361[0:0];
  _RAND_2362 = {1{`RANDOM}};
  T_38110_1_wakeup_delay = _RAND_2362[1:0];
  _RAND_2363 = {1{`RANDOM}};
  T_38110_1_allocate_brtag = _RAND_2363[0:0];
  _RAND_2364 = {1{`RANDOM}};
  T_38110_1_is_br_or_jmp = _RAND_2364[0:0];
  _RAND_2365 = {1{`RANDOM}};
  T_38110_1_is_jump = _RAND_2365[0:0];
  _RAND_2366 = {1{`RANDOM}};
  T_38110_1_is_jal = _RAND_2366[0:0];
  _RAND_2367 = {1{`RANDOM}};
  T_38110_1_is_ret = _RAND_2367[0:0];
  _RAND_2368 = {1{`RANDOM}};
  T_38110_1_is_call = _RAND_2368[0:0];
  _RAND_2369 = {1{`RANDOM}};
  T_38110_1_br_mask = _RAND_2369[7:0];
  _RAND_2370 = {1{`RANDOM}};
  T_38110_1_br_tag = _RAND_2370[2:0];
  _RAND_2371 = {1{`RANDOM}};
  T_38110_1_br_prediction_bpd_predict_val = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  T_38110_1_br_prediction_bpd_predict_taken = _RAND_2372[0:0];
  _RAND_2373 = {1{`RANDOM}};
  T_38110_1_br_prediction_btb_hit = _RAND_2373[0:0];
  _RAND_2374 = {1{`RANDOM}};
  T_38110_1_br_prediction_btb_predicted = _RAND_2374[0:0];
  _RAND_2375 = {1{`RANDOM}};
  T_38110_1_br_prediction_is_br_or_jalr = _RAND_2375[0:0];
  _RAND_2376 = {1{`RANDOM}};
  T_38110_1_stat_brjmp_mispredicted = _RAND_2376[0:0];
  _RAND_2377 = {1{`RANDOM}};
  T_38110_1_stat_btb_made_pred = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  T_38110_1_stat_btb_mispredicted = _RAND_2378[0:0];
  _RAND_2379 = {1{`RANDOM}};
  T_38110_1_stat_bpd_made_pred = _RAND_2379[0:0];
  _RAND_2380 = {1{`RANDOM}};
  T_38110_1_stat_bpd_mispredicted = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  T_38110_1_fetch_pc_lob = _RAND_2381[2:0];
  _RAND_2382 = {1{`RANDOM}};
  T_38110_1_imm_packed = _RAND_2382[19:0];
  _RAND_2383 = {1{`RANDOM}};
  T_38110_1_csr_addr = _RAND_2383[11:0];
  _RAND_2384 = {1{`RANDOM}};
  T_38110_1_rob_idx = _RAND_2384[5:0];
  _RAND_2385 = {1{`RANDOM}};
  T_38110_1_ldq_idx = _RAND_2385[3:0];
  _RAND_2386 = {1{`RANDOM}};
  T_38110_1_stq_idx = _RAND_2386[3:0];
  _RAND_2387 = {1{`RANDOM}};
  T_38110_1_brob_idx = _RAND_2387[4:0];
  _RAND_2388 = {1{`RANDOM}};
  T_38110_1_pdst = _RAND_2388[6:0];
  _RAND_2389 = {1{`RANDOM}};
  T_38110_1_pop1 = _RAND_2389[6:0];
  _RAND_2390 = {1{`RANDOM}};
  T_38110_1_pop2 = _RAND_2390[6:0];
  _RAND_2391 = {1{`RANDOM}};
  T_38110_1_pop3 = _RAND_2391[6:0];
  _RAND_2392 = {1{`RANDOM}};
  T_38110_1_prs1_busy = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  T_38110_1_prs2_busy = _RAND_2393[0:0];
  _RAND_2394 = {1{`RANDOM}};
  T_38110_1_prs3_busy = _RAND_2394[0:0];
  _RAND_2395 = {1{`RANDOM}};
  T_38110_1_stale_pdst = _RAND_2395[6:0];
  _RAND_2396 = {1{`RANDOM}};
  T_38110_1_exception = _RAND_2396[0:0];
  _RAND_2397 = {2{`RANDOM}};
  T_38110_1_exc_cause = _RAND_2397[63:0];
  _RAND_2398 = {1{`RANDOM}};
  T_38110_1_bypassable = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  T_38110_1_mem_cmd = _RAND_2399[3:0];
  _RAND_2400 = {1{`RANDOM}};
  T_38110_1_mem_typ = _RAND_2400[2:0];
  _RAND_2401 = {1{`RANDOM}};
  T_38110_1_is_fence = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  T_38110_1_is_fencei = _RAND_2402[0:0];
  _RAND_2403 = {1{`RANDOM}};
  T_38110_1_is_store = _RAND_2403[0:0];
  _RAND_2404 = {1{`RANDOM}};
  T_38110_1_is_amo = _RAND_2404[0:0];
  _RAND_2405 = {1{`RANDOM}};
  T_38110_1_is_load = _RAND_2405[0:0];
  _RAND_2406 = {1{`RANDOM}};
  T_38110_1_is_unique = _RAND_2406[0:0];
  _RAND_2407 = {1{`RANDOM}};
  T_38110_1_flush_on_commit = _RAND_2407[0:0];
  _RAND_2408 = {1{`RANDOM}};
  T_38110_1_ldst = _RAND_2408[5:0];
  _RAND_2409 = {1{`RANDOM}};
  T_38110_1_lrs1 = _RAND_2409[5:0];
  _RAND_2410 = {1{`RANDOM}};
  T_38110_1_lrs2 = _RAND_2410[5:0];
  _RAND_2411 = {1{`RANDOM}};
  T_38110_1_lrs3 = _RAND_2411[5:0];
  _RAND_2412 = {1{`RANDOM}};
  T_38110_1_ldst_val = _RAND_2412[0:0];
  _RAND_2413 = {1{`RANDOM}};
  T_38110_1_dst_rtype = _RAND_2413[1:0];
  _RAND_2414 = {1{`RANDOM}};
  T_38110_1_lrs1_rtype = _RAND_2414[1:0];
  _RAND_2415 = {1{`RANDOM}};
  T_38110_1_lrs2_rtype = _RAND_2415[1:0];
  _RAND_2416 = {1{`RANDOM}};
  T_38110_1_frs3_en = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  T_38110_1_fp_val = _RAND_2417[0:0];
  _RAND_2418 = {1{`RANDOM}};
  T_38110_1_fp_single = _RAND_2418[0:0];
  _RAND_2419 = {1{`RANDOM}};
  T_38110_1_xcpt_if = _RAND_2419[0:0];
  _RAND_2420 = {1{`RANDOM}};
  T_38110_1_replay_if = _RAND_2420[0:0];
  _RAND_2421 = {2{`RANDOM}};
  T_38110_1_debug_wdata = _RAND_2421[63:0];
  _RAND_2422 = {1{`RANDOM}};
  T_38110_1_debug_events_fetch_seq = _RAND_2422[31:0];
  _RAND_2423 = {1{`RANDOM}};
  T_38110_2_valid = _RAND_2423[0:0];
  _RAND_2424 = {1{`RANDOM}};
  T_38110_2_iw_state = _RAND_2424[1:0];
  _RAND_2425 = {1{`RANDOM}};
  T_38110_2_uopc = _RAND_2425[8:0];
  _RAND_2426 = {1{`RANDOM}};
  T_38110_2_inst = _RAND_2426[31:0];
  _RAND_2427 = {2{`RANDOM}};
  T_38110_2_pc = _RAND_2427[39:0];
  _RAND_2428 = {1{`RANDOM}};
  T_38110_2_fu_code = _RAND_2428[7:0];
  _RAND_2429 = {1{`RANDOM}};
  T_38110_2_ctrl_br_type = _RAND_2429[3:0];
  _RAND_2430 = {1{`RANDOM}};
  T_38110_2_ctrl_op1_sel = _RAND_2430[1:0];
  _RAND_2431 = {1{`RANDOM}};
  T_38110_2_ctrl_op2_sel = _RAND_2431[2:0];
  _RAND_2432 = {1{`RANDOM}};
  T_38110_2_ctrl_imm_sel = _RAND_2432[2:0];
  _RAND_2433 = {1{`RANDOM}};
  T_38110_2_ctrl_op_fcn = _RAND_2433[3:0];
  _RAND_2434 = {1{`RANDOM}};
  T_38110_2_ctrl_fcn_dw = _RAND_2434[0:0];
  _RAND_2435 = {1{`RANDOM}};
  T_38110_2_ctrl_rf_wen = _RAND_2435[0:0];
  _RAND_2436 = {1{`RANDOM}};
  T_38110_2_ctrl_csr_cmd = _RAND_2436[2:0];
  _RAND_2437 = {1{`RANDOM}};
  T_38110_2_ctrl_is_load = _RAND_2437[0:0];
  _RAND_2438 = {1{`RANDOM}};
  T_38110_2_ctrl_is_sta = _RAND_2438[0:0];
  _RAND_2439 = {1{`RANDOM}};
  T_38110_2_ctrl_is_std = _RAND_2439[0:0];
  _RAND_2440 = {1{`RANDOM}};
  T_38110_2_wakeup_delay = _RAND_2440[1:0];
  _RAND_2441 = {1{`RANDOM}};
  T_38110_2_allocate_brtag = _RAND_2441[0:0];
  _RAND_2442 = {1{`RANDOM}};
  T_38110_2_is_br_or_jmp = _RAND_2442[0:0];
  _RAND_2443 = {1{`RANDOM}};
  T_38110_2_is_jump = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  T_38110_2_is_jal = _RAND_2444[0:0];
  _RAND_2445 = {1{`RANDOM}};
  T_38110_2_is_ret = _RAND_2445[0:0];
  _RAND_2446 = {1{`RANDOM}};
  T_38110_2_is_call = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  T_38110_2_br_mask = _RAND_2447[7:0];
  _RAND_2448 = {1{`RANDOM}};
  T_38110_2_br_tag = _RAND_2448[2:0];
  _RAND_2449 = {1{`RANDOM}};
  T_38110_2_br_prediction_bpd_predict_val = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  T_38110_2_br_prediction_bpd_predict_taken = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  T_38110_2_br_prediction_btb_hit = _RAND_2451[0:0];
  _RAND_2452 = {1{`RANDOM}};
  T_38110_2_br_prediction_btb_predicted = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  T_38110_2_br_prediction_is_br_or_jalr = _RAND_2453[0:0];
  _RAND_2454 = {1{`RANDOM}};
  T_38110_2_stat_brjmp_mispredicted = _RAND_2454[0:0];
  _RAND_2455 = {1{`RANDOM}};
  T_38110_2_stat_btb_made_pred = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  T_38110_2_stat_btb_mispredicted = _RAND_2456[0:0];
  _RAND_2457 = {1{`RANDOM}};
  T_38110_2_stat_bpd_made_pred = _RAND_2457[0:0];
  _RAND_2458 = {1{`RANDOM}};
  T_38110_2_stat_bpd_mispredicted = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  T_38110_2_fetch_pc_lob = _RAND_2459[2:0];
  _RAND_2460 = {1{`RANDOM}};
  T_38110_2_imm_packed = _RAND_2460[19:0];
  _RAND_2461 = {1{`RANDOM}};
  T_38110_2_csr_addr = _RAND_2461[11:0];
  _RAND_2462 = {1{`RANDOM}};
  T_38110_2_rob_idx = _RAND_2462[5:0];
  _RAND_2463 = {1{`RANDOM}};
  T_38110_2_ldq_idx = _RAND_2463[3:0];
  _RAND_2464 = {1{`RANDOM}};
  T_38110_2_stq_idx = _RAND_2464[3:0];
  _RAND_2465 = {1{`RANDOM}};
  T_38110_2_brob_idx = _RAND_2465[4:0];
  _RAND_2466 = {1{`RANDOM}};
  T_38110_2_pdst = _RAND_2466[6:0];
  _RAND_2467 = {1{`RANDOM}};
  T_38110_2_pop1 = _RAND_2467[6:0];
  _RAND_2468 = {1{`RANDOM}};
  T_38110_2_pop2 = _RAND_2468[6:0];
  _RAND_2469 = {1{`RANDOM}};
  T_38110_2_pop3 = _RAND_2469[6:0];
  _RAND_2470 = {1{`RANDOM}};
  T_38110_2_prs1_busy = _RAND_2470[0:0];
  _RAND_2471 = {1{`RANDOM}};
  T_38110_2_prs2_busy = _RAND_2471[0:0];
  _RAND_2472 = {1{`RANDOM}};
  T_38110_2_prs3_busy = _RAND_2472[0:0];
  _RAND_2473 = {1{`RANDOM}};
  T_38110_2_stale_pdst = _RAND_2473[6:0];
  _RAND_2474 = {1{`RANDOM}};
  T_38110_2_exception = _RAND_2474[0:0];
  _RAND_2475 = {2{`RANDOM}};
  T_38110_2_exc_cause = _RAND_2475[63:0];
  _RAND_2476 = {1{`RANDOM}};
  T_38110_2_bypassable = _RAND_2476[0:0];
  _RAND_2477 = {1{`RANDOM}};
  T_38110_2_mem_cmd = _RAND_2477[3:0];
  _RAND_2478 = {1{`RANDOM}};
  T_38110_2_mem_typ = _RAND_2478[2:0];
  _RAND_2479 = {1{`RANDOM}};
  T_38110_2_is_fence = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  T_38110_2_is_fencei = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  T_38110_2_is_store = _RAND_2481[0:0];
  _RAND_2482 = {1{`RANDOM}};
  T_38110_2_is_amo = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  T_38110_2_is_load = _RAND_2483[0:0];
  _RAND_2484 = {1{`RANDOM}};
  T_38110_2_is_unique = _RAND_2484[0:0];
  _RAND_2485 = {1{`RANDOM}};
  T_38110_2_flush_on_commit = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  T_38110_2_ldst = _RAND_2486[5:0];
  _RAND_2487 = {1{`RANDOM}};
  T_38110_2_lrs1 = _RAND_2487[5:0];
  _RAND_2488 = {1{`RANDOM}};
  T_38110_2_lrs2 = _RAND_2488[5:0];
  _RAND_2489 = {1{`RANDOM}};
  T_38110_2_lrs3 = _RAND_2489[5:0];
  _RAND_2490 = {1{`RANDOM}};
  T_38110_2_ldst_val = _RAND_2490[0:0];
  _RAND_2491 = {1{`RANDOM}};
  T_38110_2_dst_rtype = _RAND_2491[1:0];
  _RAND_2492 = {1{`RANDOM}};
  T_38110_2_lrs1_rtype = _RAND_2492[1:0];
  _RAND_2493 = {1{`RANDOM}};
  T_38110_2_lrs2_rtype = _RAND_2493[1:0];
  _RAND_2494 = {1{`RANDOM}};
  T_38110_2_frs3_en = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  T_38110_2_fp_val = _RAND_2495[0:0];
  _RAND_2496 = {1{`RANDOM}};
  T_38110_2_fp_single = _RAND_2496[0:0];
  _RAND_2497 = {1{`RANDOM}};
  T_38110_2_xcpt_if = _RAND_2497[0:0];
  _RAND_2498 = {1{`RANDOM}};
  T_38110_2_replay_if = _RAND_2498[0:0];
  _RAND_2499 = {2{`RANDOM}};
  T_38110_2_debug_wdata = _RAND_2499[63:0];
  _RAND_2500 = {1{`RANDOM}};
  T_38110_2_debug_events_fetch_seq = _RAND_2500[31:0];
  _RAND_2501 = {1{`RANDOM}};
  T_38110_3_valid = _RAND_2501[0:0];
  _RAND_2502 = {1{`RANDOM}};
  T_38110_3_iw_state = _RAND_2502[1:0];
  _RAND_2503 = {1{`RANDOM}};
  T_38110_3_uopc = _RAND_2503[8:0];
  _RAND_2504 = {1{`RANDOM}};
  T_38110_3_inst = _RAND_2504[31:0];
  _RAND_2505 = {2{`RANDOM}};
  T_38110_3_pc = _RAND_2505[39:0];
  _RAND_2506 = {1{`RANDOM}};
  T_38110_3_fu_code = _RAND_2506[7:0];
  _RAND_2507 = {1{`RANDOM}};
  T_38110_3_ctrl_br_type = _RAND_2507[3:0];
  _RAND_2508 = {1{`RANDOM}};
  T_38110_3_ctrl_op1_sel = _RAND_2508[1:0];
  _RAND_2509 = {1{`RANDOM}};
  T_38110_3_ctrl_op2_sel = _RAND_2509[2:0];
  _RAND_2510 = {1{`RANDOM}};
  T_38110_3_ctrl_imm_sel = _RAND_2510[2:0];
  _RAND_2511 = {1{`RANDOM}};
  T_38110_3_ctrl_op_fcn = _RAND_2511[3:0];
  _RAND_2512 = {1{`RANDOM}};
  T_38110_3_ctrl_fcn_dw = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  T_38110_3_ctrl_rf_wen = _RAND_2513[0:0];
  _RAND_2514 = {1{`RANDOM}};
  T_38110_3_ctrl_csr_cmd = _RAND_2514[2:0];
  _RAND_2515 = {1{`RANDOM}};
  T_38110_3_ctrl_is_load = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  T_38110_3_ctrl_is_sta = _RAND_2516[0:0];
  _RAND_2517 = {1{`RANDOM}};
  T_38110_3_ctrl_is_std = _RAND_2517[0:0];
  _RAND_2518 = {1{`RANDOM}};
  T_38110_3_wakeup_delay = _RAND_2518[1:0];
  _RAND_2519 = {1{`RANDOM}};
  T_38110_3_allocate_brtag = _RAND_2519[0:0];
  _RAND_2520 = {1{`RANDOM}};
  T_38110_3_is_br_or_jmp = _RAND_2520[0:0];
  _RAND_2521 = {1{`RANDOM}};
  T_38110_3_is_jump = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  T_38110_3_is_jal = _RAND_2522[0:0];
  _RAND_2523 = {1{`RANDOM}};
  T_38110_3_is_ret = _RAND_2523[0:0];
  _RAND_2524 = {1{`RANDOM}};
  T_38110_3_is_call = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  T_38110_3_br_mask = _RAND_2525[7:0];
  _RAND_2526 = {1{`RANDOM}};
  T_38110_3_br_tag = _RAND_2526[2:0];
  _RAND_2527 = {1{`RANDOM}};
  T_38110_3_br_prediction_bpd_predict_val = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  T_38110_3_br_prediction_bpd_predict_taken = _RAND_2528[0:0];
  _RAND_2529 = {1{`RANDOM}};
  T_38110_3_br_prediction_btb_hit = _RAND_2529[0:0];
  _RAND_2530 = {1{`RANDOM}};
  T_38110_3_br_prediction_btb_predicted = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  T_38110_3_br_prediction_is_br_or_jalr = _RAND_2531[0:0];
  _RAND_2532 = {1{`RANDOM}};
  T_38110_3_stat_brjmp_mispredicted = _RAND_2532[0:0];
  _RAND_2533 = {1{`RANDOM}};
  T_38110_3_stat_btb_made_pred = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  T_38110_3_stat_btb_mispredicted = _RAND_2534[0:0];
  _RAND_2535 = {1{`RANDOM}};
  T_38110_3_stat_bpd_made_pred = _RAND_2535[0:0];
  _RAND_2536 = {1{`RANDOM}};
  T_38110_3_stat_bpd_mispredicted = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  T_38110_3_fetch_pc_lob = _RAND_2537[2:0];
  _RAND_2538 = {1{`RANDOM}};
  T_38110_3_imm_packed = _RAND_2538[19:0];
  _RAND_2539 = {1{`RANDOM}};
  T_38110_3_csr_addr = _RAND_2539[11:0];
  _RAND_2540 = {1{`RANDOM}};
  T_38110_3_rob_idx = _RAND_2540[5:0];
  _RAND_2541 = {1{`RANDOM}};
  T_38110_3_ldq_idx = _RAND_2541[3:0];
  _RAND_2542 = {1{`RANDOM}};
  T_38110_3_stq_idx = _RAND_2542[3:0];
  _RAND_2543 = {1{`RANDOM}};
  T_38110_3_brob_idx = _RAND_2543[4:0];
  _RAND_2544 = {1{`RANDOM}};
  T_38110_3_pdst = _RAND_2544[6:0];
  _RAND_2545 = {1{`RANDOM}};
  T_38110_3_pop1 = _RAND_2545[6:0];
  _RAND_2546 = {1{`RANDOM}};
  T_38110_3_pop2 = _RAND_2546[6:0];
  _RAND_2547 = {1{`RANDOM}};
  T_38110_3_pop3 = _RAND_2547[6:0];
  _RAND_2548 = {1{`RANDOM}};
  T_38110_3_prs1_busy = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  T_38110_3_prs2_busy = _RAND_2549[0:0];
  _RAND_2550 = {1{`RANDOM}};
  T_38110_3_prs3_busy = _RAND_2550[0:0];
  _RAND_2551 = {1{`RANDOM}};
  T_38110_3_stale_pdst = _RAND_2551[6:0];
  _RAND_2552 = {1{`RANDOM}};
  T_38110_3_exception = _RAND_2552[0:0];
  _RAND_2553 = {2{`RANDOM}};
  T_38110_3_exc_cause = _RAND_2553[63:0];
  _RAND_2554 = {1{`RANDOM}};
  T_38110_3_bypassable = _RAND_2554[0:0];
  _RAND_2555 = {1{`RANDOM}};
  T_38110_3_mem_cmd = _RAND_2555[3:0];
  _RAND_2556 = {1{`RANDOM}};
  T_38110_3_mem_typ = _RAND_2556[2:0];
  _RAND_2557 = {1{`RANDOM}};
  T_38110_3_is_fence = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  T_38110_3_is_fencei = _RAND_2558[0:0];
  _RAND_2559 = {1{`RANDOM}};
  T_38110_3_is_store = _RAND_2559[0:0];
  _RAND_2560 = {1{`RANDOM}};
  T_38110_3_is_amo = _RAND_2560[0:0];
  _RAND_2561 = {1{`RANDOM}};
  T_38110_3_is_load = _RAND_2561[0:0];
  _RAND_2562 = {1{`RANDOM}};
  T_38110_3_is_unique = _RAND_2562[0:0];
  _RAND_2563 = {1{`RANDOM}};
  T_38110_3_flush_on_commit = _RAND_2563[0:0];
  _RAND_2564 = {1{`RANDOM}};
  T_38110_3_ldst = _RAND_2564[5:0];
  _RAND_2565 = {1{`RANDOM}};
  T_38110_3_lrs1 = _RAND_2565[5:0];
  _RAND_2566 = {1{`RANDOM}};
  T_38110_3_lrs2 = _RAND_2566[5:0];
  _RAND_2567 = {1{`RANDOM}};
  T_38110_3_lrs3 = _RAND_2567[5:0];
  _RAND_2568 = {1{`RANDOM}};
  T_38110_3_ldst_val = _RAND_2568[0:0];
  _RAND_2569 = {1{`RANDOM}};
  T_38110_3_dst_rtype = _RAND_2569[1:0];
  _RAND_2570 = {1{`RANDOM}};
  T_38110_3_lrs1_rtype = _RAND_2570[1:0];
  _RAND_2571 = {1{`RANDOM}};
  T_38110_3_lrs2_rtype = _RAND_2571[1:0];
  _RAND_2572 = {1{`RANDOM}};
  T_38110_3_frs3_en = _RAND_2572[0:0];
  _RAND_2573 = {1{`RANDOM}};
  T_38110_3_fp_val = _RAND_2573[0:0];
  _RAND_2574 = {1{`RANDOM}};
  T_38110_3_fp_single = _RAND_2574[0:0];
  _RAND_2575 = {1{`RANDOM}};
  T_38110_3_xcpt_if = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  T_38110_3_replay_if = _RAND_2576[0:0];
  _RAND_2577 = {2{`RANDOM}};
  T_38110_3_debug_wdata = _RAND_2577[63:0];
  _RAND_2578 = {1{`RANDOM}};
  T_38110_3_debug_events_fetch_seq = _RAND_2578[31:0];
  _RAND_2579 = {1{`RANDOM}};
  T_38110_4_valid = _RAND_2579[0:0];
  _RAND_2580 = {1{`RANDOM}};
  T_38110_4_iw_state = _RAND_2580[1:0];
  _RAND_2581 = {1{`RANDOM}};
  T_38110_4_uopc = _RAND_2581[8:0];
  _RAND_2582 = {1{`RANDOM}};
  T_38110_4_inst = _RAND_2582[31:0];
  _RAND_2583 = {2{`RANDOM}};
  T_38110_4_pc = _RAND_2583[39:0];
  _RAND_2584 = {1{`RANDOM}};
  T_38110_4_fu_code = _RAND_2584[7:0];
  _RAND_2585 = {1{`RANDOM}};
  T_38110_4_ctrl_br_type = _RAND_2585[3:0];
  _RAND_2586 = {1{`RANDOM}};
  T_38110_4_ctrl_op1_sel = _RAND_2586[1:0];
  _RAND_2587 = {1{`RANDOM}};
  T_38110_4_ctrl_op2_sel = _RAND_2587[2:0];
  _RAND_2588 = {1{`RANDOM}};
  T_38110_4_ctrl_imm_sel = _RAND_2588[2:0];
  _RAND_2589 = {1{`RANDOM}};
  T_38110_4_ctrl_op_fcn = _RAND_2589[3:0];
  _RAND_2590 = {1{`RANDOM}};
  T_38110_4_ctrl_fcn_dw = _RAND_2590[0:0];
  _RAND_2591 = {1{`RANDOM}};
  T_38110_4_ctrl_rf_wen = _RAND_2591[0:0];
  _RAND_2592 = {1{`RANDOM}};
  T_38110_4_ctrl_csr_cmd = _RAND_2592[2:0];
  _RAND_2593 = {1{`RANDOM}};
  T_38110_4_ctrl_is_load = _RAND_2593[0:0];
  _RAND_2594 = {1{`RANDOM}};
  T_38110_4_ctrl_is_sta = _RAND_2594[0:0];
  _RAND_2595 = {1{`RANDOM}};
  T_38110_4_ctrl_is_std = _RAND_2595[0:0];
  _RAND_2596 = {1{`RANDOM}};
  T_38110_4_wakeup_delay = _RAND_2596[1:0];
  _RAND_2597 = {1{`RANDOM}};
  T_38110_4_allocate_brtag = _RAND_2597[0:0];
  _RAND_2598 = {1{`RANDOM}};
  T_38110_4_is_br_or_jmp = _RAND_2598[0:0];
  _RAND_2599 = {1{`RANDOM}};
  T_38110_4_is_jump = _RAND_2599[0:0];
  _RAND_2600 = {1{`RANDOM}};
  T_38110_4_is_jal = _RAND_2600[0:0];
  _RAND_2601 = {1{`RANDOM}};
  T_38110_4_is_ret = _RAND_2601[0:0];
  _RAND_2602 = {1{`RANDOM}};
  T_38110_4_is_call = _RAND_2602[0:0];
  _RAND_2603 = {1{`RANDOM}};
  T_38110_4_br_mask = _RAND_2603[7:0];
  _RAND_2604 = {1{`RANDOM}};
  T_38110_4_br_tag = _RAND_2604[2:0];
  _RAND_2605 = {1{`RANDOM}};
  T_38110_4_br_prediction_bpd_predict_val = _RAND_2605[0:0];
  _RAND_2606 = {1{`RANDOM}};
  T_38110_4_br_prediction_bpd_predict_taken = _RAND_2606[0:0];
  _RAND_2607 = {1{`RANDOM}};
  T_38110_4_br_prediction_btb_hit = _RAND_2607[0:0];
  _RAND_2608 = {1{`RANDOM}};
  T_38110_4_br_prediction_btb_predicted = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  T_38110_4_br_prediction_is_br_or_jalr = _RAND_2609[0:0];
  _RAND_2610 = {1{`RANDOM}};
  T_38110_4_stat_brjmp_mispredicted = _RAND_2610[0:0];
  _RAND_2611 = {1{`RANDOM}};
  T_38110_4_stat_btb_made_pred = _RAND_2611[0:0];
  _RAND_2612 = {1{`RANDOM}};
  T_38110_4_stat_btb_mispredicted = _RAND_2612[0:0];
  _RAND_2613 = {1{`RANDOM}};
  T_38110_4_stat_bpd_made_pred = _RAND_2613[0:0];
  _RAND_2614 = {1{`RANDOM}};
  T_38110_4_stat_bpd_mispredicted = _RAND_2614[0:0];
  _RAND_2615 = {1{`RANDOM}};
  T_38110_4_fetch_pc_lob = _RAND_2615[2:0];
  _RAND_2616 = {1{`RANDOM}};
  T_38110_4_imm_packed = _RAND_2616[19:0];
  _RAND_2617 = {1{`RANDOM}};
  T_38110_4_csr_addr = _RAND_2617[11:0];
  _RAND_2618 = {1{`RANDOM}};
  T_38110_4_rob_idx = _RAND_2618[5:0];
  _RAND_2619 = {1{`RANDOM}};
  T_38110_4_ldq_idx = _RAND_2619[3:0];
  _RAND_2620 = {1{`RANDOM}};
  T_38110_4_stq_idx = _RAND_2620[3:0];
  _RAND_2621 = {1{`RANDOM}};
  T_38110_4_brob_idx = _RAND_2621[4:0];
  _RAND_2622 = {1{`RANDOM}};
  T_38110_4_pdst = _RAND_2622[6:0];
  _RAND_2623 = {1{`RANDOM}};
  T_38110_4_pop1 = _RAND_2623[6:0];
  _RAND_2624 = {1{`RANDOM}};
  T_38110_4_pop2 = _RAND_2624[6:0];
  _RAND_2625 = {1{`RANDOM}};
  T_38110_4_pop3 = _RAND_2625[6:0];
  _RAND_2626 = {1{`RANDOM}};
  T_38110_4_prs1_busy = _RAND_2626[0:0];
  _RAND_2627 = {1{`RANDOM}};
  T_38110_4_prs2_busy = _RAND_2627[0:0];
  _RAND_2628 = {1{`RANDOM}};
  T_38110_4_prs3_busy = _RAND_2628[0:0];
  _RAND_2629 = {1{`RANDOM}};
  T_38110_4_stale_pdst = _RAND_2629[6:0];
  _RAND_2630 = {1{`RANDOM}};
  T_38110_4_exception = _RAND_2630[0:0];
  _RAND_2631 = {2{`RANDOM}};
  T_38110_4_exc_cause = _RAND_2631[63:0];
  _RAND_2632 = {1{`RANDOM}};
  T_38110_4_bypassable = _RAND_2632[0:0];
  _RAND_2633 = {1{`RANDOM}};
  T_38110_4_mem_cmd = _RAND_2633[3:0];
  _RAND_2634 = {1{`RANDOM}};
  T_38110_4_mem_typ = _RAND_2634[2:0];
  _RAND_2635 = {1{`RANDOM}};
  T_38110_4_is_fence = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  T_38110_4_is_fencei = _RAND_2636[0:0];
  _RAND_2637 = {1{`RANDOM}};
  T_38110_4_is_store = _RAND_2637[0:0];
  _RAND_2638 = {1{`RANDOM}};
  T_38110_4_is_amo = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  T_38110_4_is_load = _RAND_2639[0:0];
  _RAND_2640 = {1{`RANDOM}};
  T_38110_4_is_unique = _RAND_2640[0:0];
  _RAND_2641 = {1{`RANDOM}};
  T_38110_4_flush_on_commit = _RAND_2641[0:0];
  _RAND_2642 = {1{`RANDOM}};
  T_38110_4_ldst = _RAND_2642[5:0];
  _RAND_2643 = {1{`RANDOM}};
  T_38110_4_lrs1 = _RAND_2643[5:0];
  _RAND_2644 = {1{`RANDOM}};
  T_38110_4_lrs2 = _RAND_2644[5:0];
  _RAND_2645 = {1{`RANDOM}};
  T_38110_4_lrs3 = _RAND_2645[5:0];
  _RAND_2646 = {1{`RANDOM}};
  T_38110_4_ldst_val = _RAND_2646[0:0];
  _RAND_2647 = {1{`RANDOM}};
  T_38110_4_dst_rtype = _RAND_2647[1:0];
  _RAND_2648 = {1{`RANDOM}};
  T_38110_4_lrs1_rtype = _RAND_2648[1:0];
  _RAND_2649 = {1{`RANDOM}};
  T_38110_4_lrs2_rtype = _RAND_2649[1:0];
  _RAND_2650 = {1{`RANDOM}};
  T_38110_4_frs3_en = _RAND_2650[0:0];
  _RAND_2651 = {1{`RANDOM}};
  T_38110_4_fp_val = _RAND_2651[0:0];
  _RAND_2652 = {1{`RANDOM}};
  T_38110_4_fp_single = _RAND_2652[0:0];
  _RAND_2653 = {1{`RANDOM}};
  T_38110_4_xcpt_if = _RAND_2653[0:0];
  _RAND_2654 = {1{`RANDOM}};
  T_38110_4_replay_if = _RAND_2654[0:0];
  _RAND_2655 = {2{`RANDOM}};
  T_38110_4_debug_wdata = _RAND_2655[63:0];
  _RAND_2656 = {1{`RANDOM}};
  T_38110_4_debug_events_fetch_seq = _RAND_2656[31:0];
  _RAND_2657 = {1{`RANDOM}};
  T_38110_5_valid = _RAND_2657[0:0];
  _RAND_2658 = {1{`RANDOM}};
  T_38110_5_iw_state = _RAND_2658[1:0];
  _RAND_2659 = {1{`RANDOM}};
  T_38110_5_uopc = _RAND_2659[8:0];
  _RAND_2660 = {1{`RANDOM}};
  T_38110_5_inst = _RAND_2660[31:0];
  _RAND_2661 = {2{`RANDOM}};
  T_38110_5_pc = _RAND_2661[39:0];
  _RAND_2662 = {1{`RANDOM}};
  T_38110_5_fu_code = _RAND_2662[7:0];
  _RAND_2663 = {1{`RANDOM}};
  T_38110_5_ctrl_br_type = _RAND_2663[3:0];
  _RAND_2664 = {1{`RANDOM}};
  T_38110_5_ctrl_op1_sel = _RAND_2664[1:0];
  _RAND_2665 = {1{`RANDOM}};
  T_38110_5_ctrl_op2_sel = _RAND_2665[2:0];
  _RAND_2666 = {1{`RANDOM}};
  T_38110_5_ctrl_imm_sel = _RAND_2666[2:0];
  _RAND_2667 = {1{`RANDOM}};
  T_38110_5_ctrl_op_fcn = _RAND_2667[3:0];
  _RAND_2668 = {1{`RANDOM}};
  T_38110_5_ctrl_fcn_dw = _RAND_2668[0:0];
  _RAND_2669 = {1{`RANDOM}};
  T_38110_5_ctrl_rf_wen = _RAND_2669[0:0];
  _RAND_2670 = {1{`RANDOM}};
  T_38110_5_ctrl_csr_cmd = _RAND_2670[2:0];
  _RAND_2671 = {1{`RANDOM}};
  T_38110_5_ctrl_is_load = _RAND_2671[0:0];
  _RAND_2672 = {1{`RANDOM}};
  T_38110_5_ctrl_is_sta = _RAND_2672[0:0];
  _RAND_2673 = {1{`RANDOM}};
  T_38110_5_ctrl_is_std = _RAND_2673[0:0];
  _RAND_2674 = {1{`RANDOM}};
  T_38110_5_wakeup_delay = _RAND_2674[1:0];
  _RAND_2675 = {1{`RANDOM}};
  T_38110_5_allocate_brtag = _RAND_2675[0:0];
  _RAND_2676 = {1{`RANDOM}};
  T_38110_5_is_br_or_jmp = _RAND_2676[0:0];
  _RAND_2677 = {1{`RANDOM}};
  T_38110_5_is_jump = _RAND_2677[0:0];
  _RAND_2678 = {1{`RANDOM}};
  T_38110_5_is_jal = _RAND_2678[0:0];
  _RAND_2679 = {1{`RANDOM}};
  T_38110_5_is_ret = _RAND_2679[0:0];
  _RAND_2680 = {1{`RANDOM}};
  T_38110_5_is_call = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  T_38110_5_br_mask = _RAND_2681[7:0];
  _RAND_2682 = {1{`RANDOM}};
  T_38110_5_br_tag = _RAND_2682[2:0];
  _RAND_2683 = {1{`RANDOM}};
  T_38110_5_br_prediction_bpd_predict_val = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  T_38110_5_br_prediction_bpd_predict_taken = _RAND_2684[0:0];
  _RAND_2685 = {1{`RANDOM}};
  T_38110_5_br_prediction_btb_hit = _RAND_2685[0:0];
  _RAND_2686 = {1{`RANDOM}};
  T_38110_5_br_prediction_btb_predicted = _RAND_2686[0:0];
  _RAND_2687 = {1{`RANDOM}};
  T_38110_5_br_prediction_is_br_or_jalr = _RAND_2687[0:0];
  _RAND_2688 = {1{`RANDOM}};
  T_38110_5_stat_brjmp_mispredicted = _RAND_2688[0:0];
  _RAND_2689 = {1{`RANDOM}};
  T_38110_5_stat_btb_made_pred = _RAND_2689[0:0];
  _RAND_2690 = {1{`RANDOM}};
  T_38110_5_stat_btb_mispredicted = _RAND_2690[0:0];
  _RAND_2691 = {1{`RANDOM}};
  T_38110_5_stat_bpd_made_pred = _RAND_2691[0:0];
  _RAND_2692 = {1{`RANDOM}};
  T_38110_5_stat_bpd_mispredicted = _RAND_2692[0:0];
  _RAND_2693 = {1{`RANDOM}};
  T_38110_5_fetch_pc_lob = _RAND_2693[2:0];
  _RAND_2694 = {1{`RANDOM}};
  T_38110_5_imm_packed = _RAND_2694[19:0];
  _RAND_2695 = {1{`RANDOM}};
  T_38110_5_csr_addr = _RAND_2695[11:0];
  _RAND_2696 = {1{`RANDOM}};
  T_38110_5_rob_idx = _RAND_2696[5:0];
  _RAND_2697 = {1{`RANDOM}};
  T_38110_5_ldq_idx = _RAND_2697[3:0];
  _RAND_2698 = {1{`RANDOM}};
  T_38110_5_stq_idx = _RAND_2698[3:0];
  _RAND_2699 = {1{`RANDOM}};
  T_38110_5_brob_idx = _RAND_2699[4:0];
  _RAND_2700 = {1{`RANDOM}};
  T_38110_5_pdst = _RAND_2700[6:0];
  _RAND_2701 = {1{`RANDOM}};
  T_38110_5_pop1 = _RAND_2701[6:0];
  _RAND_2702 = {1{`RANDOM}};
  T_38110_5_pop2 = _RAND_2702[6:0];
  _RAND_2703 = {1{`RANDOM}};
  T_38110_5_pop3 = _RAND_2703[6:0];
  _RAND_2704 = {1{`RANDOM}};
  T_38110_5_prs1_busy = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  T_38110_5_prs2_busy = _RAND_2705[0:0];
  _RAND_2706 = {1{`RANDOM}};
  T_38110_5_prs3_busy = _RAND_2706[0:0];
  _RAND_2707 = {1{`RANDOM}};
  T_38110_5_stale_pdst = _RAND_2707[6:0];
  _RAND_2708 = {1{`RANDOM}};
  T_38110_5_exception = _RAND_2708[0:0];
  _RAND_2709 = {2{`RANDOM}};
  T_38110_5_exc_cause = _RAND_2709[63:0];
  _RAND_2710 = {1{`RANDOM}};
  T_38110_5_bypassable = _RAND_2710[0:0];
  _RAND_2711 = {1{`RANDOM}};
  T_38110_5_mem_cmd = _RAND_2711[3:0];
  _RAND_2712 = {1{`RANDOM}};
  T_38110_5_mem_typ = _RAND_2712[2:0];
  _RAND_2713 = {1{`RANDOM}};
  T_38110_5_is_fence = _RAND_2713[0:0];
  _RAND_2714 = {1{`RANDOM}};
  T_38110_5_is_fencei = _RAND_2714[0:0];
  _RAND_2715 = {1{`RANDOM}};
  T_38110_5_is_store = _RAND_2715[0:0];
  _RAND_2716 = {1{`RANDOM}};
  T_38110_5_is_amo = _RAND_2716[0:0];
  _RAND_2717 = {1{`RANDOM}};
  T_38110_5_is_load = _RAND_2717[0:0];
  _RAND_2718 = {1{`RANDOM}};
  T_38110_5_is_unique = _RAND_2718[0:0];
  _RAND_2719 = {1{`RANDOM}};
  T_38110_5_flush_on_commit = _RAND_2719[0:0];
  _RAND_2720 = {1{`RANDOM}};
  T_38110_5_ldst = _RAND_2720[5:0];
  _RAND_2721 = {1{`RANDOM}};
  T_38110_5_lrs1 = _RAND_2721[5:0];
  _RAND_2722 = {1{`RANDOM}};
  T_38110_5_lrs2 = _RAND_2722[5:0];
  _RAND_2723 = {1{`RANDOM}};
  T_38110_5_lrs3 = _RAND_2723[5:0];
  _RAND_2724 = {1{`RANDOM}};
  T_38110_5_ldst_val = _RAND_2724[0:0];
  _RAND_2725 = {1{`RANDOM}};
  T_38110_5_dst_rtype = _RAND_2725[1:0];
  _RAND_2726 = {1{`RANDOM}};
  T_38110_5_lrs1_rtype = _RAND_2726[1:0];
  _RAND_2727 = {1{`RANDOM}};
  T_38110_5_lrs2_rtype = _RAND_2727[1:0];
  _RAND_2728 = {1{`RANDOM}};
  T_38110_5_frs3_en = _RAND_2728[0:0];
  _RAND_2729 = {1{`RANDOM}};
  T_38110_5_fp_val = _RAND_2729[0:0];
  _RAND_2730 = {1{`RANDOM}};
  T_38110_5_fp_single = _RAND_2730[0:0];
  _RAND_2731 = {1{`RANDOM}};
  T_38110_5_xcpt_if = _RAND_2731[0:0];
  _RAND_2732 = {1{`RANDOM}};
  T_38110_5_replay_if = _RAND_2732[0:0];
  _RAND_2733 = {2{`RANDOM}};
  T_38110_5_debug_wdata = _RAND_2733[63:0];
  _RAND_2734 = {1{`RANDOM}};
  T_38110_5_debug_events_fetch_seq = _RAND_2734[31:0];
  _RAND_2735 = {1{`RANDOM}};
  T_38110_6_valid = _RAND_2735[0:0];
  _RAND_2736 = {1{`RANDOM}};
  T_38110_6_iw_state = _RAND_2736[1:0];
  _RAND_2737 = {1{`RANDOM}};
  T_38110_6_uopc = _RAND_2737[8:0];
  _RAND_2738 = {1{`RANDOM}};
  T_38110_6_inst = _RAND_2738[31:0];
  _RAND_2739 = {2{`RANDOM}};
  T_38110_6_pc = _RAND_2739[39:0];
  _RAND_2740 = {1{`RANDOM}};
  T_38110_6_fu_code = _RAND_2740[7:0];
  _RAND_2741 = {1{`RANDOM}};
  T_38110_6_ctrl_br_type = _RAND_2741[3:0];
  _RAND_2742 = {1{`RANDOM}};
  T_38110_6_ctrl_op1_sel = _RAND_2742[1:0];
  _RAND_2743 = {1{`RANDOM}};
  T_38110_6_ctrl_op2_sel = _RAND_2743[2:0];
  _RAND_2744 = {1{`RANDOM}};
  T_38110_6_ctrl_imm_sel = _RAND_2744[2:0];
  _RAND_2745 = {1{`RANDOM}};
  T_38110_6_ctrl_op_fcn = _RAND_2745[3:0];
  _RAND_2746 = {1{`RANDOM}};
  T_38110_6_ctrl_fcn_dw = _RAND_2746[0:0];
  _RAND_2747 = {1{`RANDOM}};
  T_38110_6_ctrl_rf_wen = _RAND_2747[0:0];
  _RAND_2748 = {1{`RANDOM}};
  T_38110_6_ctrl_csr_cmd = _RAND_2748[2:0];
  _RAND_2749 = {1{`RANDOM}};
  T_38110_6_ctrl_is_load = _RAND_2749[0:0];
  _RAND_2750 = {1{`RANDOM}};
  T_38110_6_ctrl_is_sta = _RAND_2750[0:0];
  _RAND_2751 = {1{`RANDOM}};
  T_38110_6_ctrl_is_std = _RAND_2751[0:0];
  _RAND_2752 = {1{`RANDOM}};
  T_38110_6_wakeup_delay = _RAND_2752[1:0];
  _RAND_2753 = {1{`RANDOM}};
  T_38110_6_allocate_brtag = _RAND_2753[0:0];
  _RAND_2754 = {1{`RANDOM}};
  T_38110_6_is_br_or_jmp = _RAND_2754[0:0];
  _RAND_2755 = {1{`RANDOM}};
  T_38110_6_is_jump = _RAND_2755[0:0];
  _RAND_2756 = {1{`RANDOM}};
  T_38110_6_is_jal = _RAND_2756[0:0];
  _RAND_2757 = {1{`RANDOM}};
  T_38110_6_is_ret = _RAND_2757[0:0];
  _RAND_2758 = {1{`RANDOM}};
  T_38110_6_is_call = _RAND_2758[0:0];
  _RAND_2759 = {1{`RANDOM}};
  T_38110_6_br_mask = _RAND_2759[7:0];
  _RAND_2760 = {1{`RANDOM}};
  T_38110_6_br_tag = _RAND_2760[2:0];
  _RAND_2761 = {1{`RANDOM}};
  T_38110_6_br_prediction_bpd_predict_val = _RAND_2761[0:0];
  _RAND_2762 = {1{`RANDOM}};
  T_38110_6_br_prediction_bpd_predict_taken = _RAND_2762[0:0];
  _RAND_2763 = {1{`RANDOM}};
  T_38110_6_br_prediction_btb_hit = _RAND_2763[0:0];
  _RAND_2764 = {1{`RANDOM}};
  T_38110_6_br_prediction_btb_predicted = _RAND_2764[0:0];
  _RAND_2765 = {1{`RANDOM}};
  T_38110_6_br_prediction_is_br_or_jalr = _RAND_2765[0:0];
  _RAND_2766 = {1{`RANDOM}};
  T_38110_6_stat_brjmp_mispredicted = _RAND_2766[0:0];
  _RAND_2767 = {1{`RANDOM}};
  T_38110_6_stat_btb_made_pred = _RAND_2767[0:0];
  _RAND_2768 = {1{`RANDOM}};
  T_38110_6_stat_btb_mispredicted = _RAND_2768[0:0];
  _RAND_2769 = {1{`RANDOM}};
  T_38110_6_stat_bpd_made_pred = _RAND_2769[0:0];
  _RAND_2770 = {1{`RANDOM}};
  T_38110_6_stat_bpd_mispredicted = _RAND_2770[0:0];
  _RAND_2771 = {1{`RANDOM}};
  T_38110_6_fetch_pc_lob = _RAND_2771[2:0];
  _RAND_2772 = {1{`RANDOM}};
  T_38110_6_imm_packed = _RAND_2772[19:0];
  _RAND_2773 = {1{`RANDOM}};
  T_38110_6_csr_addr = _RAND_2773[11:0];
  _RAND_2774 = {1{`RANDOM}};
  T_38110_6_rob_idx = _RAND_2774[5:0];
  _RAND_2775 = {1{`RANDOM}};
  T_38110_6_ldq_idx = _RAND_2775[3:0];
  _RAND_2776 = {1{`RANDOM}};
  T_38110_6_stq_idx = _RAND_2776[3:0];
  _RAND_2777 = {1{`RANDOM}};
  T_38110_6_brob_idx = _RAND_2777[4:0];
  _RAND_2778 = {1{`RANDOM}};
  T_38110_6_pdst = _RAND_2778[6:0];
  _RAND_2779 = {1{`RANDOM}};
  T_38110_6_pop1 = _RAND_2779[6:0];
  _RAND_2780 = {1{`RANDOM}};
  T_38110_6_pop2 = _RAND_2780[6:0];
  _RAND_2781 = {1{`RANDOM}};
  T_38110_6_pop3 = _RAND_2781[6:0];
  _RAND_2782 = {1{`RANDOM}};
  T_38110_6_prs1_busy = _RAND_2782[0:0];
  _RAND_2783 = {1{`RANDOM}};
  T_38110_6_prs2_busy = _RAND_2783[0:0];
  _RAND_2784 = {1{`RANDOM}};
  T_38110_6_prs3_busy = _RAND_2784[0:0];
  _RAND_2785 = {1{`RANDOM}};
  T_38110_6_stale_pdst = _RAND_2785[6:0];
  _RAND_2786 = {1{`RANDOM}};
  T_38110_6_exception = _RAND_2786[0:0];
  _RAND_2787 = {2{`RANDOM}};
  T_38110_6_exc_cause = _RAND_2787[63:0];
  _RAND_2788 = {1{`RANDOM}};
  T_38110_6_bypassable = _RAND_2788[0:0];
  _RAND_2789 = {1{`RANDOM}};
  T_38110_6_mem_cmd = _RAND_2789[3:0];
  _RAND_2790 = {1{`RANDOM}};
  T_38110_6_mem_typ = _RAND_2790[2:0];
  _RAND_2791 = {1{`RANDOM}};
  T_38110_6_is_fence = _RAND_2791[0:0];
  _RAND_2792 = {1{`RANDOM}};
  T_38110_6_is_fencei = _RAND_2792[0:0];
  _RAND_2793 = {1{`RANDOM}};
  T_38110_6_is_store = _RAND_2793[0:0];
  _RAND_2794 = {1{`RANDOM}};
  T_38110_6_is_amo = _RAND_2794[0:0];
  _RAND_2795 = {1{`RANDOM}};
  T_38110_6_is_load = _RAND_2795[0:0];
  _RAND_2796 = {1{`RANDOM}};
  T_38110_6_is_unique = _RAND_2796[0:0];
  _RAND_2797 = {1{`RANDOM}};
  T_38110_6_flush_on_commit = _RAND_2797[0:0];
  _RAND_2798 = {1{`RANDOM}};
  T_38110_6_ldst = _RAND_2798[5:0];
  _RAND_2799 = {1{`RANDOM}};
  T_38110_6_lrs1 = _RAND_2799[5:0];
  _RAND_2800 = {1{`RANDOM}};
  T_38110_6_lrs2 = _RAND_2800[5:0];
  _RAND_2801 = {1{`RANDOM}};
  T_38110_6_lrs3 = _RAND_2801[5:0];
  _RAND_2802 = {1{`RANDOM}};
  T_38110_6_ldst_val = _RAND_2802[0:0];
  _RAND_2803 = {1{`RANDOM}};
  T_38110_6_dst_rtype = _RAND_2803[1:0];
  _RAND_2804 = {1{`RANDOM}};
  T_38110_6_lrs1_rtype = _RAND_2804[1:0];
  _RAND_2805 = {1{`RANDOM}};
  T_38110_6_lrs2_rtype = _RAND_2805[1:0];
  _RAND_2806 = {1{`RANDOM}};
  T_38110_6_frs3_en = _RAND_2806[0:0];
  _RAND_2807 = {1{`RANDOM}};
  T_38110_6_fp_val = _RAND_2807[0:0];
  _RAND_2808 = {1{`RANDOM}};
  T_38110_6_fp_single = _RAND_2808[0:0];
  _RAND_2809 = {1{`RANDOM}};
  T_38110_6_xcpt_if = _RAND_2809[0:0];
  _RAND_2810 = {1{`RANDOM}};
  T_38110_6_replay_if = _RAND_2810[0:0];
  _RAND_2811 = {2{`RANDOM}};
  T_38110_6_debug_wdata = _RAND_2811[63:0];
  _RAND_2812 = {1{`RANDOM}};
  T_38110_6_debug_events_fetch_seq = _RAND_2812[31:0];
  _RAND_2813 = {1{`RANDOM}};
  T_38110_7_valid = _RAND_2813[0:0];
  _RAND_2814 = {1{`RANDOM}};
  T_38110_7_iw_state = _RAND_2814[1:0];
  _RAND_2815 = {1{`RANDOM}};
  T_38110_7_uopc = _RAND_2815[8:0];
  _RAND_2816 = {1{`RANDOM}};
  T_38110_7_inst = _RAND_2816[31:0];
  _RAND_2817 = {2{`RANDOM}};
  T_38110_7_pc = _RAND_2817[39:0];
  _RAND_2818 = {1{`RANDOM}};
  T_38110_7_fu_code = _RAND_2818[7:0];
  _RAND_2819 = {1{`RANDOM}};
  T_38110_7_ctrl_br_type = _RAND_2819[3:0];
  _RAND_2820 = {1{`RANDOM}};
  T_38110_7_ctrl_op1_sel = _RAND_2820[1:0];
  _RAND_2821 = {1{`RANDOM}};
  T_38110_7_ctrl_op2_sel = _RAND_2821[2:0];
  _RAND_2822 = {1{`RANDOM}};
  T_38110_7_ctrl_imm_sel = _RAND_2822[2:0];
  _RAND_2823 = {1{`RANDOM}};
  T_38110_7_ctrl_op_fcn = _RAND_2823[3:0];
  _RAND_2824 = {1{`RANDOM}};
  T_38110_7_ctrl_fcn_dw = _RAND_2824[0:0];
  _RAND_2825 = {1{`RANDOM}};
  T_38110_7_ctrl_rf_wen = _RAND_2825[0:0];
  _RAND_2826 = {1{`RANDOM}};
  T_38110_7_ctrl_csr_cmd = _RAND_2826[2:0];
  _RAND_2827 = {1{`RANDOM}};
  T_38110_7_ctrl_is_load = _RAND_2827[0:0];
  _RAND_2828 = {1{`RANDOM}};
  T_38110_7_ctrl_is_sta = _RAND_2828[0:0];
  _RAND_2829 = {1{`RANDOM}};
  T_38110_7_ctrl_is_std = _RAND_2829[0:0];
  _RAND_2830 = {1{`RANDOM}};
  T_38110_7_wakeup_delay = _RAND_2830[1:0];
  _RAND_2831 = {1{`RANDOM}};
  T_38110_7_allocate_brtag = _RAND_2831[0:0];
  _RAND_2832 = {1{`RANDOM}};
  T_38110_7_is_br_or_jmp = _RAND_2832[0:0];
  _RAND_2833 = {1{`RANDOM}};
  T_38110_7_is_jump = _RAND_2833[0:0];
  _RAND_2834 = {1{`RANDOM}};
  T_38110_7_is_jal = _RAND_2834[0:0];
  _RAND_2835 = {1{`RANDOM}};
  T_38110_7_is_ret = _RAND_2835[0:0];
  _RAND_2836 = {1{`RANDOM}};
  T_38110_7_is_call = _RAND_2836[0:0];
  _RAND_2837 = {1{`RANDOM}};
  T_38110_7_br_mask = _RAND_2837[7:0];
  _RAND_2838 = {1{`RANDOM}};
  T_38110_7_br_tag = _RAND_2838[2:0];
  _RAND_2839 = {1{`RANDOM}};
  T_38110_7_br_prediction_bpd_predict_val = _RAND_2839[0:0];
  _RAND_2840 = {1{`RANDOM}};
  T_38110_7_br_prediction_bpd_predict_taken = _RAND_2840[0:0];
  _RAND_2841 = {1{`RANDOM}};
  T_38110_7_br_prediction_btb_hit = _RAND_2841[0:0];
  _RAND_2842 = {1{`RANDOM}};
  T_38110_7_br_prediction_btb_predicted = _RAND_2842[0:0];
  _RAND_2843 = {1{`RANDOM}};
  T_38110_7_br_prediction_is_br_or_jalr = _RAND_2843[0:0];
  _RAND_2844 = {1{`RANDOM}};
  T_38110_7_stat_brjmp_mispredicted = _RAND_2844[0:0];
  _RAND_2845 = {1{`RANDOM}};
  T_38110_7_stat_btb_made_pred = _RAND_2845[0:0];
  _RAND_2846 = {1{`RANDOM}};
  T_38110_7_stat_btb_mispredicted = _RAND_2846[0:0];
  _RAND_2847 = {1{`RANDOM}};
  T_38110_7_stat_bpd_made_pred = _RAND_2847[0:0];
  _RAND_2848 = {1{`RANDOM}};
  T_38110_7_stat_bpd_mispredicted = _RAND_2848[0:0];
  _RAND_2849 = {1{`RANDOM}};
  T_38110_7_fetch_pc_lob = _RAND_2849[2:0];
  _RAND_2850 = {1{`RANDOM}};
  T_38110_7_imm_packed = _RAND_2850[19:0];
  _RAND_2851 = {1{`RANDOM}};
  T_38110_7_csr_addr = _RAND_2851[11:0];
  _RAND_2852 = {1{`RANDOM}};
  T_38110_7_rob_idx = _RAND_2852[5:0];
  _RAND_2853 = {1{`RANDOM}};
  T_38110_7_ldq_idx = _RAND_2853[3:0];
  _RAND_2854 = {1{`RANDOM}};
  T_38110_7_stq_idx = _RAND_2854[3:0];
  _RAND_2855 = {1{`RANDOM}};
  T_38110_7_brob_idx = _RAND_2855[4:0];
  _RAND_2856 = {1{`RANDOM}};
  T_38110_7_pdst = _RAND_2856[6:0];
  _RAND_2857 = {1{`RANDOM}};
  T_38110_7_pop1 = _RAND_2857[6:0];
  _RAND_2858 = {1{`RANDOM}};
  T_38110_7_pop2 = _RAND_2858[6:0];
  _RAND_2859 = {1{`RANDOM}};
  T_38110_7_pop3 = _RAND_2859[6:0];
  _RAND_2860 = {1{`RANDOM}};
  T_38110_7_prs1_busy = _RAND_2860[0:0];
  _RAND_2861 = {1{`RANDOM}};
  T_38110_7_prs2_busy = _RAND_2861[0:0];
  _RAND_2862 = {1{`RANDOM}};
  T_38110_7_prs3_busy = _RAND_2862[0:0];
  _RAND_2863 = {1{`RANDOM}};
  T_38110_7_stale_pdst = _RAND_2863[6:0];
  _RAND_2864 = {1{`RANDOM}};
  T_38110_7_exception = _RAND_2864[0:0];
  _RAND_2865 = {2{`RANDOM}};
  T_38110_7_exc_cause = _RAND_2865[63:0];
  _RAND_2866 = {1{`RANDOM}};
  T_38110_7_bypassable = _RAND_2866[0:0];
  _RAND_2867 = {1{`RANDOM}};
  T_38110_7_mem_cmd = _RAND_2867[3:0];
  _RAND_2868 = {1{`RANDOM}};
  T_38110_7_mem_typ = _RAND_2868[2:0];
  _RAND_2869 = {1{`RANDOM}};
  T_38110_7_is_fence = _RAND_2869[0:0];
  _RAND_2870 = {1{`RANDOM}};
  T_38110_7_is_fencei = _RAND_2870[0:0];
  _RAND_2871 = {1{`RANDOM}};
  T_38110_7_is_store = _RAND_2871[0:0];
  _RAND_2872 = {1{`RANDOM}};
  T_38110_7_is_amo = _RAND_2872[0:0];
  _RAND_2873 = {1{`RANDOM}};
  T_38110_7_is_load = _RAND_2873[0:0];
  _RAND_2874 = {1{`RANDOM}};
  T_38110_7_is_unique = _RAND_2874[0:0];
  _RAND_2875 = {1{`RANDOM}};
  T_38110_7_flush_on_commit = _RAND_2875[0:0];
  _RAND_2876 = {1{`RANDOM}};
  T_38110_7_ldst = _RAND_2876[5:0];
  _RAND_2877 = {1{`RANDOM}};
  T_38110_7_lrs1 = _RAND_2877[5:0];
  _RAND_2878 = {1{`RANDOM}};
  T_38110_7_lrs2 = _RAND_2878[5:0];
  _RAND_2879 = {1{`RANDOM}};
  T_38110_7_lrs3 = _RAND_2879[5:0];
  _RAND_2880 = {1{`RANDOM}};
  T_38110_7_ldst_val = _RAND_2880[0:0];
  _RAND_2881 = {1{`RANDOM}};
  T_38110_7_dst_rtype = _RAND_2881[1:0];
  _RAND_2882 = {1{`RANDOM}};
  T_38110_7_lrs1_rtype = _RAND_2882[1:0];
  _RAND_2883 = {1{`RANDOM}};
  T_38110_7_lrs2_rtype = _RAND_2883[1:0];
  _RAND_2884 = {1{`RANDOM}};
  T_38110_7_frs3_en = _RAND_2884[0:0];
  _RAND_2885 = {1{`RANDOM}};
  T_38110_7_fp_val = _RAND_2885[0:0];
  _RAND_2886 = {1{`RANDOM}};
  T_38110_7_fp_single = _RAND_2886[0:0];
  _RAND_2887 = {1{`RANDOM}};
  T_38110_7_xcpt_if = _RAND_2887[0:0];
  _RAND_2888 = {1{`RANDOM}};
  T_38110_7_replay_if = _RAND_2888[0:0];
  _RAND_2889 = {2{`RANDOM}};
  T_38110_7_debug_wdata = _RAND_2889[63:0];
  _RAND_2890 = {1{`RANDOM}};
  T_38110_7_debug_events_fetch_seq = _RAND_2890[31:0];
  _RAND_2891 = {1{`RANDOM}};
  T_38110_8_valid = _RAND_2891[0:0];
  _RAND_2892 = {1{`RANDOM}};
  T_38110_8_iw_state = _RAND_2892[1:0];
  _RAND_2893 = {1{`RANDOM}};
  T_38110_8_uopc = _RAND_2893[8:0];
  _RAND_2894 = {1{`RANDOM}};
  T_38110_8_inst = _RAND_2894[31:0];
  _RAND_2895 = {2{`RANDOM}};
  T_38110_8_pc = _RAND_2895[39:0];
  _RAND_2896 = {1{`RANDOM}};
  T_38110_8_fu_code = _RAND_2896[7:0];
  _RAND_2897 = {1{`RANDOM}};
  T_38110_8_ctrl_br_type = _RAND_2897[3:0];
  _RAND_2898 = {1{`RANDOM}};
  T_38110_8_ctrl_op1_sel = _RAND_2898[1:0];
  _RAND_2899 = {1{`RANDOM}};
  T_38110_8_ctrl_op2_sel = _RAND_2899[2:0];
  _RAND_2900 = {1{`RANDOM}};
  T_38110_8_ctrl_imm_sel = _RAND_2900[2:0];
  _RAND_2901 = {1{`RANDOM}};
  T_38110_8_ctrl_op_fcn = _RAND_2901[3:0];
  _RAND_2902 = {1{`RANDOM}};
  T_38110_8_ctrl_fcn_dw = _RAND_2902[0:0];
  _RAND_2903 = {1{`RANDOM}};
  T_38110_8_ctrl_rf_wen = _RAND_2903[0:0];
  _RAND_2904 = {1{`RANDOM}};
  T_38110_8_ctrl_csr_cmd = _RAND_2904[2:0];
  _RAND_2905 = {1{`RANDOM}};
  T_38110_8_ctrl_is_load = _RAND_2905[0:0];
  _RAND_2906 = {1{`RANDOM}};
  T_38110_8_ctrl_is_sta = _RAND_2906[0:0];
  _RAND_2907 = {1{`RANDOM}};
  T_38110_8_ctrl_is_std = _RAND_2907[0:0];
  _RAND_2908 = {1{`RANDOM}};
  T_38110_8_wakeup_delay = _RAND_2908[1:0];
  _RAND_2909 = {1{`RANDOM}};
  T_38110_8_allocate_brtag = _RAND_2909[0:0];
  _RAND_2910 = {1{`RANDOM}};
  T_38110_8_is_br_or_jmp = _RAND_2910[0:0];
  _RAND_2911 = {1{`RANDOM}};
  T_38110_8_is_jump = _RAND_2911[0:0];
  _RAND_2912 = {1{`RANDOM}};
  T_38110_8_is_jal = _RAND_2912[0:0];
  _RAND_2913 = {1{`RANDOM}};
  T_38110_8_is_ret = _RAND_2913[0:0];
  _RAND_2914 = {1{`RANDOM}};
  T_38110_8_is_call = _RAND_2914[0:0];
  _RAND_2915 = {1{`RANDOM}};
  T_38110_8_br_mask = _RAND_2915[7:0];
  _RAND_2916 = {1{`RANDOM}};
  T_38110_8_br_tag = _RAND_2916[2:0];
  _RAND_2917 = {1{`RANDOM}};
  T_38110_8_br_prediction_bpd_predict_val = _RAND_2917[0:0];
  _RAND_2918 = {1{`RANDOM}};
  T_38110_8_br_prediction_bpd_predict_taken = _RAND_2918[0:0];
  _RAND_2919 = {1{`RANDOM}};
  T_38110_8_br_prediction_btb_hit = _RAND_2919[0:0];
  _RAND_2920 = {1{`RANDOM}};
  T_38110_8_br_prediction_btb_predicted = _RAND_2920[0:0];
  _RAND_2921 = {1{`RANDOM}};
  T_38110_8_br_prediction_is_br_or_jalr = _RAND_2921[0:0];
  _RAND_2922 = {1{`RANDOM}};
  T_38110_8_stat_brjmp_mispredicted = _RAND_2922[0:0];
  _RAND_2923 = {1{`RANDOM}};
  T_38110_8_stat_btb_made_pred = _RAND_2923[0:0];
  _RAND_2924 = {1{`RANDOM}};
  T_38110_8_stat_btb_mispredicted = _RAND_2924[0:0];
  _RAND_2925 = {1{`RANDOM}};
  T_38110_8_stat_bpd_made_pred = _RAND_2925[0:0];
  _RAND_2926 = {1{`RANDOM}};
  T_38110_8_stat_bpd_mispredicted = _RAND_2926[0:0];
  _RAND_2927 = {1{`RANDOM}};
  T_38110_8_fetch_pc_lob = _RAND_2927[2:0];
  _RAND_2928 = {1{`RANDOM}};
  T_38110_8_imm_packed = _RAND_2928[19:0];
  _RAND_2929 = {1{`RANDOM}};
  T_38110_8_csr_addr = _RAND_2929[11:0];
  _RAND_2930 = {1{`RANDOM}};
  T_38110_8_rob_idx = _RAND_2930[5:0];
  _RAND_2931 = {1{`RANDOM}};
  T_38110_8_ldq_idx = _RAND_2931[3:0];
  _RAND_2932 = {1{`RANDOM}};
  T_38110_8_stq_idx = _RAND_2932[3:0];
  _RAND_2933 = {1{`RANDOM}};
  T_38110_8_brob_idx = _RAND_2933[4:0];
  _RAND_2934 = {1{`RANDOM}};
  T_38110_8_pdst = _RAND_2934[6:0];
  _RAND_2935 = {1{`RANDOM}};
  T_38110_8_pop1 = _RAND_2935[6:0];
  _RAND_2936 = {1{`RANDOM}};
  T_38110_8_pop2 = _RAND_2936[6:0];
  _RAND_2937 = {1{`RANDOM}};
  T_38110_8_pop3 = _RAND_2937[6:0];
  _RAND_2938 = {1{`RANDOM}};
  T_38110_8_prs1_busy = _RAND_2938[0:0];
  _RAND_2939 = {1{`RANDOM}};
  T_38110_8_prs2_busy = _RAND_2939[0:0];
  _RAND_2940 = {1{`RANDOM}};
  T_38110_8_prs3_busy = _RAND_2940[0:0];
  _RAND_2941 = {1{`RANDOM}};
  T_38110_8_stale_pdst = _RAND_2941[6:0];
  _RAND_2942 = {1{`RANDOM}};
  T_38110_8_exception = _RAND_2942[0:0];
  _RAND_2943 = {2{`RANDOM}};
  T_38110_8_exc_cause = _RAND_2943[63:0];
  _RAND_2944 = {1{`RANDOM}};
  T_38110_8_bypassable = _RAND_2944[0:0];
  _RAND_2945 = {1{`RANDOM}};
  T_38110_8_mem_cmd = _RAND_2945[3:0];
  _RAND_2946 = {1{`RANDOM}};
  T_38110_8_mem_typ = _RAND_2946[2:0];
  _RAND_2947 = {1{`RANDOM}};
  T_38110_8_is_fence = _RAND_2947[0:0];
  _RAND_2948 = {1{`RANDOM}};
  T_38110_8_is_fencei = _RAND_2948[0:0];
  _RAND_2949 = {1{`RANDOM}};
  T_38110_8_is_store = _RAND_2949[0:0];
  _RAND_2950 = {1{`RANDOM}};
  T_38110_8_is_amo = _RAND_2950[0:0];
  _RAND_2951 = {1{`RANDOM}};
  T_38110_8_is_load = _RAND_2951[0:0];
  _RAND_2952 = {1{`RANDOM}};
  T_38110_8_is_unique = _RAND_2952[0:0];
  _RAND_2953 = {1{`RANDOM}};
  T_38110_8_flush_on_commit = _RAND_2953[0:0];
  _RAND_2954 = {1{`RANDOM}};
  T_38110_8_ldst = _RAND_2954[5:0];
  _RAND_2955 = {1{`RANDOM}};
  T_38110_8_lrs1 = _RAND_2955[5:0];
  _RAND_2956 = {1{`RANDOM}};
  T_38110_8_lrs2 = _RAND_2956[5:0];
  _RAND_2957 = {1{`RANDOM}};
  T_38110_8_lrs3 = _RAND_2957[5:0];
  _RAND_2958 = {1{`RANDOM}};
  T_38110_8_ldst_val = _RAND_2958[0:0];
  _RAND_2959 = {1{`RANDOM}};
  T_38110_8_dst_rtype = _RAND_2959[1:0];
  _RAND_2960 = {1{`RANDOM}};
  T_38110_8_lrs1_rtype = _RAND_2960[1:0];
  _RAND_2961 = {1{`RANDOM}};
  T_38110_8_lrs2_rtype = _RAND_2961[1:0];
  _RAND_2962 = {1{`RANDOM}};
  T_38110_8_frs3_en = _RAND_2962[0:0];
  _RAND_2963 = {1{`RANDOM}};
  T_38110_8_fp_val = _RAND_2963[0:0];
  _RAND_2964 = {1{`RANDOM}};
  T_38110_8_fp_single = _RAND_2964[0:0];
  _RAND_2965 = {1{`RANDOM}};
  T_38110_8_xcpt_if = _RAND_2965[0:0];
  _RAND_2966 = {1{`RANDOM}};
  T_38110_8_replay_if = _RAND_2966[0:0];
  _RAND_2967 = {2{`RANDOM}};
  T_38110_8_debug_wdata = _RAND_2967[63:0];
  _RAND_2968 = {1{`RANDOM}};
  T_38110_8_debug_events_fetch_seq = _RAND_2968[31:0];
  _RAND_2969 = {1{`RANDOM}};
  T_38110_9_valid = _RAND_2969[0:0];
  _RAND_2970 = {1{`RANDOM}};
  T_38110_9_iw_state = _RAND_2970[1:0];
  _RAND_2971 = {1{`RANDOM}};
  T_38110_9_uopc = _RAND_2971[8:0];
  _RAND_2972 = {1{`RANDOM}};
  T_38110_9_inst = _RAND_2972[31:0];
  _RAND_2973 = {2{`RANDOM}};
  T_38110_9_pc = _RAND_2973[39:0];
  _RAND_2974 = {1{`RANDOM}};
  T_38110_9_fu_code = _RAND_2974[7:0];
  _RAND_2975 = {1{`RANDOM}};
  T_38110_9_ctrl_br_type = _RAND_2975[3:0];
  _RAND_2976 = {1{`RANDOM}};
  T_38110_9_ctrl_op1_sel = _RAND_2976[1:0];
  _RAND_2977 = {1{`RANDOM}};
  T_38110_9_ctrl_op2_sel = _RAND_2977[2:0];
  _RAND_2978 = {1{`RANDOM}};
  T_38110_9_ctrl_imm_sel = _RAND_2978[2:0];
  _RAND_2979 = {1{`RANDOM}};
  T_38110_9_ctrl_op_fcn = _RAND_2979[3:0];
  _RAND_2980 = {1{`RANDOM}};
  T_38110_9_ctrl_fcn_dw = _RAND_2980[0:0];
  _RAND_2981 = {1{`RANDOM}};
  T_38110_9_ctrl_rf_wen = _RAND_2981[0:0];
  _RAND_2982 = {1{`RANDOM}};
  T_38110_9_ctrl_csr_cmd = _RAND_2982[2:0];
  _RAND_2983 = {1{`RANDOM}};
  T_38110_9_ctrl_is_load = _RAND_2983[0:0];
  _RAND_2984 = {1{`RANDOM}};
  T_38110_9_ctrl_is_sta = _RAND_2984[0:0];
  _RAND_2985 = {1{`RANDOM}};
  T_38110_9_ctrl_is_std = _RAND_2985[0:0];
  _RAND_2986 = {1{`RANDOM}};
  T_38110_9_wakeup_delay = _RAND_2986[1:0];
  _RAND_2987 = {1{`RANDOM}};
  T_38110_9_allocate_brtag = _RAND_2987[0:0];
  _RAND_2988 = {1{`RANDOM}};
  T_38110_9_is_br_or_jmp = _RAND_2988[0:0];
  _RAND_2989 = {1{`RANDOM}};
  T_38110_9_is_jump = _RAND_2989[0:0];
  _RAND_2990 = {1{`RANDOM}};
  T_38110_9_is_jal = _RAND_2990[0:0];
  _RAND_2991 = {1{`RANDOM}};
  T_38110_9_is_ret = _RAND_2991[0:0];
  _RAND_2992 = {1{`RANDOM}};
  T_38110_9_is_call = _RAND_2992[0:0];
  _RAND_2993 = {1{`RANDOM}};
  T_38110_9_br_mask = _RAND_2993[7:0];
  _RAND_2994 = {1{`RANDOM}};
  T_38110_9_br_tag = _RAND_2994[2:0];
  _RAND_2995 = {1{`RANDOM}};
  T_38110_9_br_prediction_bpd_predict_val = _RAND_2995[0:0];
  _RAND_2996 = {1{`RANDOM}};
  T_38110_9_br_prediction_bpd_predict_taken = _RAND_2996[0:0];
  _RAND_2997 = {1{`RANDOM}};
  T_38110_9_br_prediction_btb_hit = _RAND_2997[0:0];
  _RAND_2998 = {1{`RANDOM}};
  T_38110_9_br_prediction_btb_predicted = _RAND_2998[0:0];
  _RAND_2999 = {1{`RANDOM}};
  T_38110_9_br_prediction_is_br_or_jalr = _RAND_2999[0:0];
  _RAND_3000 = {1{`RANDOM}};
  T_38110_9_stat_brjmp_mispredicted = _RAND_3000[0:0];
  _RAND_3001 = {1{`RANDOM}};
  T_38110_9_stat_btb_made_pred = _RAND_3001[0:0];
  _RAND_3002 = {1{`RANDOM}};
  T_38110_9_stat_btb_mispredicted = _RAND_3002[0:0];
  _RAND_3003 = {1{`RANDOM}};
  T_38110_9_stat_bpd_made_pred = _RAND_3003[0:0];
  _RAND_3004 = {1{`RANDOM}};
  T_38110_9_stat_bpd_mispredicted = _RAND_3004[0:0];
  _RAND_3005 = {1{`RANDOM}};
  T_38110_9_fetch_pc_lob = _RAND_3005[2:0];
  _RAND_3006 = {1{`RANDOM}};
  T_38110_9_imm_packed = _RAND_3006[19:0];
  _RAND_3007 = {1{`RANDOM}};
  T_38110_9_csr_addr = _RAND_3007[11:0];
  _RAND_3008 = {1{`RANDOM}};
  T_38110_9_rob_idx = _RAND_3008[5:0];
  _RAND_3009 = {1{`RANDOM}};
  T_38110_9_ldq_idx = _RAND_3009[3:0];
  _RAND_3010 = {1{`RANDOM}};
  T_38110_9_stq_idx = _RAND_3010[3:0];
  _RAND_3011 = {1{`RANDOM}};
  T_38110_9_brob_idx = _RAND_3011[4:0];
  _RAND_3012 = {1{`RANDOM}};
  T_38110_9_pdst = _RAND_3012[6:0];
  _RAND_3013 = {1{`RANDOM}};
  T_38110_9_pop1 = _RAND_3013[6:0];
  _RAND_3014 = {1{`RANDOM}};
  T_38110_9_pop2 = _RAND_3014[6:0];
  _RAND_3015 = {1{`RANDOM}};
  T_38110_9_pop3 = _RAND_3015[6:0];
  _RAND_3016 = {1{`RANDOM}};
  T_38110_9_prs1_busy = _RAND_3016[0:0];
  _RAND_3017 = {1{`RANDOM}};
  T_38110_9_prs2_busy = _RAND_3017[0:0];
  _RAND_3018 = {1{`RANDOM}};
  T_38110_9_prs3_busy = _RAND_3018[0:0];
  _RAND_3019 = {1{`RANDOM}};
  T_38110_9_stale_pdst = _RAND_3019[6:0];
  _RAND_3020 = {1{`RANDOM}};
  T_38110_9_exception = _RAND_3020[0:0];
  _RAND_3021 = {2{`RANDOM}};
  T_38110_9_exc_cause = _RAND_3021[63:0];
  _RAND_3022 = {1{`RANDOM}};
  T_38110_9_bypassable = _RAND_3022[0:0];
  _RAND_3023 = {1{`RANDOM}};
  T_38110_9_mem_cmd = _RAND_3023[3:0];
  _RAND_3024 = {1{`RANDOM}};
  T_38110_9_mem_typ = _RAND_3024[2:0];
  _RAND_3025 = {1{`RANDOM}};
  T_38110_9_is_fence = _RAND_3025[0:0];
  _RAND_3026 = {1{`RANDOM}};
  T_38110_9_is_fencei = _RAND_3026[0:0];
  _RAND_3027 = {1{`RANDOM}};
  T_38110_9_is_store = _RAND_3027[0:0];
  _RAND_3028 = {1{`RANDOM}};
  T_38110_9_is_amo = _RAND_3028[0:0];
  _RAND_3029 = {1{`RANDOM}};
  T_38110_9_is_load = _RAND_3029[0:0];
  _RAND_3030 = {1{`RANDOM}};
  T_38110_9_is_unique = _RAND_3030[0:0];
  _RAND_3031 = {1{`RANDOM}};
  T_38110_9_flush_on_commit = _RAND_3031[0:0];
  _RAND_3032 = {1{`RANDOM}};
  T_38110_9_ldst = _RAND_3032[5:0];
  _RAND_3033 = {1{`RANDOM}};
  T_38110_9_lrs1 = _RAND_3033[5:0];
  _RAND_3034 = {1{`RANDOM}};
  T_38110_9_lrs2 = _RAND_3034[5:0];
  _RAND_3035 = {1{`RANDOM}};
  T_38110_9_lrs3 = _RAND_3035[5:0];
  _RAND_3036 = {1{`RANDOM}};
  T_38110_9_ldst_val = _RAND_3036[0:0];
  _RAND_3037 = {1{`RANDOM}};
  T_38110_9_dst_rtype = _RAND_3037[1:0];
  _RAND_3038 = {1{`RANDOM}};
  T_38110_9_lrs1_rtype = _RAND_3038[1:0];
  _RAND_3039 = {1{`RANDOM}};
  T_38110_9_lrs2_rtype = _RAND_3039[1:0];
  _RAND_3040 = {1{`RANDOM}};
  T_38110_9_frs3_en = _RAND_3040[0:0];
  _RAND_3041 = {1{`RANDOM}};
  T_38110_9_fp_val = _RAND_3041[0:0];
  _RAND_3042 = {1{`RANDOM}};
  T_38110_9_fp_single = _RAND_3042[0:0];
  _RAND_3043 = {1{`RANDOM}};
  T_38110_9_xcpt_if = _RAND_3043[0:0];
  _RAND_3044 = {1{`RANDOM}};
  T_38110_9_replay_if = _RAND_3044[0:0];
  _RAND_3045 = {2{`RANDOM}};
  T_38110_9_debug_wdata = _RAND_3045[63:0];
  _RAND_3046 = {1{`RANDOM}};
  T_38110_9_debug_events_fetch_seq = _RAND_3046[31:0];
  _RAND_3047 = {1{`RANDOM}};
  T_38110_10_valid = _RAND_3047[0:0];
  _RAND_3048 = {1{`RANDOM}};
  T_38110_10_iw_state = _RAND_3048[1:0];
  _RAND_3049 = {1{`RANDOM}};
  T_38110_10_uopc = _RAND_3049[8:0];
  _RAND_3050 = {1{`RANDOM}};
  T_38110_10_inst = _RAND_3050[31:0];
  _RAND_3051 = {2{`RANDOM}};
  T_38110_10_pc = _RAND_3051[39:0];
  _RAND_3052 = {1{`RANDOM}};
  T_38110_10_fu_code = _RAND_3052[7:0];
  _RAND_3053 = {1{`RANDOM}};
  T_38110_10_ctrl_br_type = _RAND_3053[3:0];
  _RAND_3054 = {1{`RANDOM}};
  T_38110_10_ctrl_op1_sel = _RAND_3054[1:0];
  _RAND_3055 = {1{`RANDOM}};
  T_38110_10_ctrl_op2_sel = _RAND_3055[2:0];
  _RAND_3056 = {1{`RANDOM}};
  T_38110_10_ctrl_imm_sel = _RAND_3056[2:0];
  _RAND_3057 = {1{`RANDOM}};
  T_38110_10_ctrl_op_fcn = _RAND_3057[3:0];
  _RAND_3058 = {1{`RANDOM}};
  T_38110_10_ctrl_fcn_dw = _RAND_3058[0:0];
  _RAND_3059 = {1{`RANDOM}};
  T_38110_10_ctrl_rf_wen = _RAND_3059[0:0];
  _RAND_3060 = {1{`RANDOM}};
  T_38110_10_ctrl_csr_cmd = _RAND_3060[2:0];
  _RAND_3061 = {1{`RANDOM}};
  T_38110_10_ctrl_is_load = _RAND_3061[0:0];
  _RAND_3062 = {1{`RANDOM}};
  T_38110_10_ctrl_is_sta = _RAND_3062[0:0];
  _RAND_3063 = {1{`RANDOM}};
  T_38110_10_ctrl_is_std = _RAND_3063[0:0];
  _RAND_3064 = {1{`RANDOM}};
  T_38110_10_wakeup_delay = _RAND_3064[1:0];
  _RAND_3065 = {1{`RANDOM}};
  T_38110_10_allocate_brtag = _RAND_3065[0:0];
  _RAND_3066 = {1{`RANDOM}};
  T_38110_10_is_br_or_jmp = _RAND_3066[0:0];
  _RAND_3067 = {1{`RANDOM}};
  T_38110_10_is_jump = _RAND_3067[0:0];
  _RAND_3068 = {1{`RANDOM}};
  T_38110_10_is_jal = _RAND_3068[0:0];
  _RAND_3069 = {1{`RANDOM}};
  T_38110_10_is_ret = _RAND_3069[0:0];
  _RAND_3070 = {1{`RANDOM}};
  T_38110_10_is_call = _RAND_3070[0:0];
  _RAND_3071 = {1{`RANDOM}};
  T_38110_10_br_mask = _RAND_3071[7:0];
  _RAND_3072 = {1{`RANDOM}};
  T_38110_10_br_tag = _RAND_3072[2:0];
  _RAND_3073 = {1{`RANDOM}};
  T_38110_10_br_prediction_bpd_predict_val = _RAND_3073[0:0];
  _RAND_3074 = {1{`RANDOM}};
  T_38110_10_br_prediction_bpd_predict_taken = _RAND_3074[0:0];
  _RAND_3075 = {1{`RANDOM}};
  T_38110_10_br_prediction_btb_hit = _RAND_3075[0:0];
  _RAND_3076 = {1{`RANDOM}};
  T_38110_10_br_prediction_btb_predicted = _RAND_3076[0:0];
  _RAND_3077 = {1{`RANDOM}};
  T_38110_10_br_prediction_is_br_or_jalr = _RAND_3077[0:0];
  _RAND_3078 = {1{`RANDOM}};
  T_38110_10_stat_brjmp_mispredicted = _RAND_3078[0:0];
  _RAND_3079 = {1{`RANDOM}};
  T_38110_10_stat_btb_made_pred = _RAND_3079[0:0];
  _RAND_3080 = {1{`RANDOM}};
  T_38110_10_stat_btb_mispredicted = _RAND_3080[0:0];
  _RAND_3081 = {1{`RANDOM}};
  T_38110_10_stat_bpd_made_pred = _RAND_3081[0:0];
  _RAND_3082 = {1{`RANDOM}};
  T_38110_10_stat_bpd_mispredicted = _RAND_3082[0:0];
  _RAND_3083 = {1{`RANDOM}};
  T_38110_10_fetch_pc_lob = _RAND_3083[2:0];
  _RAND_3084 = {1{`RANDOM}};
  T_38110_10_imm_packed = _RAND_3084[19:0];
  _RAND_3085 = {1{`RANDOM}};
  T_38110_10_csr_addr = _RAND_3085[11:0];
  _RAND_3086 = {1{`RANDOM}};
  T_38110_10_rob_idx = _RAND_3086[5:0];
  _RAND_3087 = {1{`RANDOM}};
  T_38110_10_ldq_idx = _RAND_3087[3:0];
  _RAND_3088 = {1{`RANDOM}};
  T_38110_10_stq_idx = _RAND_3088[3:0];
  _RAND_3089 = {1{`RANDOM}};
  T_38110_10_brob_idx = _RAND_3089[4:0];
  _RAND_3090 = {1{`RANDOM}};
  T_38110_10_pdst = _RAND_3090[6:0];
  _RAND_3091 = {1{`RANDOM}};
  T_38110_10_pop1 = _RAND_3091[6:0];
  _RAND_3092 = {1{`RANDOM}};
  T_38110_10_pop2 = _RAND_3092[6:0];
  _RAND_3093 = {1{`RANDOM}};
  T_38110_10_pop3 = _RAND_3093[6:0];
  _RAND_3094 = {1{`RANDOM}};
  T_38110_10_prs1_busy = _RAND_3094[0:0];
  _RAND_3095 = {1{`RANDOM}};
  T_38110_10_prs2_busy = _RAND_3095[0:0];
  _RAND_3096 = {1{`RANDOM}};
  T_38110_10_prs3_busy = _RAND_3096[0:0];
  _RAND_3097 = {1{`RANDOM}};
  T_38110_10_stale_pdst = _RAND_3097[6:0];
  _RAND_3098 = {1{`RANDOM}};
  T_38110_10_exception = _RAND_3098[0:0];
  _RAND_3099 = {2{`RANDOM}};
  T_38110_10_exc_cause = _RAND_3099[63:0];
  _RAND_3100 = {1{`RANDOM}};
  T_38110_10_bypassable = _RAND_3100[0:0];
  _RAND_3101 = {1{`RANDOM}};
  T_38110_10_mem_cmd = _RAND_3101[3:0];
  _RAND_3102 = {1{`RANDOM}};
  T_38110_10_mem_typ = _RAND_3102[2:0];
  _RAND_3103 = {1{`RANDOM}};
  T_38110_10_is_fence = _RAND_3103[0:0];
  _RAND_3104 = {1{`RANDOM}};
  T_38110_10_is_fencei = _RAND_3104[0:0];
  _RAND_3105 = {1{`RANDOM}};
  T_38110_10_is_store = _RAND_3105[0:0];
  _RAND_3106 = {1{`RANDOM}};
  T_38110_10_is_amo = _RAND_3106[0:0];
  _RAND_3107 = {1{`RANDOM}};
  T_38110_10_is_load = _RAND_3107[0:0];
  _RAND_3108 = {1{`RANDOM}};
  T_38110_10_is_unique = _RAND_3108[0:0];
  _RAND_3109 = {1{`RANDOM}};
  T_38110_10_flush_on_commit = _RAND_3109[0:0];
  _RAND_3110 = {1{`RANDOM}};
  T_38110_10_ldst = _RAND_3110[5:0];
  _RAND_3111 = {1{`RANDOM}};
  T_38110_10_lrs1 = _RAND_3111[5:0];
  _RAND_3112 = {1{`RANDOM}};
  T_38110_10_lrs2 = _RAND_3112[5:0];
  _RAND_3113 = {1{`RANDOM}};
  T_38110_10_lrs3 = _RAND_3113[5:0];
  _RAND_3114 = {1{`RANDOM}};
  T_38110_10_ldst_val = _RAND_3114[0:0];
  _RAND_3115 = {1{`RANDOM}};
  T_38110_10_dst_rtype = _RAND_3115[1:0];
  _RAND_3116 = {1{`RANDOM}};
  T_38110_10_lrs1_rtype = _RAND_3116[1:0];
  _RAND_3117 = {1{`RANDOM}};
  T_38110_10_lrs2_rtype = _RAND_3117[1:0];
  _RAND_3118 = {1{`RANDOM}};
  T_38110_10_frs3_en = _RAND_3118[0:0];
  _RAND_3119 = {1{`RANDOM}};
  T_38110_10_fp_val = _RAND_3119[0:0];
  _RAND_3120 = {1{`RANDOM}};
  T_38110_10_fp_single = _RAND_3120[0:0];
  _RAND_3121 = {1{`RANDOM}};
  T_38110_10_xcpt_if = _RAND_3121[0:0];
  _RAND_3122 = {1{`RANDOM}};
  T_38110_10_replay_if = _RAND_3122[0:0];
  _RAND_3123 = {2{`RANDOM}};
  T_38110_10_debug_wdata = _RAND_3123[63:0];
  _RAND_3124 = {1{`RANDOM}};
  T_38110_10_debug_events_fetch_seq = _RAND_3124[31:0];
  _RAND_3125 = {1{`RANDOM}};
  T_38110_11_valid = _RAND_3125[0:0];
  _RAND_3126 = {1{`RANDOM}};
  T_38110_11_iw_state = _RAND_3126[1:0];
  _RAND_3127 = {1{`RANDOM}};
  T_38110_11_uopc = _RAND_3127[8:0];
  _RAND_3128 = {1{`RANDOM}};
  T_38110_11_inst = _RAND_3128[31:0];
  _RAND_3129 = {2{`RANDOM}};
  T_38110_11_pc = _RAND_3129[39:0];
  _RAND_3130 = {1{`RANDOM}};
  T_38110_11_fu_code = _RAND_3130[7:0];
  _RAND_3131 = {1{`RANDOM}};
  T_38110_11_ctrl_br_type = _RAND_3131[3:0];
  _RAND_3132 = {1{`RANDOM}};
  T_38110_11_ctrl_op1_sel = _RAND_3132[1:0];
  _RAND_3133 = {1{`RANDOM}};
  T_38110_11_ctrl_op2_sel = _RAND_3133[2:0];
  _RAND_3134 = {1{`RANDOM}};
  T_38110_11_ctrl_imm_sel = _RAND_3134[2:0];
  _RAND_3135 = {1{`RANDOM}};
  T_38110_11_ctrl_op_fcn = _RAND_3135[3:0];
  _RAND_3136 = {1{`RANDOM}};
  T_38110_11_ctrl_fcn_dw = _RAND_3136[0:0];
  _RAND_3137 = {1{`RANDOM}};
  T_38110_11_ctrl_rf_wen = _RAND_3137[0:0];
  _RAND_3138 = {1{`RANDOM}};
  T_38110_11_ctrl_csr_cmd = _RAND_3138[2:0];
  _RAND_3139 = {1{`RANDOM}};
  T_38110_11_ctrl_is_load = _RAND_3139[0:0];
  _RAND_3140 = {1{`RANDOM}};
  T_38110_11_ctrl_is_sta = _RAND_3140[0:0];
  _RAND_3141 = {1{`RANDOM}};
  T_38110_11_ctrl_is_std = _RAND_3141[0:0];
  _RAND_3142 = {1{`RANDOM}};
  T_38110_11_wakeup_delay = _RAND_3142[1:0];
  _RAND_3143 = {1{`RANDOM}};
  T_38110_11_allocate_brtag = _RAND_3143[0:0];
  _RAND_3144 = {1{`RANDOM}};
  T_38110_11_is_br_or_jmp = _RAND_3144[0:0];
  _RAND_3145 = {1{`RANDOM}};
  T_38110_11_is_jump = _RAND_3145[0:0];
  _RAND_3146 = {1{`RANDOM}};
  T_38110_11_is_jal = _RAND_3146[0:0];
  _RAND_3147 = {1{`RANDOM}};
  T_38110_11_is_ret = _RAND_3147[0:0];
  _RAND_3148 = {1{`RANDOM}};
  T_38110_11_is_call = _RAND_3148[0:0];
  _RAND_3149 = {1{`RANDOM}};
  T_38110_11_br_mask = _RAND_3149[7:0];
  _RAND_3150 = {1{`RANDOM}};
  T_38110_11_br_tag = _RAND_3150[2:0];
  _RAND_3151 = {1{`RANDOM}};
  T_38110_11_br_prediction_bpd_predict_val = _RAND_3151[0:0];
  _RAND_3152 = {1{`RANDOM}};
  T_38110_11_br_prediction_bpd_predict_taken = _RAND_3152[0:0];
  _RAND_3153 = {1{`RANDOM}};
  T_38110_11_br_prediction_btb_hit = _RAND_3153[0:0];
  _RAND_3154 = {1{`RANDOM}};
  T_38110_11_br_prediction_btb_predicted = _RAND_3154[0:0];
  _RAND_3155 = {1{`RANDOM}};
  T_38110_11_br_prediction_is_br_or_jalr = _RAND_3155[0:0];
  _RAND_3156 = {1{`RANDOM}};
  T_38110_11_stat_brjmp_mispredicted = _RAND_3156[0:0];
  _RAND_3157 = {1{`RANDOM}};
  T_38110_11_stat_btb_made_pred = _RAND_3157[0:0];
  _RAND_3158 = {1{`RANDOM}};
  T_38110_11_stat_btb_mispredicted = _RAND_3158[0:0];
  _RAND_3159 = {1{`RANDOM}};
  T_38110_11_stat_bpd_made_pred = _RAND_3159[0:0];
  _RAND_3160 = {1{`RANDOM}};
  T_38110_11_stat_bpd_mispredicted = _RAND_3160[0:0];
  _RAND_3161 = {1{`RANDOM}};
  T_38110_11_fetch_pc_lob = _RAND_3161[2:0];
  _RAND_3162 = {1{`RANDOM}};
  T_38110_11_imm_packed = _RAND_3162[19:0];
  _RAND_3163 = {1{`RANDOM}};
  T_38110_11_csr_addr = _RAND_3163[11:0];
  _RAND_3164 = {1{`RANDOM}};
  T_38110_11_rob_idx = _RAND_3164[5:0];
  _RAND_3165 = {1{`RANDOM}};
  T_38110_11_ldq_idx = _RAND_3165[3:0];
  _RAND_3166 = {1{`RANDOM}};
  T_38110_11_stq_idx = _RAND_3166[3:0];
  _RAND_3167 = {1{`RANDOM}};
  T_38110_11_brob_idx = _RAND_3167[4:0];
  _RAND_3168 = {1{`RANDOM}};
  T_38110_11_pdst = _RAND_3168[6:0];
  _RAND_3169 = {1{`RANDOM}};
  T_38110_11_pop1 = _RAND_3169[6:0];
  _RAND_3170 = {1{`RANDOM}};
  T_38110_11_pop2 = _RAND_3170[6:0];
  _RAND_3171 = {1{`RANDOM}};
  T_38110_11_pop3 = _RAND_3171[6:0];
  _RAND_3172 = {1{`RANDOM}};
  T_38110_11_prs1_busy = _RAND_3172[0:0];
  _RAND_3173 = {1{`RANDOM}};
  T_38110_11_prs2_busy = _RAND_3173[0:0];
  _RAND_3174 = {1{`RANDOM}};
  T_38110_11_prs3_busy = _RAND_3174[0:0];
  _RAND_3175 = {1{`RANDOM}};
  T_38110_11_stale_pdst = _RAND_3175[6:0];
  _RAND_3176 = {1{`RANDOM}};
  T_38110_11_exception = _RAND_3176[0:0];
  _RAND_3177 = {2{`RANDOM}};
  T_38110_11_exc_cause = _RAND_3177[63:0];
  _RAND_3178 = {1{`RANDOM}};
  T_38110_11_bypassable = _RAND_3178[0:0];
  _RAND_3179 = {1{`RANDOM}};
  T_38110_11_mem_cmd = _RAND_3179[3:0];
  _RAND_3180 = {1{`RANDOM}};
  T_38110_11_mem_typ = _RAND_3180[2:0];
  _RAND_3181 = {1{`RANDOM}};
  T_38110_11_is_fence = _RAND_3181[0:0];
  _RAND_3182 = {1{`RANDOM}};
  T_38110_11_is_fencei = _RAND_3182[0:0];
  _RAND_3183 = {1{`RANDOM}};
  T_38110_11_is_store = _RAND_3183[0:0];
  _RAND_3184 = {1{`RANDOM}};
  T_38110_11_is_amo = _RAND_3184[0:0];
  _RAND_3185 = {1{`RANDOM}};
  T_38110_11_is_load = _RAND_3185[0:0];
  _RAND_3186 = {1{`RANDOM}};
  T_38110_11_is_unique = _RAND_3186[0:0];
  _RAND_3187 = {1{`RANDOM}};
  T_38110_11_flush_on_commit = _RAND_3187[0:0];
  _RAND_3188 = {1{`RANDOM}};
  T_38110_11_ldst = _RAND_3188[5:0];
  _RAND_3189 = {1{`RANDOM}};
  T_38110_11_lrs1 = _RAND_3189[5:0];
  _RAND_3190 = {1{`RANDOM}};
  T_38110_11_lrs2 = _RAND_3190[5:0];
  _RAND_3191 = {1{`RANDOM}};
  T_38110_11_lrs3 = _RAND_3191[5:0];
  _RAND_3192 = {1{`RANDOM}};
  T_38110_11_ldst_val = _RAND_3192[0:0];
  _RAND_3193 = {1{`RANDOM}};
  T_38110_11_dst_rtype = _RAND_3193[1:0];
  _RAND_3194 = {1{`RANDOM}};
  T_38110_11_lrs1_rtype = _RAND_3194[1:0];
  _RAND_3195 = {1{`RANDOM}};
  T_38110_11_lrs2_rtype = _RAND_3195[1:0];
  _RAND_3196 = {1{`RANDOM}};
  T_38110_11_frs3_en = _RAND_3196[0:0];
  _RAND_3197 = {1{`RANDOM}};
  T_38110_11_fp_val = _RAND_3197[0:0];
  _RAND_3198 = {1{`RANDOM}};
  T_38110_11_fp_single = _RAND_3198[0:0];
  _RAND_3199 = {1{`RANDOM}};
  T_38110_11_xcpt_if = _RAND_3199[0:0];
  _RAND_3200 = {1{`RANDOM}};
  T_38110_11_replay_if = _RAND_3200[0:0];
  _RAND_3201 = {2{`RANDOM}};
  T_38110_11_debug_wdata = _RAND_3201[63:0];
  _RAND_3202 = {1{`RANDOM}};
  T_38110_11_debug_events_fetch_seq = _RAND_3202[31:0];
  _RAND_3203 = {1{`RANDOM}};
  T_38110_12_valid = _RAND_3203[0:0];
  _RAND_3204 = {1{`RANDOM}};
  T_38110_12_iw_state = _RAND_3204[1:0];
  _RAND_3205 = {1{`RANDOM}};
  T_38110_12_uopc = _RAND_3205[8:0];
  _RAND_3206 = {1{`RANDOM}};
  T_38110_12_inst = _RAND_3206[31:0];
  _RAND_3207 = {2{`RANDOM}};
  T_38110_12_pc = _RAND_3207[39:0];
  _RAND_3208 = {1{`RANDOM}};
  T_38110_12_fu_code = _RAND_3208[7:0];
  _RAND_3209 = {1{`RANDOM}};
  T_38110_12_ctrl_br_type = _RAND_3209[3:0];
  _RAND_3210 = {1{`RANDOM}};
  T_38110_12_ctrl_op1_sel = _RAND_3210[1:0];
  _RAND_3211 = {1{`RANDOM}};
  T_38110_12_ctrl_op2_sel = _RAND_3211[2:0];
  _RAND_3212 = {1{`RANDOM}};
  T_38110_12_ctrl_imm_sel = _RAND_3212[2:0];
  _RAND_3213 = {1{`RANDOM}};
  T_38110_12_ctrl_op_fcn = _RAND_3213[3:0];
  _RAND_3214 = {1{`RANDOM}};
  T_38110_12_ctrl_fcn_dw = _RAND_3214[0:0];
  _RAND_3215 = {1{`RANDOM}};
  T_38110_12_ctrl_rf_wen = _RAND_3215[0:0];
  _RAND_3216 = {1{`RANDOM}};
  T_38110_12_ctrl_csr_cmd = _RAND_3216[2:0];
  _RAND_3217 = {1{`RANDOM}};
  T_38110_12_ctrl_is_load = _RAND_3217[0:0];
  _RAND_3218 = {1{`RANDOM}};
  T_38110_12_ctrl_is_sta = _RAND_3218[0:0];
  _RAND_3219 = {1{`RANDOM}};
  T_38110_12_ctrl_is_std = _RAND_3219[0:0];
  _RAND_3220 = {1{`RANDOM}};
  T_38110_12_wakeup_delay = _RAND_3220[1:0];
  _RAND_3221 = {1{`RANDOM}};
  T_38110_12_allocate_brtag = _RAND_3221[0:0];
  _RAND_3222 = {1{`RANDOM}};
  T_38110_12_is_br_or_jmp = _RAND_3222[0:0];
  _RAND_3223 = {1{`RANDOM}};
  T_38110_12_is_jump = _RAND_3223[0:0];
  _RAND_3224 = {1{`RANDOM}};
  T_38110_12_is_jal = _RAND_3224[0:0];
  _RAND_3225 = {1{`RANDOM}};
  T_38110_12_is_ret = _RAND_3225[0:0];
  _RAND_3226 = {1{`RANDOM}};
  T_38110_12_is_call = _RAND_3226[0:0];
  _RAND_3227 = {1{`RANDOM}};
  T_38110_12_br_mask = _RAND_3227[7:0];
  _RAND_3228 = {1{`RANDOM}};
  T_38110_12_br_tag = _RAND_3228[2:0];
  _RAND_3229 = {1{`RANDOM}};
  T_38110_12_br_prediction_bpd_predict_val = _RAND_3229[0:0];
  _RAND_3230 = {1{`RANDOM}};
  T_38110_12_br_prediction_bpd_predict_taken = _RAND_3230[0:0];
  _RAND_3231 = {1{`RANDOM}};
  T_38110_12_br_prediction_btb_hit = _RAND_3231[0:0];
  _RAND_3232 = {1{`RANDOM}};
  T_38110_12_br_prediction_btb_predicted = _RAND_3232[0:0];
  _RAND_3233 = {1{`RANDOM}};
  T_38110_12_br_prediction_is_br_or_jalr = _RAND_3233[0:0];
  _RAND_3234 = {1{`RANDOM}};
  T_38110_12_stat_brjmp_mispredicted = _RAND_3234[0:0];
  _RAND_3235 = {1{`RANDOM}};
  T_38110_12_stat_btb_made_pred = _RAND_3235[0:0];
  _RAND_3236 = {1{`RANDOM}};
  T_38110_12_stat_btb_mispredicted = _RAND_3236[0:0];
  _RAND_3237 = {1{`RANDOM}};
  T_38110_12_stat_bpd_made_pred = _RAND_3237[0:0];
  _RAND_3238 = {1{`RANDOM}};
  T_38110_12_stat_bpd_mispredicted = _RAND_3238[0:0];
  _RAND_3239 = {1{`RANDOM}};
  T_38110_12_fetch_pc_lob = _RAND_3239[2:0];
  _RAND_3240 = {1{`RANDOM}};
  T_38110_12_imm_packed = _RAND_3240[19:0];
  _RAND_3241 = {1{`RANDOM}};
  T_38110_12_csr_addr = _RAND_3241[11:0];
  _RAND_3242 = {1{`RANDOM}};
  T_38110_12_rob_idx = _RAND_3242[5:0];
  _RAND_3243 = {1{`RANDOM}};
  T_38110_12_ldq_idx = _RAND_3243[3:0];
  _RAND_3244 = {1{`RANDOM}};
  T_38110_12_stq_idx = _RAND_3244[3:0];
  _RAND_3245 = {1{`RANDOM}};
  T_38110_12_brob_idx = _RAND_3245[4:0];
  _RAND_3246 = {1{`RANDOM}};
  T_38110_12_pdst = _RAND_3246[6:0];
  _RAND_3247 = {1{`RANDOM}};
  T_38110_12_pop1 = _RAND_3247[6:0];
  _RAND_3248 = {1{`RANDOM}};
  T_38110_12_pop2 = _RAND_3248[6:0];
  _RAND_3249 = {1{`RANDOM}};
  T_38110_12_pop3 = _RAND_3249[6:0];
  _RAND_3250 = {1{`RANDOM}};
  T_38110_12_prs1_busy = _RAND_3250[0:0];
  _RAND_3251 = {1{`RANDOM}};
  T_38110_12_prs2_busy = _RAND_3251[0:0];
  _RAND_3252 = {1{`RANDOM}};
  T_38110_12_prs3_busy = _RAND_3252[0:0];
  _RAND_3253 = {1{`RANDOM}};
  T_38110_12_stale_pdst = _RAND_3253[6:0];
  _RAND_3254 = {1{`RANDOM}};
  T_38110_12_exception = _RAND_3254[0:0];
  _RAND_3255 = {2{`RANDOM}};
  T_38110_12_exc_cause = _RAND_3255[63:0];
  _RAND_3256 = {1{`RANDOM}};
  T_38110_12_bypassable = _RAND_3256[0:0];
  _RAND_3257 = {1{`RANDOM}};
  T_38110_12_mem_cmd = _RAND_3257[3:0];
  _RAND_3258 = {1{`RANDOM}};
  T_38110_12_mem_typ = _RAND_3258[2:0];
  _RAND_3259 = {1{`RANDOM}};
  T_38110_12_is_fence = _RAND_3259[0:0];
  _RAND_3260 = {1{`RANDOM}};
  T_38110_12_is_fencei = _RAND_3260[0:0];
  _RAND_3261 = {1{`RANDOM}};
  T_38110_12_is_store = _RAND_3261[0:0];
  _RAND_3262 = {1{`RANDOM}};
  T_38110_12_is_amo = _RAND_3262[0:0];
  _RAND_3263 = {1{`RANDOM}};
  T_38110_12_is_load = _RAND_3263[0:0];
  _RAND_3264 = {1{`RANDOM}};
  T_38110_12_is_unique = _RAND_3264[0:0];
  _RAND_3265 = {1{`RANDOM}};
  T_38110_12_flush_on_commit = _RAND_3265[0:0];
  _RAND_3266 = {1{`RANDOM}};
  T_38110_12_ldst = _RAND_3266[5:0];
  _RAND_3267 = {1{`RANDOM}};
  T_38110_12_lrs1 = _RAND_3267[5:0];
  _RAND_3268 = {1{`RANDOM}};
  T_38110_12_lrs2 = _RAND_3268[5:0];
  _RAND_3269 = {1{`RANDOM}};
  T_38110_12_lrs3 = _RAND_3269[5:0];
  _RAND_3270 = {1{`RANDOM}};
  T_38110_12_ldst_val = _RAND_3270[0:0];
  _RAND_3271 = {1{`RANDOM}};
  T_38110_12_dst_rtype = _RAND_3271[1:0];
  _RAND_3272 = {1{`RANDOM}};
  T_38110_12_lrs1_rtype = _RAND_3272[1:0];
  _RAND_3273 = {1{`RANDOM}};
  T_38110_12_lrs2_rtype = _RAND_3273[1:0];
  _RAND_3274 = {1{`RANDOM}};
  T_38110_12_frs3_en = _RAND_3274[0:0];
  _RAND_3275 = {1{`RANDOM}};
  T_38110_12_fp_val = _RAND_3275[0:0];
  _RAND_3276 = {1{`RANDOM}};
  T_38110_12_fp_single = _RAND_3276[0:0];
  _RAND_3277 = {1{`RANDOM}};
  T_38110_12_xcpt_if = _RAND_3277[0:0];
  _RAND_3278 = {1{`RANDOM}};
  T_38110_12_replay_if = _RAND_3278[0:0];
  _RAND_3279 = {2{`RANDOM}};
  T_38110_12_debug_wdata = _RAND_3279[63:0];
  _RAND_3280 = {1{`RANDOM}};
  T_38110_12_debug_events_fetch_seq = _RAND_3280[31:0];
  _RAND_3281 = {1{`RANDOM}};
  T_38110_13_valid = _RAND_3281[0:0];
  _RAND_3282 = {1{`RANDOM}};
  T_38110_13_iw_state = _RAND_3282[1:0];
  _RAND_3283 = {1{`RANDOM}};
  T_38110_13_uopc = _RAND_3283[8:0];
  _RAND_3284 = {1{`RANDOM}};
  T_38110_13_inst = _RAND_3284[31:0];
  _RAND_3285 = {2{`RANDOM}};
  T_38110_13_pc = _RAND_3285[39:0];
  _RAND_3286 = {1{`RANDOM}};
  T_38110_13_fu_code = _RAND_3286[7:0];
  _RAND_3287 = {1{`RANDOM}};
  T_38110_13_ctrl_br_type = _RAND_3287[3:0];
  _RAND_3288 = {1{`RANDOM}};
  T_38110_13_ctrl_op1_sel = _RAND_3288[1:0];
  _RAND_3289 = {1{`RANDOM}};
  T_38110_13_ctrl_op2_sel = _RAND_3289[2:0];
  _RAND_3290 = {1{`RANDOM}};
  T_38110_13_ctrl_imm_sel = _RAND_3290[2:0];
  _RAND_3291 = {1{`RANDOM}};
  T_38110_13_ctrl_op_fcn = _RAND_3291[3:0];
  _RAND_3292 = {1{`RANDOM}};
  T_38110_13_ctrl_fcn_dw = _RAND_3292[0:0];
  _RAND_3293 = {1{`RANDOM}};
  T_38110_13_ctrl_rf_wen = _RAND_3293[0:0];
  _RAND_3294 = {1{`RANDOM}};
  T_38110_13_ctrl_csr_cmd = _RAND_3294[2:0];
  _RAND_3295 = {1{`RANDOM}};
  T_38110_13_ctrl_is_load = _RAND_3295[0:0];
  _RAND_3296 = {1{`RANDOM}};
  T_38110_13_ctrl_is_sta = _RAND_3296[0:0];
  _RAND_3297 = {1{`RANDOM}};
  T_38110_13_ctrl_is_std = _RAND_3297[0:0];
  _RAND_3298 = {1{`RANDOM}};
  T_38110_13_wakeup_delay = _RAND_3298[1:0];
  _RAND_3299 = {1{`RANDOM}};
  T_38110_13_allocate_brtag = _RAND_3299[0:0];
  _RAND_3300 = {1{`RANDOM}};
  T_38110_13_is_br_or_jmp = _RAND_3300[0:0];
  _RAND_3301 = {1{`RANDOM}};
  T_38110_13_is_jump = _RAND_3301[0:0];
  _RAND_3302 = {1{`RANDOM}};
  T_38110_13_is_jal = _RAND_3302[0:0];
  _RAND_3303 = {1{`RANDOM}};
  T_38110_13_is_ret = _RAND_3303[0:0];
  _RAND_3304 = {1{`RANDOM}};
  T_38110_13_is_call = _RAND_3304[0:0];
  _RAND_3305 = {1{`RANDOM}};
  T_38110_13_br_mask = _RAND_3305[7:0];
  _RAND_3306 = {1{`RANDOM}};
  T_38110_13_br_tag = _RAND_3306[2:0];
  _RAND_3307 = {1{`RANDOM}};
  T_38110_13_br_prediction_bpd_predict_val = _RAND_3307[0:0];
  _RAND_3308 = {1{`RANDOM}};
  T_38110_13_br_prediction_bpd_predict_taken = _RAND_3308[0:0];
  _RAND_3309 = {1{`RANDOM}};
  T_38110_13_br_prediction_btb_hit = _RAND_3309[0:0];
  _RAND_3310 = {1{`RANDOM}};
  T_38110_13_br_prediction_btb_predicted = _RAND_3310[0:0];
  _RAND_3311 = {1{`RANDOM}};
  T_38110_13_br_prediction_is_br_or_jalr = _RAND_3311[0:0];
  _RAND_3312 = {1{`RANDOM}};
  T_38110_13_stat_brjmp_mispredicted = _RAND_3312[0:0];
  _RAND_3313 = {1{`RANDOM}};
  T_38110_13_stat_btb_made_pred = _RAND_3313[0:0];
  _RAND_3314 = {1{`RANDOM}};
  T_38110_13_stat_btb_mispredicted = _RAND_3314[0:0];
  _RAND_3315 = {1{`RANDOM}};
  T_38110_13_stat_bpd_made_pred = _RAND_3315[0:0];
  _RAND_3316 = {1{`RANDOM}};
  T_38110_13_stat_bpd_mispredicted = _RAND_3316[0:0];
  _RAND_3317 = {1{`RANDOM}};
  T_38110_13_fetch_pc_lob = _RAND_3317[2:0];
  _RAND_3318 = {1{`RANDOM}};
  T_38110_13_imm_packed = _RAND_3318[19:0];
  _RAND_3319 = {1{`RANDOM}};
  T_38110_13_csr_addr = _RAND_3319[11:0];
  _RAND_3320 = {1{`RANDOM}};
  T_38110_13_rob_idx = _RAND_3320[5:0];
  _RAND_3321 = {1{`RANDOM}};
  T_38110_13_ldq_idx = _RAND_3321[3:0];
  _RAND_3322 = {1{`RANDOM}};
  T_38110_13_stq_idx = _RAND_3322[3:0];
  _RAND_3323 = {1{`RANDOM}};
  T_38110_13_brob_idx = _RAND_3323[4:0];
  _RAND_3324 = {1{`RANDOM}};
  T_38110_13_pdst = _RAND_3324[6:0];
  _RAND_3325 = {1{`RANDOM}};
  T_38110_13_pop1 = _RAND_3325[6:0];
  _RAND_3326 = {1{`RANDOM}};
  T_38110_13_pop2 = _RAND_3326[6:0];
  _RAND_3327 = {1{`RANDOM}};
  T_38110_13_pop3 = _RAND_3327[6:0];
  _RAND_3328 = {1{`RANDOM}};
  T_38110_13_prs1_busy = _RAND_3328[0:0];
  _RAND_3329 = {1{`RANDOM}};
  T_38110_13_prs2_busy = _RAND_3329[0:0];
  _RAND_3330 = {1{`RANDOM}};
  T_38110_13_prs3_busy = _RAND_3330[0:0];
  _RAND_3331 = {1{`RANDOM}};
  T_38110_13_stale_pdst = _RAND_3331[6:0];
  _RAND_3332 = {1{`RANDOM}};
  T_38110_13_exception = _RAND_3332[0:0];
  _RAND_3333 = {2{`RANDOM}};
  T_38110_13_exc_cause = _RAND_3333[63:0];
  _RAND_3334 = {1{`RANDOM}};
  T_38110_13_bypassable = _RAND_3334[0:0];
  _RAND_3335 = {1{`RANDOM}};
  T_38110_13_mem_cmd = _RAND_3335[3:0];
  _RAND_3336 = {1{`RANDOM}};
  T_38110_13_mem_typ = _RAND_3336[2:0];
  _RAND_3337 = {1{`RANDOM}};
  T_38110_13_is_fence = _RAND_3337[0:0];
  _RAND_3338 = {1{`RANDOM}};
  T_38110_13_is_fencei = _RAND_3338[0:0];
  _RAND_3339 = {1{`RANDOM}};
  T_38110_13_is_store = _RAND_3339[0:0];
  _RAND_3340 = {1{`RANDOM}};
  T_38110_13_is_amo = _RAND_3340[0:0];
  _RAND_3341 = {1{`RANDOM}};
  T_38110_13_is_load = _RAND_3341[0:0];
  _RAND_3342 = {1{`RANDOM}};
  T_38110_13_is_unique = _RAND_3342[0:0];
  _RAND_3343 = {1{`RANDOM}};
  T_38110_13_flush_on_commit = _RAND_3343[0:0];
  _RAND_3344 = {1{`RANDOM}};
  T_38110_13_ldst = _RAND_3344[5:0];
  _RAND_3345 = {1{`RANDOM}};
  T_38110_13_lrs1 = _RAND_3345[5:0];
  _RAND_3346 = {1{`RANDOM}};
  T_38110_13_lrs2 = _RAND_3346[5:0];
  _RAND_3347 = {1{`RANDOM}};
  T_38110_13_lrs3 = _RAND_3347[5:0];
  _RAND_3348 = {1{`RANDOM}};
  T_38110_13_ldst_val = _RAND_3348[0:0];
  _RAND_3349 = {1{`RANDOM}};
  T_38110_13_dst_rtype = _RAND_3349[1:0];
  _RAND_3350 = {1{`RANDOM}};
  T_38110_13_lrs1_rtype = _RAND_3350[1:0];
  _RAND_3351 = {1{`RANDOM}};
  T_38110_13_lrs2_rtype = _RAND_3351[1:0];
  _RAND_3352 = {1{`RANDOM}};
  T_38110_13_frs3_en = _RAND_3352[0:0];
  _RAND_3353 = {1{`RANDOM}};
  T_38110_13_fp_val = _RAND_3353[0:0];
  _RAND_3354 = {1{`RANDOM}};
  T_38110_13_fp_single = _RAND_3354[0:0];
  _RAND_3355 = {1{`RANDOM}};
  T_38110_13_xcpt_if = _RAND_3355[0:0];
  _RAND_3356 = {1{`RANDOM}};
  T_38110_13_replay_if = _RAND_3356[0:0];
  _RAND_3357 = {2{`RANDOM}};
  T_38110_13_debug_wdata = _RAND_3357[63:0];
  _RAND_3358 = {1{`RANDOM}};
  T_38110_13_debug_events_fetch_seq = _RAND_3358[31:0];
  _RAND_3359 = {1{`RANDOM}};
  T_38110_14_valid = _RAND_3359[0:0];
  _RAND_3360 = {1{`RANDOM}};
  T_38110_14_iw_state = _RAND_3360[1:0];
  _RAND_3361 = {1{`RANDOM}};
  T_38110_14_uopc = _RAND_3361[8:0];
  _RAND_3362 = {1{`RANDOM}};
  T_38110_14_inst = _RAND_3362[31:0];
  _RAND_3363 = {2{`RANDOM}};
  T_38110_14_pc = _RAND_3363[39:0];
  _RAND_3364 = {1{`RANDOM}};
  T_38110_14_fu_code = _RAND_3364[7:0];
  _RAND_3365 = {1{`RANDOM}};
  T_38110_14_ctrl_br_type = _RAND_3365[3:0];
  _RAND_3366 = {1{`RANDOM}};
  T_38110_14_ctrl_op1_sel = _RAND_3366[1:0];
  _RAND_3367 = {1{`RANDOM}};
  T_38110_14_ctrl_op2_sel = _RAND_3367[2:0];
  _RAND_3368 = {1{`RANDOM}};
  T_38110_14_ctrl_imm_sel = _RAND_3368[2:0];
  _RAND_3369 = {1{`RANDOM}};
  T_38110_14_ctrl_op_fcn = _RAND_3369[3:0];
  _RAND_3370 = {1{`RANDOM}};
  T_38110_14_ctrl_fcn_dw = _RAND_3370[0:0];
  _RAND_3371 = {1{`RANDOM}};
  T_38110_14_ctrl_rf_wen = _RAND_3371[0:0];
  _RAND_3372 = {1{`RANDOM}};
  T_38110_14_ctrl_csr_cmd = _RAND_3372[2:0];
  _RAND_3373 = {1{`RANDOM}};
  T_38110_14_ctrl_is_load = _RAND_3373[0:0];
  _RAND_3374 = {1{`RANDOM}};
  T_38110_14_ctrl_is_sta = _RAND_3374[0:0];
  _RAND_3375 = {1{`RANDOM}};
  T_38110_14_ctrl_is_std = _RAND_3375[0:0];
  _RAND_3376 = {1{`RANDOM}};
  T_38110_14_wakeup_delay = _RAND_3376[1:0];
  _RAND_3377 = {1{`RANDOM}};
  T_38110_14_allocate_brtag = _RAND_3377[0:0];
  _RAND_3378 = {1{`RANDOM}};
  T_38110_14_is_br_or_jmp = _RAND_3378[0:0];
  _RAND_3379 = {1{`RANDOM}};
  T_38110_14_is_jump = _RAND_3379[0:0];
  _RAND_3380 = {1{`RANDOM}};
  T_38110_14_is_jal = _RAND_3380[0:0];
  _RAND_3381 = {1{`RANDOM}};
  T_38110_14_is_ret = _RAND_3381[0:0];
  _RAND_3382 = {1{`RANDOM}};
  T_38110_14_is_call = _RAND_3382[0:0];
  _RAND_3383 = {1{`RANDOM}};
  T_38110_14_br_mask = _RAND_3383[7:0];
  _RAND_3384 = {1{`RANDOM}};
  T_38110_14_br_tag = _RAND_3384[2:0];
  _RAND_3385 = {1{`RANDOM}};
  T_38110_14_br_prediction_bpd_predict_val = _RAND_3385[0:0];
  _RAND_3386 = {1{`RANDOM}};
  T_38110_14_br_prediction_bpd_predict_taken = _RAND_3386[0:0];
  _RAND_3387 = {1{`RANDOM}};
  T_38110_14_br_prediction_btb_hit = _RAND_3387[0:0];
  _RAND_3388 = {1{`RANDOM}};
  T_38110_14_br_prediction_btb_predicted = _RAND_3388[0:0];
  _RAND_3389 = {1{`RANDOM}};
  T_38110_14_br_prediction_is_br_or_jalr = _RAND_3389[0:0];
  _RAND_3390 = {1{`RANDOM}};
  T_38110_14_stat_brjmp_mispredicted = _RAND_3390[0:0];
  _RAND_3391 = {1{`RANDOM}};
  T_38110_14_stat_btb_made_pred = _RAND_3391[0:0];
  _RAND_3392 = {1{`RANDOM}};
  T_38110_14_stat_btb_mispredicted = _RAND_3392[0:0];
  _RAND_3393 = {1{`RANDOM}};
  T_38110_14_stat_bpd_made_pred = _RAND_3393[0:0];
  _RAND_3394 = {1{`RANDOM}};
  T_38110_14_stat_bpd_mispredicted = _RAND_3394[0:0];
  _RAND_3395 = {1{`RANDOM}};
  T_38110_14_fetch_pc_lob = _RAND_3395[2:0];
  _RAND_3396 = {1{`RANDOM}};
  T_38110_14_imm_packed = _RAND_3396[19:0];
  _RAND_3397 = {1{`RANDOM}};
  T_38110_14_csr_addr = _RAND_3397[11:0];
  _RAND_3398 = {1{`RANDOM}};
  T_38110_14_rob_idx = _RAND_3398[5:0];
  _RAND_3399 = {1{`RANDOM}};
  T_38110_14_ldq_idx = _RAND_3399[3:0];
  _RAND_3400 = {1{`RANDOM}};
  T_38110_14_stq_idx = _RAND_3400[3:0];
  _RAND_3401 = {1{`RANDOM}};
  T_38110_14_brob_idx = _RAND_3401[4:0];
  _RAND_3402 = {1{`RANDOM}};
  T_38110_14_pdst = _RAND_3402[6:0];
  _RAND_3403 = {1{`RANDOM}};
  T_38110_14_pop1 = _RAND_3403[6:0];
  _RAND_3404 = {1{`RANDOM}};
  T_38110_14_pop2 = _RAND_3404[6:0];
  _RAND_3405 = {1{`RANDOM}};
  T_38110_14_pop3 = _RAND_3405[6:0];
  _RAND_3406 = {1{`RANDOM}};
  T_38110_14_prs1_busy = _RAND_3406[0:0];
  _RAND_3407 = {1{`RANDOM}};
  T_38110_14_prs2_busy = _RAND_3407[0:0];
  _RAND_3408 = {1{`RANDOM}};
  T_38110_14_prs3_busy = _RAND_3408[0:0];
  _RAND_3409 = {1{`RANDOM}};
  T_38110_14_stale_pdst = _RAND_3409[6:0];
  _RAND_3410 = {1{`RANDOM}};
  T_38110_14_exception = _RAND_3410[0:0];
  _RAND_3411 = {2{`RANDOM}};
  T_38110_14_exc_cause = _RAND_3411[63:0];
  _RAND_3412 = {1{`RANDOM}};
  T_38110_14_bypassable = _RAND_3412[0:0];
  _RAND_3413 = {1{`RANDOM}};
  T_38110_14_mem_cmd = _RAND_3413[3:0];
  _RAND_3414 = {1{`RANDOM}};
  T_38110_14_mem_typ = _RAND_3414[2:0];
  _RAND_3415 = {1{`RANDOM}};
  T_38110_14_is_fence = _RAND_3415[0:0];
  _RAND_3416 = {1{`RANDOM}};
  T_38110_14_is_fencei = _RAND_3416[0:0];
  _RAND_3417 = {1{`RANDOM}};
  T_38110_14_is_store = _RAND_3417[0:0];
  _RAND_3418 = {1{`RANDOM}};
  T_38110_14_is_amo = _RAND_3418[0:0];
  _RAND_3419 = {1{`RANDOM}};
  T_38110_14_is_load = _RAND_3419[0:0];
  _RAND_3420 = {1{`RANDOM}};
  T_38110_14_is_unique = _RAND_3420[0:0];
  _RAND_3421 = {1{`RANDOM}};
  T_38110_14_flush_on_commit = _RAND_3421[0:0];
  _RAND_3422 = {1{`RANDOM}};
  T_38110_14_ldst = _RAND_3422[5:0];
  _RAND_3423 = {1{`RANDOM}};
  T_38110_14_lrs1 = _RAND_3423[5:0];
  _RAND_3424 = {1{`RANDOM}};
  T_38110_14_lrs2 = _RAND_3424[5:0];
  _RAND_3425 = {1{`RANDOM}};
  T_38110_14_lrs3 = _RAND_3425[5:0];
  _RAND_3426 = {1{`RANDOM}};
  T_38110_14_ldst_val = _RAND_3426[0:0];
  _RAND_3427 = {1{`RANDOM}};
  T_38110_14_dst_rtype = _RAND_3427[1:0];
  _RAND_3428 = {1{`RANDOM}};
  T_38110_14_lrs1_rtype = _RAND_3428[1:0];
  _RAND_3429 = {1{`RANDOM}};
  T_38110_14_lrs2_rtype = _RAND_3429[1:0];
  _RAND_3430 = {1{`RANDOM}};
  T_38110_14_frs3_en = _RAND_3430[0:0];
  _RAND_3431 = {1{`RANDOM}};
  T_38110_14_fp_val = _RAND_3431[0:0];
  _RAND_3432 = {1{`RANDOM}};
  T_38110_14_fp_single = _RAND_3432[0:0];
  _RAND_3433 = {1{`RANDOM}};
  T_38110_14_xcpt_if = _RAND_3433[0:0];
  _RAND_3434 = {1{`RANDOM}};
  T_38110_14_replay_if = _RAND_3434[0:0];
  _RAND_3435 = {2{`RANDOM}};
  T_38110_14_debug_wdata = _RAND_3435[63:0];
  _RAND_3436 = {1{`RANDOM}};
  T_38110_14_debug_events_fetch_seq = _RAND_3436[31:0];
  _RAND_3437 = {1{`RANDOM}};
  T_38110_15_valid = _RAND_3437[0:0];
  _RAND_3438 = {1{`RANDOM}};
  T_38110_15_iw_state = _RAND_3438[1:0];
  _RAND_3439 = {1{`RANDOM}};
  T_38110_15_uopc = _RAND_3439[8:0];
  _RAND_3440 = {1{`RANDOM}};
  T_38110_15_inst = _RAND_3440[31:0];
  _RAND_3441 = {2{`RANDOM}};
  T_38110_15_pc = _RAND_3441[39:0];
  _RAND_3442 = {1{`RANDOM}};
  T_38110_15_fu_code = _RAND_3442[7:0];
  _RAND_3443 = {1{`RANDOM}};
  T_38110_15_ctrl_br_type = _RAND_3443[3:0];
  _RAND_3444 = {1{`RANDOM}};
  T_38110_15_ctrl_op1_sel = _RAND_3444[1:0];
  _RAND_3445 = {1{`RANDOM}};
  T_38110_15_ctrl_op2_sel = _RAND_3445[2:0];
  _RAND_3446 = {1{`RANDOM}};
  T_38110_15_ctrl_imm_sel = _RAND_3446[2:0];
  _RAND_3447 = {1{`RANDOM}};
  T_38110_15_ctrl_op_fcn = _RAND_3447[3:0];
  _RAND_3448 = {1{`RANDOM}};
  T_38110_15_ctrl_fcn_dw = _RAND_3448[0:0];
  _RAND_3449 = {1{`RANDOM}};
  T_38110_15_ctrl_rf_wen = _RAND_3449[0:0];
  _RAND_3450 = {1{`RANDOM}};
  T_38110_15_ctrl_csr_cmd = _RAND_3450[2:0];
  _RAND_3451 = {1{`RANDOM}};
  T_38110_15_ctrl_is_load = _RAND_3451[0:0];
  _RAND_3452 = {1{`RANDOM}};
  T_38110_15_ctrl_is_sta = _RAND_3452[0:0];
  _RAND_3453 = {1{`RANDOM}};
  T_38110_15_ctrl_is_std = _RAND_3453[0:0];
  _RAND_3454 = {1{`RANDOM}};
  T_38110_15_wakeup_delay = _RAND_3454[1:0];
  _RAND_3455 = {1{`RANDOM}};
  T_38110_15_allocate_brtag = _RAND_3455[0:0];
  _RAND_3456 = {1{`RANDOM}};
  T_38110_15_is_br_or_jmp = _RAND_3456[0:0];
  _RAND_3457 = {1{`RANDOM}};
  T_38110_15_is_jump = _RAND_3457[0:0];
  _RAND_3458 = {1{`RANDOM}};
  T_38110_15_is_jal = _RAND_3458[0:0];
  _RAND_3459 = {1{`RANDOM}};
  T_38110_15_is_ret = _RAND_3459[0:0];
  _RAND_3460 = {1{`RANDOM}};
  T_38110_15_is_call = _RAND_3460[0:0];
  _RAND_3461 = {1{`RANDOM}};
  T_38110_15_br_mask = _RAND_3461[7:0];
  _RAND_3462 = {1{`RANDOM}};
  T_38110_15_br_tag = _RAND_3462[2:0];
  _RAND_3463 = {1{`RANDOM}};
  T_38110_15_br_prediction_bpd_predict_val = _RAND_3463[0:0];
  _RAND_3464 = {1{`RANDOM}};
  T_38110_15_br_prediction_bpd_predict_taken = _RAND_3464[0:0];
  _RAND_3465 = {1{`RANDOM}};
  T_38110_15_br_prediction_btb_hit = _RAND_3465[0:0];
  _RAND_3466 = {1{`RANDOM}};
  T_38110_15_br_prediction_btb_predicted = _RAND_3466[0:0];
  _RAND_3467 = {1{`RANDOM}};
  T_38110_15_br_prediction_is_br_or_jalr = _RAND_3467[0:0];
  _RAND_3468 = {1{`RANDOM}};
  T_38110_15_stat_brjmp_mispredicted = _RAND_3468[0:0];
  _RAND_3469 = {1{`RANDOM}};
  T_38110_15_stat_btb_made_pred = _RAND_3469[0:0];
  _RAND_3470 = {1{`RANDOM}};
  T_38110_15_stat_btb_mispredicted = _RAND_3470[0:0];
  _RAND_3471 = {1{`RANDOM}};
  T_38110_15_stat_bpd_made_pred = _RAND_3471[0:0];
  _RAND_3472 = {1{`RANDOM}};
  T_38110_15_stat_bpd_mispredicted = _RAND_3472[0:0];
  _RAND_3473 = {1{`RANDOM}};
  T_38110_15_fetch_pc_lob = _RAND_3473[2:0];
  _RAND_3474 = {1{`RANDOM}};
  T_38110_15_imm_packed = _RAND_3474[19:0];
  _RAND_3475 = {1{`RANDOM}};
  T_38110_15_csr_addr = _RAND_3475[11:0];
  _RAND_3476 = {1{`RANDOM}};
  T_38110_15_rob_idx = _RAND_3476[5:0];
  _RAND_3477 = {1{`RANDOM}};
  T_38110_15_ldq_idx = _RAND_3477[3:0];
  _RAND_3478 = {1{`RANDOM}};
  T_38110_15_stq_idx = _RAND_3478[3:0];
  _RAND_3479 = {1{`RANDOM}};
  T_38110_15_brob_idx = _RAND_3479[4:0];
  _RAND_3480 = {1{`RANDOM}};
  T_38110_15_pdst = _RAND_3480[6:0];
  _RAND_3481 = {1{`RANDOM}};
  T_38110_15_pop1 = _RAND_3481[6:0];
  _RAND_3482 = {1{`RANDOM}};
  T_38110_15_pop2 = _RAND_3482[6:0];
  _RAND_3483 = {1{`RANDOM}};
  T_38110_15_pop3 = _RAND_3483[6:0];
  _RAND_3484 = {1{`RANDOM}};
  T_38110_15_prs1_busy = _RAND_3484[0:0];
  _RAND_3485 = {1{`RANDOM}};
  T_38110_15_prs2_busy = _RAND_3485[0:0];
  _RAND_3486 = {1{`RANDOM}};
  T_38110_15_prs3_busy = _RAND_3486[0:0];
  _RAND_3487 = {1{`RANDOM}};
  T_38110_15_stale_pdst = _RAND_3487[6:0];
  _RAND_3488 = {1{`RANDOM}};
  T_38110_15_exception = _RAND_3488[0:0];
  _RAND_3489 = {2{`RANDOM}};
  T_38110_15_exc_cause = _RAND_3489[63:0];
  _RAND_3490 = {1{`RANDOM}};
  T_38110_15_bypassable = _RAND_3490[0:0];
  _RAND_3491 = {1{`RANDOM}};
  T_38110_15_mem_cmd = _RAND_3491[3:0];
  _RAND_3492 = {1{`RANDOM}};
  T_38110_15_mem_typ = _RAND_3492[2:0];
  _RAND_3493 = {1{`RANDOM}};
  T_38110_15_is_fence = _RAND_3493[0:0];
  _RAND_3494 = {1{`RANDOM}};
  T_38110_15_is_fencei = _RAND_3494[0:0];
  _RAND_3495 = {1{`RANDOM}};
  T_38110_15_is_store = _RAND_3495[0:0];
  _RAND_3496 = {1{`RANDOM}};
  T_38110_15_is_amo = _RAND_3496[0:0];
  _RAND_3497 = {1{`RANDOM}};
  T_38110_15_is_load = _RAND_3497[0:0];
  _RAND_3498 = {1{`RANDOM}};
  T_38110_15_is_unique = _RAND_3498[0:0];
  _RAND_3499 = {1{`RANDOM}};
  T_38110_15_flush_on_commit = _RAND_3499[0:0];
  _RAND_3500 = {1{`RANDOM}};
  T_38110_15_ldst = _RAND_3500[5:0];
  _RAND_3501 = {1{`RANDOM}};
  T_38110_15_lrs1 = _RAND_3501[5:0];
  _RAND_3502 = {1{`RANDOM}};
  T_38110_15_lrs2 = _RAND_3502[5:0];
  _RAND_3503 = {1{`RANDOM}};
  T_38110_15_lrs3 = _RAND_3503[5:0];
  _RAND_3504 = {1{`RANDOM}};
  T_38110_15_ldst_val = _RAND_3504[0:0];
  _RAND_3505 = {1{`RANDOM}};
  T_38110_15_dst_rtype = _RAND_3505[1:0];
  _RAND_3506 = {1{`RANDOM}};
  T_38110_15_lrs1_rtype = _RAND_3506[1:0];
  _RAND_3507 = {1{`RANDOM}};
  T_38110_15_lrs2_rtype = _RAND_3507[1:0];
  _RAND_3508 = {1{`RANDOM}};
  T_38110_15_frs3_en = _RAND_3508[0:0];
  _RAND_3509 = {1{`RANDOM}};
  T_38110_15_fp_val = _RAND_3509[0:0];
  _RAND_3510 = {1{`RANDOM}};
  T_38110_15_fp_single = _RAND_3510[0:0];
  _RAND_3511 = {1{`RANDOM}};
  T_38110_15_xcpt_if = _RAND_3511[0:0];
  _RAND_3512 = {1{`RANDOM}};
  T_38110_15_replay_if = _RAND_3512[0:0];
  _RAND_3513 = {2{`RANDOM}};
  T_38110_15_debug_wdata = _RAND_3513[63:0];
  _RAND_3514 = {1{`RANDOM}};
  T_38110_15_debug_events_fetch_seq = _RAND_3514[31:0];
  _RAND_3515 = {1{`RANDOM}};
  T_38110_16_valid = _RAND_3515[0:0];
  _RAND_3516 = {1{`RANDOM}};
  T_38110_16_iw_state = _RAND_3516[1:0];
  _RAND_3517 = {1{`RANDOM}};
  T_38110_16_uopc = _RAND_3517[8:0];
  _RAND_3518 = {1{`RANDOM}};
  T_38110_16_inst = _RAND_3518[31:0];
  _RAND_3519 = {2{`RANDOM}};
  T_38110_16_pc = _RAND_3519[39:0];
  _RAND_3520 = {1{`RANDOM}};
  T_38110_16_fu_code = _RAND_3520[7:0];
  _RAND_3521 = {1{`RANDOM}};
  T_38110_16_ctrl_br_type = _RAND_3521[3:0];
  _RAND_3522 = {1{`RANDOM}};
  T_38110_16_ctrl_op1_sel = _RAND_3522[1:0];
  _RAND_3523 = {1{`RANDOM}};
  T_38110_16_ctrl_op2_sel = _RAND_3523[2:0];
  _RAND_3524 = {1{`RANDOM}};
  T_38110_16_ctrl_imm_sel = _RAND_3524[2:0];
  _RAND_3525 = {1{`RANDOM}};
  T_38110_16_ctrl_op_fcn = _RAND_3525[3:0];
  _RAND_3526 = {1{`RANDOM}};
  T_38110_16_ctrl_fcn_dw = _RAND_3526[0:0];
  _RAND_3527 = {1{`RANDOM}};
  T_38110_16_ctrl_rf_wen = _RAND_3527[0:0];
  _RAND_3528 = {1{`RANDOM}};
  T_38110_16_ctrl_csr_cmd = _RAND_3528[2:0];
  _RAND_3529 = {1{`RANDOM}};
  T_38110_16_ctrl_is_load = _RAND_3529[0:0];
  _RAND_3530 = {1{`RANDOM}};
  T_38110_16_ctrl_is_sta = _RAND_3530[0:0];
  _RAND_3531 = {1{`RANDOM}};
  T_38110_16_ctrl_is_std = _RAND_3531[0:0];
  _RAND_3532 = {1{`RANDOM}};
  T_38110_16_wakeup_delay = _RAND_3532[1:0];
  _RAND_3533 = {1{`RANDOM}};
  T_38110_16_allocate_brtag = _RAND_3533[0:0];
  _RAND_3534 = {1{`RANDOM}};
  T_38110_16_is_br_or_jmp = _RAND_3534[0:0];
  _RAND_3535 = {1{`RANDOM}};
  T_38110_16_is_jump = _RAND_3535[0:0];
  _RAND_3536 = {1{`RANDOM}};
  T_38110_16_is_jal = _RAND_3536[0:0];
  _RAND_3537 = {1{`RANDOM}};
  T_38110_16_is_ret = _RAND_3537[0:0];
  _RAND_3538 = {1{`RANDOM}};
  T_38110_16_is_call = _RAND_3538[0:0];
  _RAND_3539 = {1{`RANDOM}};
  T_38110_16_br_mask = _RAND_3539[7:0];
  _RAND_3540 = {1{`RANDOM}};
  T_38110_16_br_tag = _RAND_3540[2:0];
  _RAND_3541 = {1{`RANDOM}};
  T_38110_16_br_prediction_bpd_predict_val = _RAND_3541[0:0];
  _RAND_3542 = {1{`RANDOM}};
  T_38110_16_br_prediction_bpd_predict_taken = _RAND_3542[0:0];
  _RAND_3543 = {1{`RANDOM}};
  T_38110_16_br_prediction_btb_hit = _RAND_3543[0:0];
  _RAND_3544 = {1{`RANDOM}};
  T_38110_16_br_prediction_btb_predicted = _RAND_3544[0:0];
  _RAND_3545 = {1{`RANDOM}};
  T_38110_16_br_prediction_is_br_or_jalr = _RAND_3545[0:0];
  _RAND_3546 = {1{`RANDOM}};
  T_38110_16_stat_brjmp_mispredicted = _RAND_3546[0:0];
  _RAND_3547 = {1{`RANDOM}};
  T_38110_16_stat_btb_made_pred = _RAND_3547[0:0];
  _RAND_3548 = {1{`RANDOM}};
  T_38110_16_stat_btb_mispredicted = _RAND_3548[0:0];
  _RAND_3549 = {1{`RANDOM}};
  T_38110_16_stat_bpd_made_pred = _RAND_3549[0:0];
  _RAND_3550 = {1{`RANDOM}};
  T_38110_16_stat_bpd_mispredicted = _RAND_3550[0:0];
  _RAND_3551 = {1{`RANDOM}};
  T_38110_16_fetch_pc_lob = _RAND_3551[2:0];
  _RAND_3552 = {1{`RANDOM}};
  T_38110_16_imm_packed = _RAND_3552[19:0];
  _RAND_3553 = {1{`RANDOM}};
  T_38110_16_csr_addr = _RAND_3553[11:0];
  _RAND_3554 = {1{`RANDOM}};
  T_38110_16_rob_idx = _RAND_3554[5:0];
  _RAND_3555 = {1{`RANDOM}};
  T_38110_16_ldq_idx = _RAND_3555[3:0];
  _RAND_3556 = {1{`RANDOM}};
  T_38110_16_stq_idx = _RAND_3556[3:0];
  _RAND_3557 = {1{`RANDOM}};
  T_38110_16_brob_idx = _RAND_3557[4:0];
  _RAND_3558 = {1{`RANDOM}};
  T_38110_16_pdst = _RAND_3558[6:0];
  _RAND_3559 = {1{`RANDOM}};
  T_38110_16_pop1 = _RAND_3559[6:0];
  _RAND_3560 = {1{`RANDOM}};
  T_38110_16_pop2 = _RAND_3560[6:0];
  _RAND_3561 = {1{`RANDOM}};
  T_38110_16_pop3 = _RAND_3561[6:0];
  _RAND_3562 = {1{`RANDOM}};
  T_38110_16_prs1_busy = _RAND_3562[0:0];
  _RAND_3563 = {1{`RANDOM}};
  T_38110_16_prs2_busy = _RAND_3563[0:0];
  _RAND_3564 = {1{`RANDOM}};
  T_38110_16_prs3_busy = _RAND_3564[0:0];
  _RAND_3565 = {1{`RANDOM}};
  T_38110_16_stale_pdst = _RAND_3565[6:0];
  _RAND_3566 = {1{`RANDOM}};
  T_38110_16_exception = _RAND_3566[0:0];
  _RAND_3567 = {2{`RANDOM}};
  T_38110_16_exc_cause = _RAND_3567[63:0];
  _RAND_3568 = {1{`RANDOM}};
  T_38110_16_bypassable = _RAND_3568[0:0];
  _RAND_3569 = {1{`RANDOM}};
  T_38110_16_mem_cmd = _RAND_3569[3:0];
  _RAND_3570 = {1{`RANDOM}};
  T_38110_16_mem_typ = _RAND_3570[2:0];
  _RAND_3571 = {1{`RANDOM}};
  T_38110_16_is_fence = _RAND_3571[0:0];
  _RAND_3572 = {1{`RANDOM}};
  T_38110_16_is_fencei = _RAND_3572[0:0];
  _RAND_3573 = {1{`RANDOM}};
  T_38110_16_is_store = _RAND_3573[0:0];
  _RAND_3574 = {1{`RANDOM}};
  T_38110_16_is_amo = _RAND_3574[0:0];
  _RAND_3575 = {1{`RANDOM}};
  T_38110_16_is_load = _RAND_3575[0:0];
  _RAND_3576 = {1{`RANDOM}};
  T_38110_16_is_unique = _RAND_3576[0:0];
  _RAND_3577 = {1{`RANDOM}};
  T_38110_16_flush_on_commit = _RAND_3577[0:0];
  _RAND_3578 = {1{`RANDOM}};
  T_38110_16_ldst = _RAND_3578[5:0];
  _RAND_3579 = {1{`RANDOM}};
  T_38110_16_lrs1 = _RAND_3579[5:0];
  _RAND_3580 = {1{`RANDOM}};
  T_38110_16_lrs2 = _RAND_3580[5:0];
  _RAND_3581 = {1{`RANDOM}};
  T_38110_16_lrs3 = _RAND_3581[5:0];
  _RAND_3582 = {1{`RANDOM}};
  T_38110_16_ldst_val = _RAND_3582[0:0];
  _RAND_3583 = {1{`RANDOM}};
  T_38110_16_dst_rtype = _RAND_3583[1:0];
  _RAND_3584 = {1{`RANDOM}};
  T_38110_16_lrs1_rtype = _RAND_3584[1:0];
  _RAND_3585 = {1{`RANDOM}};
  T_38110_16_lrs2_rtype = _RAND_3585[1:0];
  _RAND_3586 = {1{`RANDOM}};
  T_38110_16_frs3_en = _RAND_3586[0:0];
  _RAND_3587 = {1{`RANDOM}};
  T_38110_16_fp_val = _RAND_3587[0:0];
  _RAND_3588 = {1{`RANDOM}};
  T_38110_16_fp_single = _RAND_3588[0:0];
  _RAND_3589 = {1{`RANDOM}};
  T_38110_16_xcpt_if = _RAND_3589[0:0];
  _RAND_3590 = {1{`RANDOM}};
  T_38110_16_replay_if = _RAND_3590[0:0];
  _RAND_3591 = {2{`RANDOM}};
  T_38110_16_debug_wdata = _RAND_3591[63:0];
  _RAND_3592 = {1{`RANDOM}};
  T_38110_16_debug_events_fetch_seq = _RAND_3592[31:0];
  _RAND_3593 = {1{`RANDOM}};
  T_38110_17_valid = _RAND_3593[0:0];
  _RAND_3594 = {1{`RANDOM}};
  T_38110_17_iw_state = _RAND_3594[1:0];
  _RAND_3595 = {1{`RANDOM}};
  T_38110_17_uopc = _RAND_3595[8:0];
  _RAND_3596 = {1{`RANDOM}};
  T_38110_17_inst = _RAND_3596[31:0];
  _RAND_3597 = {2{`RANDOM}};
  T_38110_17_pc = _RAND_3597[39:0];
  _RAND_3598 = {1{`RANDOM}};
  T_38110_17_fu_code = _RAND_3598[7:0];
  _RAND_3599 = {1{`RANDOM}};
  T_38110_17_ctrl_br_type = _RAND_3599[3:0];
  _RAND_3600 = {1{`RANDOM}};
  T_38110_17_ctrl_op1_sel = _RAND_3600[1:0];
  _RAND_3601 = {1{`RANDOM}};
  T_38110_17_ctrl_op2_sel = _RAND_3601[2:0];
  _RAND_3602 = {1{`RANDOM}};
  T_38110_17_ctrl_imm_sel = _RAND_3602[2:0];
  _RAND_3603 = {1{`RANDOM}};
  T_38110_17_ctrl_op_fcn = _RAND_3603[3:0];
  _RAND_3604 = {1{`RANDOM}};
  T_38110_17_ctrl_fcn_dw = _RAND_3604[0:0];
  _RAND_3605 = {1{`RANDOM}};
  T_38110_17_ctrl_rf_wen = _RAND_3605[0:0];
  _RAND_3606 = {1{`RANDOM}};
  T_38110_17_ctrl_csr_cmd = _RAND_3606[2:0];
  _RAND_3607 = {1{`RANDOM}};
  T_38110_17_ctrl_is_load = _RAND_3607[0:0];
  _RAND_3608 = {1{`RANDOM}};
  T_38110_17_ctrl_is_sta = _RAND_3608[0:0];
  _RAND_3609 = {1{`RANDOM}};
  T_38110_17_ctrl_is_std = _RAND_3609[0:0];
  _RAND_3610 = {1{`RANDOM}};
  T_38110_17_wakeup_delay = _RAND_3610[1:0];
  _RAND_3611 = {1{`RANDOM}};
  T_38110_17_allocate_brtag = _RAND_3611[0:0];
  _RAND_3612 = {1{`RANDOM}};
  T_38110_17_is_br_or_jmp = _RAND_3612[0:0];
  _RAND_3613 = {1{`RANDOM}};
  T_38110_17_is_jump = _RAND_3613[0:0];
  _RAND_3614 = {1{`RANDOM}};
  T_38110_17_is_jal = _RAND_3614[0:0];
  _RAND_3615 = {1{`RANDOM}};
  T_38110_17_is_ret = _RAND_3615[0:0];
  _RAND_3616 = {1{`RANDOM}};
  T_38110_17_is_call = _RAND_3616[0:0];
  _RAND_3617 = {1{`RANDOM}};
  T_38110_17_br_mask = _RAND_3617[7:0];
  _RAND_3618 = {1{`RANDOM}};
  T_38110_17_br_tag = _RAND_3618[2:0];
  _RAND_3619 = {1{`RANDOM}};
  T_38110_17_br_prediction_bpd_predict_val = _RAND_3619[0:0];
  _RAND_3620 = {1{`RANDOM}};
  T_38110_17_br_prediction_bpd_predict_taken = _RAND_3620[0:0];
  _RAND_3621 = {1{`RANDOM}};
  T_38110_17_br_prediction_btb_hit = _RAND_3621[0:0];
  _RAND_3622 = {1{`RANDOM}};
  T_38110_17_br_prediction_btb_predicted = _RAND_3622[0:0];
  _RAND_3623 = {1{`RANDOM}};
  T_38110_17_br_prediction_is_br_or_jalr = _RAND_3623[0:0];
  _RAND_3624 = {1{`RANDOM}};
  T_38110_17_stat_brjmp_mispredicted = _RAND_3624[0:0];
  _RAND_3625 = {1{`RANDOM}};
  T_38110_17_stat_btb_made_pred = _RAND_3625[0:0];
  _RAND_3626 = {1{`RANDOM}};
  T_38110_17_stat_btb_mispredicted = _RAND_3626[0:0];
  _RAND_3627 = {1{`RANDOM}};
  T_38110_17_stat_bpd_made_pred = _RAND_3627[0:0];
  _RAND_3628 = {1{`RANDOM}};
  T_38110_17_stat_bpd_mispredicted = _RAND_3628[0:0];
  _RAND_3629 = {1{`RANDOM}};
  T_38110_17_fetch_pc_lob = _RAND_3629[2:0];
  _RAND_3630 = {1{`RANDOM}};
  T_38110_17_imm_packed = _RAND_3630[19:0];
  _RAND_3631 = {1{`RANDOM}};
  T_38110_17_csr_addr = _RAND_3631[11:0];
  _RAND_3632 = {1{`RANDOM}};
  T_38110_17_rob_idx = _RAND_3632[5:0];
  _RAND_3633 = {1{`RANDOM}};
  T_38110_17_ldq_idx = _RAND_3633[3:0];
  _RAND_3634 = {1{`RANDOM}};
  T_38110_17_stq_idx = _RAND_3634[3:0];
  _RAND_3635 = {1{`RANDOM}};
  T_38110_17_brob_idx = _RAND_3635[4:0];
  _RAND_3636 = {1{`RANDOM}};
  T_38110_17_pdst = _RAND_3636[6:0];
  _RAND_3637 = {1{`RANDOM}};
  T_38110_17_pop1 = _RAND_3637[6:0];
  _RAND_3638 = {1{`RANDOM}};
  T_38110_17_pop2 = _RAND_3638[6:0];
  _RAND_3639 = {1{`RANDOM}};
  T_38110_17_pop3 = _RAND_3639[6:0];
  _RAND_3640 = {1{`RANDOM}};
  T_38110_17_prs1_busy = _RAND_3640[0:0];
  _RAND_3641 = {1{`RANDOM}};
  T_38110_17_prs2_busy = _RAND_3641[0:0];
  _RAND_3642 = {1{`RANDOM}};
  T_38110_17_prs3_busy = _RAND_3642[0:0];
  _RAND_3643 = {1{`RANDOM}};
  T_38110_17_stale_pdst = _RAND_3643[6:0];
  _RAND_3644 = {1{`RANDOM}};
  T_38110_17_exception = _RAND_3644[0:0];
  _RAND_3645 = {2{`RANDOM}};
  T_38110_17_exc_cause = _RAND_3645[63:0];
  _RAND_3646 = {1{`RANDOM}};
  T_38110_17_bypassable = _RAND_3646[0:0];
  _RAND_3647 = {1{`RANDOM}};
  T_38110_17_mem_cmd = _RAND_3647[3:0];
  _RAND_3648 = {1{`RANDOM}};
  T_38110_17_mem_typ = _RAND_3648[2:0];
  _RAND_3649 = {1{`RANDOM}};
  T_38110_17_is_fence = _RAND_3649[0:0];
  _RAND_3650 = {1{`RANDOM}};
  T_38110_17_is_fencei = _RAND_3650[0:0];
  _RAND_3651 = {1{`RANDOM}};
  T_38110_17_is_store = _RAND_3651[0:0];
  _RAND_3652 = {1{`RANDOM}};
  T_38110_17_is_amo = _RAND_3652[0:0];
  _RAND_3653 = {1{`RANDOM}};
  T_38110_17_is_load = _RAND_3653[0:0];
  _RAND_3654 = {1{`RANDOM}};
  T_38110_17_is_unique = _RAND_3654[0:0];
  _RAND_3655 = {1{`RANDOM}};
  T_38110_17_flush_on_commit = _RAND_3655[0:0];
  _RAND_3656 = {1{`RANDOM}};
  T_38110_17_ldst = _RAND_3656[5:0];
  _RAND_3657 = {1{`RANDOM}};
  T_38110_17_lrs1 = _RAND_3657[5:0];
  _RAND_3658 = {1{`RANDOM}};
  T_38110_17_lrs2 = _RAND_3658[5:0];
  _RAND_3659 = {1{`RANDOM}};
  T_38110_17_lrs3 = _RAND_3659[5:0];
  _RAND_3660 = {1{`RANDOM}};
  T_38110_17_ldst_val = _RAND_3660[0:0];
  _RAND_3661 = {1{`RANDOM}};
  T_38110_17_dst_rtype = _RAND_3661[1:0];
  _RAND_3662 = {1{`RANDOM}};
  T_38110_17_lrs1_rtype = _RAND_3662[1:0];
  _RAND_3663 = {1{`RANDOM}};
  T_38110_17_lrs2_rtype = _RAND_3663[1:0];
  _RAND_3664 = {1{`RANDOM}};
  T_38110_17_frs3_en = _RAND_3664[0:0];
  _RAND_3665 = {1{`RANDOM}};
  T_38110_17_fp_val = _RAND_3665[0:0];
  _RAND_3666 = {1{`RANDOM}};
  T_38110_17_fp_single = _RAND_3666[0:0];
  _RAND_3667 = {1{`RANDOM}};
  T_38110_17_xcpt_if = _RAND_3667[0:0];
  _RAND_3668 = {1{`RANDOM}};
  T_38110_17_replay_if = _RAND_3668[0:0];
  _RAND_3669 = {2{`RANDOM}};
  T_38110_17_debug_wdata = _RAND_3669[63:0];
  _RAND_3670 = {1{`RANDOM}};
  T_38110_17_debug_events_fetch_seq = _RAND_3670[31:0];
  _RAND_3671 = {1{`RANDOM}};
  T_38110_18_valid = _RAND_3671[0:0];
  _RAND_3672 = {1{`RANDOM}};
  T_38110_18_iw_state = _RAND_3672[1:0];
  _RAND_3673 = {1{`RANDOM}};
  T_38110_18_uopc = _RAND_3673[8:0];
  _RAND_3674 = {1{`RANDOM}};
  T_38110_18_inst = _RAND_3674[31:0];
  _RAND_3675 = {2{`RANDOM}};
  T_38110_18_pc = _RAND_3675[39:0];
  _RAND_3676 = {1{`RANDOM}};
  T_38110_18_fu_code = _RAND_3676[7:0];
  _RAND_3677 = {1{`RANDOM}};
  T_38110_18_ctrl_br_type = _RAND_3677[3:0];
  _RAND_3678 = {1{`RANDOM}};
  T_38110_18_ctrl_op1_sel = _RAND_3678[1:0];
  _RAND_3679 = {1{`RANDOM}};
  T_38110_18_ctrl_op2_sel = _RAND_3679[2:0];
  _RAND_3680 = {1{`RANDOM}};
  T_38110_18_ctrl_imm_sel = _RAND_3680[2:0];
  _RAND_3681 = {1{`RANDOM}};
  T_38110_18_ctrl_op_fcn = _RAND_3681[3:0];
  _RAND_3682 = {1{`RANDOM}};
  T_38110_18_ctrl_fcn_dw = _RAND_3682[0:0];
  _RAND_3683 = {1{`RANDOM}};
  T_38110_18_ctrl_rf_wen = _RAND_3683[0:0];
  _RAND_3684 = {1{`RANDOM}};
  T_38110_18_ctrl_csr_cmd = _RAND_3684[2:0];
  _RAND_3685 = {1{`RANDOM}};
  T_38110_18_ctrl_is_load = _RAND_3685[0:0];
  _RAND_3686 = {1{`RANDOM}};
  T_38110_18_ctrl_is_sta = _RAND_3686[0:0];
  _RAND_3687 = {1{`RANDOM}};
  T_38110_18_ctrl_is_std = _RAND_3687[0:0];
  _RAND_3688 = {1{`RANDOM}};
  T_38110_18_wakeup_delay = _RAND_3688[1:0];
  _RAND_3689 = {1{`RANDOM}};
  T_38110_18_allocate_brtag = _RAND_3689[0:0];
  _RAND_3690 = {1{`RANDOM}};
  T_38110_18_is_br_or_jmp = _RAND_3690[0:0];
  _RAND_3691 = {1{`RANDOM}};
  T_38110_18_is_jump = _RAND_3691[0:0];
  _RAND_3692 = {1{`RANDOM}};
  T_38110_18_is_jal = _RAND_3692[0:0];
  _RAND_3693 = {1{`RANDOM}};
  T_38110_18_is_ret = _RAND_3693[0:0];
  _RAND_3694 = {1{`RANDOM}};
  T_38110_18_is_call = _RAND_3694[0:0];
  _RAND_3695 = {1{`RANDOM}};
  T_38110_18_br_mask = _RAND_3695[7:0];
  _RAND_3696 = {1{`RANDOM}};
  T_38110_18_br_tag = _RAND_3696[2:0];
  _RAND_3697 = {1{`RANDOM}};
  T_38110_18_br_prediction_bpd_predict_val = _RAND_3697[0:0];
  _RAND_3698 = {1{`RANDOM}};
  T_38110_18_br_prediction_bpd_predict_taken = _RAND_3698[0:0];
  _RAND_3699 = {1{`RANDOM}};
  T_38110_18_br_prediction_btb_hit = _RAND_3699[0:0];
  _RAND_3700 = {1{`RANDOM}};
  T_38110_18_br_prediction_btb_predicted = _RAND_3700[0:0];
  _RAND_3701 = {1{`RANDOM}};
  T_38110_18_br_prediction_is_br_or_jalr = _RAND_3701[0:0];
  _RAND_3702 = {1{`RANDOM}};
  T_38110_18_stat_brjmp_mispredicted = _RAND_3702[0:0];
  _RAND_3703 = {1{`RANDOM}};
  T_38110_18_stat_btb_made_pred = _RAND_3703[0:0];
  _RAND_3704 = {1{`RANDOM}};
  T_38110_18_stat_btb_mispredicted = _RAND_3704[0:0];
  _RAND_3705 = {1{`RANDOM}};
  T_38110_18_stat_bpd_made_pred = _RAND_3705[0:0];
  _RAND_3706 = {1{`RANDOM}};
  T_38110_18_stat_bpd_mispredicted = _RAND_3706[0:0];
  _RAND_3707 = {1{`RANDOM}};
  T_38110_18_fetch_pc_lob = _RAND_3707[2:0];
  _RAND_3708 = {1{`RANDOM}};
  T_38110_18_imm_packed = _RAND_3708[19:0];
  _RAND_3709 = {1{`RANDOM}};
  T_38110_18_csr_addr = _RAND_3709[11:0];
  _RAND_3710 = {1{`RANDOM}};
  T_38110_18_rob_idx = _RAND_3710[5:0];
  _RAND_3711 = {1{`RANDOM}};
  T_38110_18_ldq_idx = _RAND_3711[3:0];
  _RAND_3712 = {1{`RANDOM}};
  T_38110_18_stq_idx = _RAND_3712[3:0];
  _RAND_3713 = {1{`RANDOM}};
  T_38110_18_brob_idx = _RAND_3713[4:0];
  _RAND_3714 = {1{`RANDOM}};
  T_38110_18_pdst = _RAND_3714[6:0];
  _RAND_3715 = {1{`RANDOM}};
  T_38110_18_pop1 = _RAND_3715[6:0];
  _RAND_3716 = {1{`RANDOM}};
  T_38110_18_pop2 = _RAND_3716[6:0];
  _RAND_3717 = {1{`RANDOM}};
  T_38110_18_pop3 = _RAND_3717[6:0];
  _RAND_3718 = {1{`RANDOM}};
  T_38110_18_prs1_busy = _RAND_3718[0:0];
  _RAND_3719 = {1{`RANDOM}};
  T_38110_18_prs2_busy = _RAND_3719[0:0];
  _RAND_3720 = {1{`RANDOM}};
  T_38110_18_prs3_busy = _RAND_3720[0:0];
  _RAND_3721 = {1{`RANDOM}};
  T_38110_18_stale_pdst = _RAND_3721[6:0];
  _RAND_3722 = {1{`RANDOM}};
  T_38110_18_exception = _RAND_3722[0:0];
  _RAND_3723 = {2{`RANDOM}};
  T_38110_18_exc_cause = _RAND_3723[63:0];
  _RAND_3724 = {1{`RANDOM}};
  T_38110_18_bypassable = _RAND_3724[0:0];
  _RAND_3725 = {1{`RANDOM}};
  T_38110_18_mem_cmd = _RAND_3725[3:0];
  _RAND_3726 = {1{`RANDOM}};
  T_38110_18_mem_typ = _RAND_3726[2:0];
  _RAND_3727 = {1{`RANDOM}};
  T_38110_18_is_fence = _RAND_3727[0:0];
  _RAND_3728 = {1{`RANDOM}};
  T_38110_18_is_fencei = _RAND_3728[0:0];
  _RAND_3729 = {1{`RANDOM}};
  T_38110_18_is_store = _RAND_3729[0:0];
  _RAND_3730 = {1{`RANDOM}};
  T_38110_18_is_amo = _RAND_3730[0:0];
  _RAND_3731 = {1{`RANDOM}};
  T_38110_18_is_load = _RAND_3731[0:0];
  _RAND_3732 = {1{`RANDOM}};
  T_38110_18_is_unique = _RAND_3732[0:0];
  _RAND_3733 = {1{`RANDOM}};
  T_38110_18_flush_on_commit = _RAND_3733[0:0];
  _RAND_3734 = {1{`RANDOM}};
  T_38110_18_ldst = _RAND_3734[5:0];
  _RAND_3735 = {1{`RANDOM}};
  T_38110_18_lrs1 = _RAND_3735[5:0];
  _RAND_3736 = {1{`RANDOM}};
  T_38110_18_lrs2 = _RAND_3736[5:0];
  _RAND_3737 = {1{`RANDOM}};
  T_38110_18_lrs3 = _RAND_3737[5:0];
  _RAND_3738 = {1{`RANDOM}};
  T_38110_18_ldst_val = _RAND_3738[0:0];
  _RAND_3739 = {1{`RANDOM}};
  T_38110_18_dst_rtype = _RAND_3739[1:0];
  _RAND_3740 = {1{`RANDOM}};
  T_38110_18_lrs1_rtype = _RAND_3740[1:0];
  _RAND_3741 = {1{`RANDOM}};
  T_38110_18_lrs2_rtype = _RAND_3741[1:0];
  _RAND_3742 = {1{`RANDOM}};
  T_38110_18_frs3_en = _RAND_3742[0:0];
  _RAND_3743 = {1{`RANDOM}};
  T_38110_18_fp_val = _RAND_3743[0:0];
  _RAND_3744 = {1{`RANDOM}};
  T_38110_18_fp_single = _RAND_3744[0:0];
  _RAND_3745 = {1{`RANDOM}};
  T_38110_18_xcpt_if = _RAND_3745[0:0];
  _RAND_3746 = {1{`RANDOM}};
  T_38110_18_replay_if = _RAND_3746[0:0];
  _RAND_3747 = {2{`RANDOM}};
  T_38110_18_debug_wdata = _RAND_3747[63:0];
  _RAND_3748 = {1{`RANDOM}};
  T_38110_18_debug_events_fetch_seq = _RAND_3748[31:0];
  _RAND_3749 = {1{`RANDOM}};
  T_38110_19_valid = _RAND_3749[0:0];
  _RAND_3750 = {1{`RANDOM}};
  T_38110_19_iw_state = _RAND_3750[1:0];
  _RAND_3751 = {1{`RANDOM}};
  T_38110_19_uopc = _RAND_3751[8:0];
  _RAND_3752 = {1{`RANDOM}};
  T_38110_19_inst = _RAND_3752[31:0];
  _RAND_3753 = {2{`RANDOM}};
  T_38110_19_pc = _RAND_3753[39:0];
  _RAND_3754 = {1{`RANDOM}};
  T_38110_19_fu_code = _RAND_3754[7:0];
  _RAND_3755 = {1{`RANDOM}};
  T_38110_19_ctrl_br_type = _RAND_3755[3:0];
  _RAND_3756 = {1{`RANDOM}};
  T_38110_19_ctrl_op1_sel = _RAND_3756[1:0];
  _RAND_3757 = {1{`RANDOM}};
  T_38110_19_ctrl_op2_sel = _RAND_3757[2:0];
  _RAND_3758 = {1{`RANDOM}};
  T_38110_19_ctrl_imm_sel = _RAND_3758[2:0];
  _RAND_3759 = {1{`RANDOM}};
  T_38110_19_ctrl_op_fcn = _RAND_3759[3:0];
  _RAND_3760 = {1{`RANDOM}};
  T_38110_19_ctrl_fcn_dw = _RAND_3760[0:0];
  _RAND_3761 = {1{`RANDOM}};
  T_38110_19_ctrl_rf_wen = _RAND_3761[0:0];
  _RAND_3762 = {1{`RANDOM}};
  T_38110_19_ctrl_csr_cmd = _RAND_3762[2:0];
  _RAND_3763 = {1{`RANDOM}};
  T_38110_19_ctrl_is_load = _RAND_3763[0:0];
  _RAND_3764 = {1{`RANDOM}};
  T_38110_19_ctrl_is_sta = _RAND_3764[0:0];
  _RAND_3765 = {1{`RANDOM}};
  T_38110_19_ctrl_is_std = _RAND_3765[0:0];
  _RAND_3766 = {1{`RANDOM}};
  T_38110_19_wakeup_delay = _RAND_3766[1:0];
  _RAND_3767 = {1{`RANDOM}};
  T_38110_19_allocate_brtag = _RAND_3767[0:0];
  _RAND_3768 = {1{`RANDOM}};
  T_38110_19_is_br_or_jmp = _RAND_3768[0:0];
  _RAND_3769 = {1{`RANDOM}};
  T_38110_19_is_jump = _RAND_3769[0:0];
  _RAND_3770 = {1{`RANDOM}};
  T_38110_19_is_jal = _RAND_3770[0:0];
  _RAND_3771 = {1{`RANDOM}};
  T_38110_19_is_ret = _RAND_3771[0:0];
  _RAND_3772 = {1{`RANDOM}};
  T_38110_19_is_call = _RAND_3772[0:0];
  _RAND_3773 = {1{`RANDOM}};
  T_38110_19_br_mask = _RAND_3773[7:0];
  _RAND_3774 = {1{`RANDOM}};
  T_38110_19_br_tag = _RAND_3774[2:0];
  _RAND_3775 = {1{`RANDOM}};
  T_38110_19_br_prediction_bpd_predict_val = _RAND_3775[0:0];
  _RAND_3776 = {1{`RANDOM}};
  T_38110_19_br_prediction_bpd_predict_taken = _RAND_3776[0:0];
  _RAND_3777 = {1{`RANDOM}};
  T_38110_19_br_prediction_btb_hit = _RAND_3777[0:0];
  _RAND_3778 = {1{`RANDOM}};
  T_38110_19_br_prediction_btb_predicted = _RAND_3778[0:0];
  _RAND_3779 = {1{`RANDOM}};
  T_38110_19_br_prediction_is_br_or_jalr = _RAND_3779[0:0];
  _RAND_3780 = {1{`RANDOM}};
  T_38110_19_stat_brjmp_mispredicted = _RAND_3780[0:0];
  _RAND_3781 = {1{`RANDOM}};
  T_38110_19_stat_btb_made_pred = _RAND_3781[0:0];
  _RAND_3782 = {1{`RANDOM}};
  T_38110_19_stat_btb_mispredicted = _RAND_3782[0:0];
  _RAND_3783 = {1{`RANDOM}};
  T_38110_19_stat_bpd_made_pred = _RAND_3783[0:0];
  _RAND_3784 = {1{`RANDOM}};
  T_38110_19_stat_bpd_mispredicted = _RAND_3784[0:0];
  _RAND_3785 = {1{`RANDOM}};
  T_38110_19_fetch_pc_lob = _RAND_3785[2:0];
  _RAND_3786 = {1{`RANDOM}};
  T_38110_19_imm_packed = _RAND_3786[19:0];
  _RAND_3787 = {1{`RANDOM}};
  T_38110_19_csr_addr = _RAND_3787[11:0];
  _RAND_3788 = {1{`RANDOM}};
  T_38110_19_rob_idx = _RAND_3788[5:0];
  _RAND_3789 = {1{`RANDOM}};
  T_38110_19_ldq_idx = _RAND_3789[3:0];
  _RAND_3790 = {1{`RANDOM}};
  T_38110_19_stq_idx = _RAND_3790[3:0];
  _RAND_3791 = {1{`RANDOM}};
  T_38110_19_brob_idx = _RAND_3791[4:0];
  _RAND_3792 = {1{`RANDOM}};
  T_38110_19_pdst = _RAND_3792[6:0];
  _RAND_3793 = {1{`RANDOM}};
  T_38110_19_pop1 = _RAND_3793[6:0];
  _RAND_3794 = {1{`RANDOM}};
  T_38110_19_pop2 = _RAND_3794[6:0];
  _RAND_3795 = {1{`RANDOM}};
  T_38110_19_pop3 = _RAND_3795[6:0];
  _RAND_3796 = {1{`RANDOM}};
  T_38110_19_prs1_busy = _RAND_3796[0:0];
  _RAND_3797 = {1{`RANDOM}};
  T_38110_19_prs2_busy = _RAND_3797[0:0];
  _RAND_3798 = {1{`RANDOM}};
  T_38110_19_prs3_busy = _RAND_3798[0:0];
  _RAND_3799 = {1{`RANDOM}};
  T_38110_19_stale_pdst = _RAND_3799[6:0];
  _RAND_3800 = {1{`RANDOM}};
  T_38110_19_exception = _RAND_3800[0:0];
  _RAND_3801 = {2{`RANDOM}};
  T_38110_19_exc_cause = _RAND_3801[63:0];
  _RAND_3802 = {1{`RANDOM}};
  T_38110_19_bypassable = _RAND_3802[0:0];
  _RAND_3803 = {1{`RANDOM}};
  T_38110_19_mem_cmd = _RAND_3803[3:0];
  _RAND_3804 = {1{`RANDOM}};
  T_38110_19_mem_typ = _RAND_3804[2:0];
  _RAND_3805 = {1{`RANDOM}};
  T_38110_19_is_fence = _RAND_3805[0:0];
  _RAND_3806 = {1{`RANDOM}};
  T_38110_19_is_fencei = _RAND_3806[0:0];
  _RAND_3807 = {1{`RANDOM}};
  T_38110_19_is_store = _RAND_3807[0:0];
  _RAND_3808 = {1{`RANDOM}};
  T_38110_19_is_amo = _RAND_3808[0:0];
  _RAND_3809 = {1{`RANDOM}};
  T_38110_19_is_load = _RAND_3809[0:0];
  _RAND_3810 = {1{`RANDOM}};
  T_38110_19_is_unique = _RAND_3810[0:0];
  _RAND_3811 = {1{`RANDOM}};
  T_38110_19_flush_on_commit = _RAND_3811[0:0];
  _RAND_3812 = {1{`RANDOM}};
  T_38110_19_ldst = _RAND_3812[5:0];
  _RAND_3813 = {1{`RANDOM}};
  T_38110_19_lrs1 = _RAND_3813[5:0];
  _RAND_3814 = {1{`RANDOM}};
  T_38110_19_lrs2 = _RAND_3814[5:0];
  _RAND_3815 = {1{`RANDOM}};
  T_38110_19_lrs3 = _RAND_3815[5:0];
  _RAND_3816 = {1{`RANDOM}};
  T_38110_19_ldst_val = _RAND_3816[0:0];
  _RAND_3817 = {1{`RANDOM}};
  T_38110_19_dst_rtype = _RAND_3817[1:0];
  _RAND_3818 = {1{`RANDOM}};
  T_38110_19_lrs1_rtype = _RAND_3818[1:0];
  _RAND_3819 = {1{`RANDOM}};
  T_38110_19_lrs2_rtype = _RAND_3819[1:0];
  _RAND_3820 = {1{`RANDOM}};
  T_38110_19_frs3_en = _RAND_3820[0:0];
  _RAND_3821 = {1{`RANDOM}};
  T_38110_19_fp_val = _RAND_3821[0:0];
  _RAND_3822 = {1{`RANDOM}};
  T_38110_19_fp_single = _RAND_3822[0:0];
  _RAND_3823 = {1{`RANDOM}};
  T_38110_19_xcpt_if = _RAND_3823[0:0];
  _RAND_3824 = {1{`RANDOM}};
  T_38110_19_replay_if = _RAND_3824[0:0];
  _RAND_3825 = {2{`RANDOM}};
  T_38110_19_debug_wdata = _RAND_3825[63:0];
  _RAND_3826 = {1{`RANDOM}};
  T_38110_19_debug_events_fetch_seq = _RAND_3826[31:0];
  _RAND_3827 = {1{`RANDOM}};
  T_38110_20_valid = _RAND_3827[0:0];
  _RAND_3828 = {1{`RANDOM}};
  T_38110_20_iw_state = _RAND_3828[1:0];
  _RAND_3829 = {1{`RANDOM}};
  T_38110_20_uopc = _RAND_3829[8:0];
  _RAND_3830 = {1{`RANDOM}};
  T_38110_20_inst = _RAND_3830[31:0];
  _RAND_3831 = {2{`RANDOM}};
  T_38110_20_pc = _RAND_3831[39:0];
  _RAND_3832 = {1{`RANDOM}};
  T_38110_20_fu_code = _RAND_3832[7:0];
  _RAND_3833 = {1{`RANDOM}};
  T_38110_20_ctrl_br_type = _RAND_3833[3:0];
  _RAND_3834 = {1{`RANDOM}};
  T_38110_20_ctrl_op1_sel = _RAND_3834[1:0];
  _RAND_3835 = {1{`RANDOM}};
  T_38110_20_ctrl_op2_sel = _RAND_3835[2:0];
  _RAND_3836 = {1{`RANDOM}};
  T_38110_20_ctrl_imm_sel = _RAND_3836[2:0];
  _RAND_3837 = {1{`RANDOM}};
  T_38110_20_ctrl_op_fcn = _RAND_3837[3:0];
  _RAND_3838 = {1{`RANDOM}};
  T_38110_20_ctrl_fcn_dw = _RAND_3838[0:0];
  _RAND_3839 = {1{`RANDOM}};
  T_38110_20_ctrl_rf_wen = _RAND_3839[0:0];
  _RAND_3840 = {1{`RANDOM}};
  T_38110_20_ctrl_csr_cmd = _RAND_3840[2:0];
  _RAND_3841 = {1{`RANDOM}};
  T_38110_20_ctrl_is_load = _RAND_3841[0:0];
  _RAND_3842 = {1{`RANDOM}};
  T_38110_20_ctrl_is_sta = _RAND_3842[0:0];
  _RAND_3843 = {1{`RANDOM}};
  T_38110_20_ctrl_is_std = _RAND_3843[0:0];
  _RAND_3844 = {1{`RANDOM}};
  T_38110_20_wakeup_delay = _RAND_3844[1:0];
  _RAND_3845 = {1{`RANDOM}};
  T_38110_20_allocate_brtag = _RAND_3845[0:0];
  _RAND_3846 = {1{`RANDOM}};
  T_38110_20_is_br_or_jmp = _RAND_3846[0:0];
  _RAND_3847 = {1{`RANDOM}};
  T_38110_20_is_jump = _RAND_3847[0:0];
  _RAND_3848 = {1{`RANDOM}};
  T_38110_20_is_jal = _RAND_3848[0:0];
  _RAND_3849 = {1{`RANDOM}};
  T_38110_20_is_ret = _RAND_3849[0:0];
  _RAND_3850 = {1{`RANDOM}};
  T_38110_20_is_call = _RAND_3850[0:0];
  _RAND_3851 = {1{`RANDOM}};
  T_38110_20_br_mask = _RAND_3851[7:0];
  _RAND_3852 = {1{`RANDOM}};
  T_38110_20_br_tag = _RAND_3852[2:0];
  _RAND_3853 = {1{`RANDOM}};
  T_38110_20_br_prediction_bpd_predict_val = _RAND_3853[0:0];
  _RAND_3854 = {1{`RANDOM}};
  T_38110_20_br_prediction_bpd_predict_taken = _RAND_3854[0:0];
  _RAND_3855 = {1{`RANDOM}};
  T_38110_20_br_prediction_btb_hit = _RAND_3855[0:0];
  _RAND_3856 = {1{`RANDOM}};
  T_38110_20_br_prediction_btb_predicted = _RAND_3856[0:0];
  _RAND_3857 = {1{`RANDOM}};
  T_38110_20_br_prediction_is_br_or_jalr = _RAND_3857[0:0];
  _RAND_3858 = {1{`RANDOM}};
  T_38110_20_stat_brjmp_mispredicted = _RAND_3858[0:0];
  _RAND_3859 = {1{`RANDOM}};
  T_38110_20_stat_btb_made_pred = _RAND_3859[0:0];
  _RAND_3860 = {1{`RANDOM}};
  T_38110_20_stat_btb_mispredicted = _RAND_3860[0:0];
  _RAND_3861 = {1{`RANDOM}};
  T_38110_20_stat_bpd_made_pred = _RAND_3861[0:0];
  _RAND_3862 = {1{`RANDOM}};
  T_38110_20_stat_bpd_mispredicted = _RAND_3862[0:0];
  _RAND_3863 = {1{`RANDOM}};
  T_38110_20_fetch_pc_lob = _RAND_3863[2:0];
  _RAND_3864 = {1{`RANDOM}};
  T_38110_20_imm_packed = _RAND_3864[19:0];
  _RAND_3865 = {1{`RANDOM}};
  T_38110_20_csr_addr = _RAND_3865[11:0];
  _RAND_3866 = {1{`RANDOM}};
  T_38110_20_rob_idx = _RAND_3866[5:0];
  _RAND_3867 = {1{`RANDOM}};
  T_38110_20_ldq_idx = _RAND_3867[3:0];
  _RAND_3868 = {1{`RANDOM}};
  T_38110_20_stq_idx = _RAND_3868[3:0];
  _RAND_3869 = {1{`RANDOM}};
  T_38110_20_brob_idx = _RAND_3869[4:0];
  _RAND_3870 = {1{`RANDOM}};
  T_38110_20_pdst = _RAND_3870[6:0];
  _RAND_3871 = {1{`RANDOM}};
  T_38110_20_pop1 = _RAND_3871[6:0];
  _RAND_3872 = {1{`RANDOM}};
  T_38110_20_pop2 = _RAND_3872[6:0];
  _RAND_3873 = {1{`RANDOM}};
  T_38110_20_pop3 = _RAND_3873[6:0];
  _RAND_3874 = {1{`RANDOM}};
  T_38110_20_prs1_busy = _RAND_3874[0:0];
  _RAND_3875 = {1{`RANDOM}};
  T_38110_20_prs2_busy = _RAND_3875[0:0];
  _RAND_3876 = {1{`RANDOM}};
  T_38110_20_prs3_busy = _RAND_3876[0:0];
  _RAND_3877 = {1{`RANDOM}};
  T_38110_20_stale_pdst = _RAND_3877[6:0];
  _RAND_3878 = {1{`RANDOM}};
  T_38110_20_exception = _RAND_3878[0:0];
  _RAND_3879 = {2{`RANDOM}};
  T_38110_20_exc_cause = _RAND_3879[63:0];
  _RAND_3880 = {1{`RANDOM}};
  T_38110_20_bypassable = _RAND_3880[0:0];
  _RAND_3881 = {1{`RANDOM}};
  T_38110_20_mem_cmd = _RAND_3881[3:0];
  _RAND_3882 = {1{`RANDOM}};
  T_38110_20_mem_typ = _RAND_3882[2:0];
  _RAND_3883 = {1{`RANDOM}};
  T_38110_20_is_fence = _RAND_3883[0:0];
  _RAND_3884 = {1{`RANDOM}};
  T_38110_20_is_fencei = _RAND_3884[0:0];
  _RAND_3885 = {1{`RANDOM}};
  T_38110_20_is_store = _RAND_3885[0:0];
  _RAND_3886 = {1{`RANDOM}};
  T_38110_20_is_amo = _RAND_3886[0:0];
  _RAND_3887 = {1{`RANDOM}};
  T_38110_20_is_load = _RAND_3887[0:0];
  _RAND_3888 = {1{`RANDOM}};
  T_38110_20_is_unique = _RAND_3888[0:0];
  _RAND_3889 = {1{`RANDOM}};
  T_38110_20_flush_on_commit = _RAND_3889[0:0];
  _RAND_3890 = {1{`RANDOM}};
  T_38110_20_ldst = _RAND_3890[5:0];
  _RAND_3891 = {1{`RANDOM}};
  T_38110_20_lrs1 = _RAND_3891[5:0];
  _RAND_3892 = {1{`RANDOM}};
  T_38110_20_lrs2 = _RAND_3892[5:0];
  _RAND_3893 = {1{`RANDOM}};
  T_38110_20_lrs3 = _RAND_3893[5:0];
  _RAND_3894 = {1{`RANDOM}};
  T_38110_20_ldst_val = _RAND_3894[0:0];
  _RAND_3895 = {1{`RANDOM}};
  T_38110_20_dst_rtype = _RAND_3895[1:0];
  _RAND_3896 = {1{`RANDOM}};
  T_38110_20_lrs1_rtype = _RAND_3896[1:0];
  _RAND_3897 = {1{`RANDOM}};
  T_38110_20_lrs2_rtype = _RAND_3897[1:0];
  _RAND_3898 = {1{`RANDOM}};
  T_38110_20_frs3_en = _RAND_3898[0:0];
  _RAND_3899 = {1{`RANDOM}};
  T_38110_20_fp_val = _RAND_3899[0:0];
  _RAND_3900 = {1{`RANDOM}};
  T_38110_20_fp_single = _RAND_3900[0:0];
  _RAND_3901 = {1{`RANDOM}};
  T_38110_20_xcpt_if = _RAND_3901[0:0];
  _RAND_3902 = {1{`RANDOM}};
  T_38110_20_replay_if = _RAND_3902[0:0];
  _RAND_3903 = {2{`RANDOM}};
  T_38110_20_debug_wdata = _RAND_3903[63:0];
  _RAND_3904 = {1{`RANDOM}};
  T_38110_20_debug_events_fetch_seq = _RAND_3904[31:0];
  _RAND_3905 = {1{`RANDOM}};
  T_38110_21_valid = _RAND_3905[0:0];
  _RAND_3906 = {1{`RANDOM}};
  T_38110_21_iw_state = _RAND_3906[1:0];
  _RAND_3907 = {1{`RANDOM}};
  T_38110_21_uopc = _RAND_3907[8:0];
  _RAND_3908 = {1{`RANDOM}};
  T_38110_21_inst = _RAND_3908[31:0];
  _RAND_3909 = {2{`RANDOM}};
  T_38110_21_pc = _RAND_3909[39:0];
  _RAND_3910 = {1{`RANDOM}};
  T_38110_21_fu_code = _RAND_3910[7:0];
  _RAND_3911 = {1{`RANDOM}};
  T_38110_21_ctrl_br_type = _RAND_3911[3:0];
  _RAND_3912 = {1{`RANDOM}};
  T_38110_21_ctrl_op1_sel = _RAND_3912[1:0];
  _RAND_3913 = {1{`RANDOM}};
  T_38110_21_ctrl_op2_sel = _RAND_3913[2:0];
  _RAND_3914 = {1{`RANDOM}};
  T_38110_21_ctrl_imm_sel = _RAND_3914[2:0];
  _RAND_3915 = {1{`RANDOM}};
  T_38110_21_ctrl_op_fcn = _RAND_3915[3:0];
  _RAND_3916 = {1{`RANDOM}};
  T_38110_21_ctrl_fcn_dw = _RAND_3916[0:0];
  _RAND_3917 = {1{`RANDOM}};
  T_38110_21_ctrl_rf_wen = _RAND_3917[0:0];
  _RAND_3918 = {1{`RANDOM}};
  T_38110_21_ctrl_csr_cmd = _RAND_3918[2:0];
  _RAND_3919 = {1{`RANDOM}};
  T_38110_21_ctrl_is_load = _RAND_3919[0:0];
  _RAND_3920 = {1{`RANDOM}};
  T_38110_21_ctrl_is_sta = _RAND_3920[0:0];
  _RAND_3921 = {1{`RANDOM}};
  T_38110_21_ctrl_is_std = _RAND_3921[0:0];
  _RAND_3922 = {1{`RANDOM}};
  T_38110_21_wakeup_delay = _RAND_3922[1:0];
  _RAND_3923 = {1{`RANDOM}};
  T_38110_21_allocate_brtag = _RAND_3923[0:0];
  _RAND_3924 = {1{`RANDOM}};
  T_38110_21_is_br_or_jmp = _RAND_3924[0:0];
  _RAND_3925 = {1{`RANDOM}};
  T_38110_21_is_jump = _RAND_3925[0:0];
  _RAND_3926 = {1{`RANDOM}};
  T_38110_21_is_jal = _RAND_3926[0:0];
  _RAND_3927 = {1{`RANDOM}};
  T_38110_21_is_ret = _RAND_3927[0:0];
  _RAND_3928 = {1{`RANDOM}};
  T_38110_21_is_call = _RAND_3928[0:0];
  _RAND_3929 = {1{`RANDOM}};
  T_38110_21_br_mask = _RAND_3929[7:0];
  _RAND_3930 = {1{`RANDOM}};
  T_38110_21_br_tag = _RAND_3930[2:0];
  _RAND_3931 = {1{`RANDOM}};
  T_38110_21_br_prediction_bpd_predict_val = _RAND_3931[0:0];
  _RAND_3932 = {1{`RANDOM}};
  T_38110_21_br_prediction_bpd_predict_taken = _RAND_3932[0:0];
  _RAND_3933 = {1{`RANDOM}};
  T_38110_21_br_prediction_btb_hit = _RAND_3933[0:0];
  _RAND_3934 = {1{`RANDOM}};
  T_38110_21_br_prediction_btb_predicted = _RAND_3934[0:0];
  _RAND_3935 = {1{`RANDOM}};
  T_38110_21_br_prediction_is_br_or_jalr = _RAND_3935[0:0];
  _RAND_3936 = {1{`RANDOM}};
  T_38110_21_stat_brjmp_mispredicted = _RAND_3936[0:0];
  _RAND_3937 = {1{`RANDOM}};
  T_38110_21_stat_btb_made_pred = _RAND_3937[0:0];
  _RAND_3938 = {1{`RANDOM}};
  T_38110_21_stat_btb_mispredicted = _RAND_3938[0:0];
  _RAND_3939 = {1{`RANDOM}};
  T_38110_21_stat_bpd_made_pred = _RAND_3939[0:0];
  _RAND_3940 = {1{`RANDOM}};
  T_38110_21_stat_bpd_mispredicted = _RAND_3940[0:0];
  _RAND_3941 = {1{`RANDOM}};
  T_38110_21_fetch_pc_lob = _RAND_3941[2:0];
  _RAND_3942 = {1{`RANDOM}};
  T_38110_21_imm_packed = _RAND_3942[19:0];
  _RAND_3943 = {1{`RANDOM}};
  T_38110_21_csr_addr = _RAND_3943[11:0];
  _RAND_3944 = {1{`RANDOM}};
  T_38110_21_rob_idx = _RAND_3944[5:0];
  _RAND_3945 = {1{`RANDOM}};
  T_38110_21_ldq_idx = _RAND_3945[3:0];
  _RAND_3946 = {1{`RANDOM}};
  T_38110_21_stq_idx = _RAND_3946[3:0];
  _RAND_3947 = {1{`RANDOM}};
  T_38110_21_brob_idx = _RAND_3947[4:0];
  _RAND_3948 = {1{`RANDOM}};
  T_38110_21_pdst = _RAND_3948[6:0];
  _RAND_3949 = {1{`RANDOM}};
  T_38110_21_pop1 = _RAND_3949[6:0];
  _RAND_3950 = {1{`RANDOM}};
  T_38110_21_pop2 = _RAND_3950[6:0];
  _RAND_3951 = {1{`RANDOM}};
  T_38110_21_pop3 = _RAND_3951[6:0];
  _RAND_3952 = {1{`RANDOM}};
  T_38110_21_prs1_busy = _RAND_3952[0:0];
  _RAND_3953 = {1{`RANDOM}};
  T_38110_21_prs2_busy = _RAND_3953[0:0];
  _RAND_3954 = {1{`RANDOM}};
  T_38110_21_prs3_busy = _RAND_3954[0:0];
  _RAND_3955 = {1{`RANDOM}};
  T_38110_21_stale_pdst = _RAND_3955[6:0];
  _RAND_3956 = {1{`RANDOM}};
  T_38110_21_exception = _RAND_3956[0:0];
  _RAND_3957 = {2{`RANDOM}};
  T_38110_21_exc_cause = _RAND_3957[63:0];
  _RAND_3958 = {1{`RANDOM}};
  T_38110_21_bypassable = _RAND_3958[0:0];
  _RAND_3959 = {1{`RANDOM}};
  T_38110_21_mem_cmd = _RAND_3959[3:0];
  _RAND_3960 = {1{`RANDOM}};
  T_38110_21_mem_typ = _RAND_3960[2:0];
  _RAND_3961 = {1{`RANDOM}};
  T_38110_21_is_fence = _RAND_3961[0:0];
  _RAND_3962 = {1{`RANDOM}};
  T_38110_21_is_fencei = _RAND_3962[0:0];
  _RAND_3963 = {1{`RANDOM}};
  T_38110_21_is_store = _RAND_3963[0:0];
  _RAND_3964 = {1{`RANDOM}};
  T_38110_21_is_amo = _RAND_3964[0:0];
  _RAND_3965 = {1{`RANDOM}};
  T_38110_21_is_load = _RAND_3965[0:0];
  _RAND_3966 = {1{`RANDOM}};
  T_38110_21_is_unique = _RAND_3966[0:0];
  _RAND_3967 = {1{`RANDOM}};
  T_38110_21_flush_on_commit = _RAND_3967[0:0];
  _RAND_3968 = {1{`RANDOM}};
  T_38110_21_ldst = _RAND_3968[5:0];
  _RAND_3969 = {1{`RANDOM}};
  T_38110_21_lrs1 = _RAND_3969[5:0];
  _RAND_3970 = {1{`RANDOM}};
  T_38110_21_lrs2 = _RAND_3970[5:0];
  _RAND_3971 = {1{`RANDOM}};
  T_38110_21_lrs3 = _RAND_3971[5:0];
  _RAND_3972 = {1{`RANDOM}};
  T_38110_21_ldst_val = _RAND_3972[0:0];
  _RAND_3973 = {1{`RANDOM}};
  T_38110_21_dst_rtype = _RAND_3973[1:0];
  _RAND_3974 = {1{`RANDOM}};
  T_38110_21_lrs1_rtype = _RAND_3974[1:0];
  _RAND_3975 = {1{`RANDOM}};
  T_38110_21_lrs2_rtype = _RAND_3975[1:0];
  _RAND_3976 = {1{`RANDOM}};
  T_38110_21_frs3_en = _RAND_3976[0:0];
  _RAND_3977 = {1{`RANDOM}};
  T_38110_21_fp_val = _RAND_3977[0:0];
  _RAND_3978 = {1{`RANDOM}};
  T_38110_21_fp_single = _RAND_3978[0:0];
  _RAND_3979 = {1{`RANDOM}};
  T_38110_21_xcpt_if = _RAND_3979[0:0];
  _RAND_3980 = {1{`RANDOM}};
  T_38110_21_replay_if = _RAND_3980[0:0];
  _RAND_3981 = {2{`RANDOM}};
  T_38110_21_debug_wdata = _RAND_3981[63:0];
  _RAND_3982 = {1{`RANDOM}};
  T_38110_21_debug_events_fetch_seq = _RAND_3982[31:0];
  _RAND_3983 = {1{`RANDOM}};
  T_38110_22_valid = _RAND_3983[0:0];
  _RAND_3984 = {1{`RANDOM}};
  T_38110_22_iw_state = _RAND_3984[1:0];
  _RAND_3985 = {1{`RANDOM}};
  T_38110_22_uopc = _RAND_3985[8:0];
  _RAND_3986 = {1{`RANDOM}};
  T_38110_22_inst = _RAND_3986[31:0];
  _RAND_3987 = {2{`RANDOM}};
  T_38110_22_pc = _RAND_3987[39:0];
  _RAND_3988 = {1{`RANDOM}};
  T_38110_22_fu_code = _RAND_3988[7:0];
  _RAND_3989 = {1{`RANDOM}};
  T_38110_22_ctrl_br_type = _RAND_3989[3:0];
  _RAND_3990 = {1{`RANDOM}};
  T_38110_22_ctrl_op1_sel = _RAND_3990[1:0];
  _RAND_3991 = {1{`RANDOM}};
  T_38110_22_ctrl_op2_sel = _RAND_3991[2:0];
  _RAND_3992 = {1{`RANDOM}};
  T_38110_22_ctrl_imm_sel = _RAND_3992[2:0];
  _RAND_3993 = {1{`RANDOM}};
  T_38110_22_ctrl_op_fcn = _RAND_3993[3:0];
  _RAND_3994 = {1{`RANDOM}};
  T_38110_22_ctrl_fcn_dw = _RAND_3994[0:0];
  _RAND_3995 = {1{`RANDOM}};
  T_38110_22_ctrl_rf_wen = _RAND_3995[0:0];
  _RAND_3996 = {1{`RANDOM}};
  T_38110_22_ctrl_csr_cmd = _RAND_3996[2:0];
  _RAND_3997 = {1{`RANDOM}};
  T_38110_22_ctrl_is_load = _RAND_3997[0:0];
  _RAND_3998 = {1{`RANDOM}};
  T_38110_22_ctrl_is_sta = _RAND_3998[0:0];
  _RAND_3999 = {1{`RANDOM}};
  T_38110_22_ctrl_is_std = _RAND_3999[0:0];
  _RAND_4000 = {1{`RANDOM}};
  T_38110_22_wakeup_delay = _RAND_4000[1:0];
  _RAND_4001 = {1{`RANDOM}};
  T_38110_22_allocate_brtag = _RAND_4001[0:0];
  _RAND_4002 = {1{`RANDOM}};
  T_38110_22_is_br_or_jmp = _RAND_4002[0:0];
  _RAND_4003 = {1{`RANDOM}};
  T_38110_22_is_jump = _RAND_4003[0:0];
  _RAND_4004 = {1{`RANDOM}};
  T_38110_22_is_jal = _RAND_4004[0:0];
  _RAND_4005 = {1{`RANDOM}};
  T_38110_22_is_ret = _RAND_4005[0:0];
  _RAND_4006 = {1{`RANDOM}};
  T_38110_22_is_call = _RAND_4006[0:0];
  _RAND_4007 = {1{`RANDOM}};
  T_38110_22_br_mask = _RAND_4007[7:0];
  _RAND_4008 = {1{`RANDOM}};
  T_38110_22_br_tag = _RAND_4008[2:0];
  _RAND_4009 = {1{`RANDOM}};
  T_38110_22_br_prediction_bpd_predict_val = _RAND_4009[0:0];
  _RAND_4010 = {1{`RANDOM}};
  T_38110_22_br_prediction_bpd_predict_taken = _RAND_4010[0:0];
  _RAND_4011 = {1{`RANDOM}};
  T_38110_22_br_prediction_btb_hit = _RAND_4011[0:0];
  _RAND_4012 = {1{`RANDOM}};
  T_38110_22_br_prediction_btb_predicted = _RAND_4012[0:0];
  _RAND_4013 = {1{`RANDOM}};
  T_38110_22_br_prediction_is_br_or_jalr = _RAND_4013[0:0];
  _RAND_4014 = {1{`RANDOM}};
  T_38110_22_stat_brjmp_mispredicted = _RAND_4014[0:0];
  _RAND_4015 = {1{`RANDOM}};
  T_38110_22_stat_btb_made_pred = _RAND_4015[0:0];
  _RAND_4016 = {1{`RANDOM}};
  T_38110_22_stat_btb_mispredicted = _RAND_4016[0:0];
  _RAND_4017 = {1{`RANDOM}};
  T_38110_22_stat_bpd_made_pred = _RAND_4017[0:0];
  _RAND_4018 = {1{`RANDOM}};
  T_38110_22_stat_bpd_mispredicted = _RAND_4018[0:0];
  _RAND_4019 = {1{`RANDOM}};
  T_38110_22_fetch_pc_lob = _RAND_4019[2:0];
  _RAND_4020 = {1{`RANDOM}};
  T_38110_22_imm_packed = _RAND_4020[19:0];
  _RAND_4021 = {1{`RANDOM}};
  T_38110_22_csr_addr = _RAND_4021[11:0];
  _RAND_4022 = {1{`RANDOM}};
  T_38110_22_rob_idx = _RAND_4022[5:0];
  _RAND_4023 = {1{`RANDOM}};
  T_38110_22_ldq_idx = _RAND_4023[3:0];
  _RAND_4024 = {1{`RANDOM}};
  T_38110_22_stq_idx = _RAND_4024[3:0];
  _RAND_4025 = {1{`RANDOM}};
  T_38110_22_brob_idx = _RAND_4025[4:0];
  _RAND_4026 = {1{`RANDOM}};
  T_38110_22_pdst = _RAND_4026[6:0];
  _RAND_4027 = {1{`RANDOM}};
  T_38110_22_pop1 = _RAND_4027[6:0];
  _RAND_4028 = {1{`RANDOM}};
  T_38110_22_pop2 = _RAND_4028[6:0];
  _RAND_4029 = {1{`RANDOM}};
  T_38110_22_pop3 = _RAND_4029[6:0];
  _RAND_4030 = {1{`RANDOM}};
  T_38110_22_prs1_busy = _RAND_4030[0:0];
  _RAND_4031 = {1{`RANDOM}};
  T_38110_22_prs2_busy = _RAND_4031[0:0];
  _RAND_4032 = {1{`RANDOM}};
  T_38110_22_prs3_busy = _RAND_4032[0:0];
  _RAND_4033 = {1{`RANDOM}};
  T_38110_22_stale_pdst = _RAND_4033[6:0];
  _RAND_4034 = {1{`RANDOM}};
  T_38110_22_exception = _RAND_4034[0:0];
  _RAND_4035 = {2{`RANDOM}};
  T_38110_22_exc_cause = _RAND_4035[63:0];
  _RAND_4036 = {1{`RANDOM}};
  T_38110_22_bypassable = _RAND_4036[0:0];
  _RAND_4037 = {1{`RANDOM}};
  T_38110_22_mem_cmd = _RAND_4037[3:0];
  _RAND_4038 = {1{`RANDOM}};
  T_38110_22_mem_typ = _RAND_4038[2:0];
  _RAND_4039 = {1{`RANDOM}};
  T_38110_22_is_fence = _RAND_4039[0:0];
  _RAND_4040 = {1{`RANDOM}};
  T_38110_22_is_fencei = _RAND_4040[0:0];
  _RAND_4041 = {1{`RANDOM}};
  T_38110_22_is_store = _RAND_4041[0:0];
  _RAND_4042 = {1{`RANDOM}};
  T_38110_22_is_amo = _RAND_4042[0:0];
  _RAND_4043 = {1{`RANDOM}};
  T_38110_22_is_load = _RAND_4043[0:0];
  _RAND_4044 = {1{`RANDOM}};
  T_38110_22_is_unique = _RAND_4044[0:0];
  _RAND_4045 = {1{`RANDOM}};
  T_38110_22_flush_on_commit = _RAND_4045[0:0];
  _RAND_4046 = {1{`RANDOM}};
  T_38110_22_ldst = _RAND_4046[5:0];
  _RAND_4047 = {1{`RANDOM}};
  T_38110_22_lrs1 = _RAND_4047[5:0];
  _RAND_4048 = {1{`RANDOM}};
  T_38110_22_lrs2 = _RAND_4048[5:0];
  _RAND_4049 = {1{`RANDOM}};
  T_38110_22_lrs3 = _RAND_4049[5:0];
  _RAND_4050 = {1{`RANDOM}};
  T_38110_22_ldst_val = _RAND_4050[0:0];
  _RAND_4051 = {1{`RANDOM}};
  T_38110_22_dst_rtype = _RAND_4051[1:0];
  _RAND_4052 = {1{`RANDOM}};
  T_38110_22_lrs1_rtype = _RAND_4052[1:0];
  _RAND_4053 = {1{`RANDOM}};
  T_38110_22_lrs2_rtype = _RAND_4053[1:0];
  _RAND_4054 = {1{`RANDOM}};
  T_38110_22_frs3_en = _RAND_4054[0:0];
  _RAND_4055 = {1{`RANDOM}};
  T_38110_22_fp_val = _RAND_4055[0:0];
  _RAND_4056 = {1{`RANDOM}};
  T_38110_22_fp_single = _RAND_4056[0:0];
  _RAND_4057 = {1{`RANDOM}};
  T_38110_22_xcpt_if = _RAND_4057[0:0];
  _RAND_4058 = {1{`RANDOM}};
  T_38110_22_replay_if = _RAND_4058[0:0];
  _RAND_4059 = {2{`RANDOM}};
  T_38110_22_debug_wdata = _RAND_4059[63:0];
  _RAND_4060 = {1{`RANDOM}};
  T_38110_22_debug_events_fetch_seq = _RAND_4060[31:0];
  _RAND_4061 = {1{`RANDOM}};
  T_38110_23_valid = _RAND_4061[0:0];
  _RAND_4062 = {1{`RANDOM}};
  T_38110_23_iw_state = _RAND_4062[1:0];
  _RAND_4063 = {1{`RANDOM}};
  T_38110_23_uopc = _RAND_4063[8:0];
  _RAND_4064 = {1{`RANDOM}};
  T_38110_23_inst = _RAND_4064[31:0];
  _RAND_4065 = {2{`RANDOM}};
  T_38110_23_pc = _RAND_4065[39:0];
  _RAND_4066 = {1{`RANDOM}};
  T_38110_23_fu_code = _RAND_4066[7:0];
  _RAND_4067 = {1{`RANDOM}};
  T_38110_23_ctrl_br_type = _RAND_4067[3:0];
  _RAND_4068 = {1{`RANDOM}};
  T_38110_23_ctrl_op1_sel = _RAND_4068[1:0];
  _RAND_4069 = {1{`RANDOM}};
  T_38110_23_ctrl_op2_sel = _RAND_4069[2:0];
  _RAND_4070 = {1{`RANDOM}};
  T_38110_23_ctrl_imm_sel = _RAND_4070[2:0];
  _RAND_4071 = {1{`RANDOM}};
  T_38110_23_ctrl_op_fcn = _RAND_4071[3:0];
  _RAND_4072 = {1{`RANDOM}};
  T_38110_23_ctrl_fcn_dw = _RAND_4072[0:0];
  _RAND_4073 = {1{`RANDOM}};
  T_38110_23_ctrl_rf_wen = _RAND_4073[0:0];
  _RAND_4074 = {1{`RANDOM}};
  T_38110_23_ctrl_csr_cmd = _RAND_4074[2:0];
  _RAND_4075 = {1{`RANDOM}};
  T_38110_23_ctrl_is_load = _RAND_4075[0:0];
  _RAND_4076 = {1{`RANDOM}};
  T_38110_23_ctrl_is_sta = _RAND_4076[0:0];
  _RAND_4077 = {1{`RANDOM}};
  T_38110_23_ctrl_is_std = _RAND_4077[0:0];
  _RAND_4078 = {1{`RANDOM}};
  T_38110_23_wakeup_delay = _RAND_4078[1:0];
  _RAND_4079 = {1{`RANDOM}};
  T_38110_23_allocate_brtag = _RAND_4079[0:0];
  _RAND_4080 = {1{`RANDOM}};
  T_38110_23_is_br_or_jmp = _RAND_4080[0:0];
  _RAND_4081 = {1{`RANDOM}};
  T_38110_23_is_jump = _RAND_4081[0:0];
  _RAND_4082 = {1{`RANDOM}};
  T_38110_23_is_jal = _RAND_4082[0:0];
  _RAND_4083 = {1{`RANDOM}};
  T_38110_23_is_ret = _RAND_4083[0:0];
  _RAND_4084 = {1{`RANDOM}};
  T_38110_23_is_call = _RAND_4084[0:0];
  _RAND_4085 = {1{`RANDOM}};
  T_38110_23_br_mask = _RAND_4085[7:0];
  _RAND_4086 = {1{`RANDOM}};
  T_38110_23_br_tag = _RAND_4086[2:0];
  _RAND_4087 = {1{`RANDOM}};
  T_38110_23_br_prediction_bpd_predict_val = _RAND_4087[0:0];
  _RAND_4088 = {1{`RANDOM}};
  T_38110_23_br_prediction_bpd_predict_taken = _RAND_4088[0:0];
  _RAND_4089 = {1{`RANDOM}};
  T_38110_23_br_prediction_btb_hit = _RAND_4089[0:0];
  _RAND_4090 = {1{`RANDOM}};
  T_38110_23_br_prediction_btb_predicted = _RAND_4090[0:0];
  _RAND_4091 = {1{`RANDOM}};
  T_38110_23_br_prediction_is_br_or_jalr = _RAND_4091[0:0];
  _RAND_4092 = {1{`RANDOM}};
  T_38110_23_stat_brjmp_mispredicted = _RAND_4092[0:0];
  _RAND_4093 = {1{`RANDOM}};
  T_38110_23_stat_btb_made_pred = _RAND_4093[0:0];
  _RAND_4094 = {1{`RANDOM}};
  T_38110_23_stat_btb_mispredicted = _RAND_4094[0:0];
  _RAND_4095 = {1{`RANDOM}};
  T_38110_23_stat_bpd_made_pred = _RAND_4095[0:0];
  _RAND_4096 = {1{`RANDOM}};
  T_38110_23_stat_bpd_mispredicted = _RAND_4096[0:0];
  _RAND_4097 = {1{`RANDOM}};
  T_38110_23_fetch_pc_lob = _RAND_4097[2:0];
  _RAND_4098 = {1{`RANDOM}};
  T_38110_23_imm_packed = _RAND_4098[19:0];
  _RAND_4099 = {1{`RANDOM}};
  T_38110_23_csr_addr = _RAND_4099[11:0];
  _RAND_4100 = {1{`RANDOM}};
  T_38110_23_rob_idx = _RAND_4100[5:0];
  _RAND_4101 = {1{`RANDOM}};
  T_38110_23_ldq_idx = _RAND_4101[3:0];
  _RAND_4102 = {1{`RANDOM}};
  T_38110_23_stq_idx = _RAND_4102[3:0];
  _RAND_4103 = {1{`RANDOM}};
  T_38110_23_brob_idx = _RAND_4103[4:0];
  _RAND_4104 = {1{`RANDOM}};
  T_38110_23_pdst = _RAND_4104[6:0];
  _RAND_4105 = {1{`RANDOM}};
  T_38110_23_pop1 = _RAND_4105[6:0];
  _RAND_4106 = {1{`RANDOM}};
  T_38110_23_pop2 = _RAND_4106[6:0];
  _RAND_4107 = {1{`RANDOM}};
  T_38110_23_pop3 = _RAND_4107[6:0];
  _RAND_4108 = {1{`RANDOM}};
  T_38110_23_prs1_busy = _RAND_4108[0:0];
  _RAND_4109 = {1{`RANDOM}};
  T_38110_23_prs2_busy = _RAND_4109[0:0];
  _RAND_4110 = {1{`RANDOM}};
  T_38110_23_prs3_busy = _RAND_4110[0:0];
  _RAND_4111 = {1{`RANDOM}};
  T_38110_23_stale_pdst = _RAND_4111[6:0];
  _RAND_4112 = {1{`RANDOM}};
  T_38110_23_exception = _RAND_4112[0:0];
  _RAND_4113 = {2{`RANDOM}};
  T_38110_23_exc_cause = _RAND_4113[63:0];
  _RAND_4114 = {1{`RANDOM}};
  T_38110_23_bypassable = _RAND_4114[0:0];
  _RAND_4115 = {1{`RANDOM}};
  T_38110_23_mem_cmd = _RAND_4115[3:0];
  _RAND_4116 = {1{`RANDOM}};
  T_38110_23_mem_typ = _RAND_4116[2:0];
  _RAND_4117 = {1{`RANDOM}};
  T_38110_23_is_fence = _RAND_4117[0:0];
  _RAND_4118 = {1{`RANDOM}};
  T_38110_23_is_fencei = _RAND_4118[0:0];
  _RAND_4119 = {1{`RANDOM}};
  T_38110_23_is_store = _RAND_4119[0:0];
  _RAND_4120 = {1{`RANDOM}};
  T_38110_23_is_amo = _RAND_4120[0:0];
  _RAND_4121 = {1{`RANDOM}};
  T_38110_23_is_load = _RAND_4121[0:0];
  _RAND_4122 = {1{`RANDOM}};
  T_38110_23_is_unique = _RAND_4122[0:0];
  _RAND_4123 = {1{`RANDOM}};
  T_38110_23_flush_on_commit = _RAND_4123[0:0];
  _RAND_4124 = {1{`RANDOM}};
  T_38110_23_ldst = _RAND_4124[5:0];
  _RAND_4125 = {1{`RANDOM}};
  T_38110_23_lrs1 = _RAND_4125[5:0];
  _RAND_4126 = {1{`RANDOM}};
  T_38110_23_lrs2 = _RAND_4126[5:0];
  _RAND_4127 = {1{`RANDOM}};
  T_38110_23_lrs3 = _RAND_4127[5:0];
  _RAND_4128 = {1{`RANDOM}};
  T_38110_23_ldst_val = _RAND_4128[0:0];
  _RAND_4129 = {1{`RANDOM}};
  T_38110_23_dst_rtype = _RAND_4129[1:0];
  _RAND_4130 = {1{`RANDOM}};
  T_38110_23_lrs1_rtype = _RAND_4130[1:0];
  _RAND_4131 = {1{`RANDOM}};
  T_38110_23_lrs2_rtype = _RAND_4131[1:0];
  _RAND_4132 = {1{`RANDOM}};
  T_38110_23_frs3_en = _RAND_4132[0:0];
  _RAND_4133 = {1{`RANDOM}};
  T_38110_23_fp_val = _RAND_4133[0:0];
  _RAND_4134 = {1{`RANDOM}};
  T_38110_23_fp_single = _RAND_4134[0:0];
  _RAND_4135 = {1{`RANDOM}};
  T_38110_23_xcpt_if = _RAND_4135[0:0];
  _RAND_4136 = {1{`RANDOM}};
  T_38110_23_replay_if = _RAND_4136[0:0];
  _RAND_4137 = {2{`RANDOM}};
  T_38110_23_debug_wdata = _RAND_4137[63:0];
  _RAND_4138 = {1{`RANDOM}};
  T_38110_23_debug_events_fetch_seq = _RAND_4138[31:0];
  _RAND_4139 = {1{`RANDOM}};
  T_47576 = _RAND_4139[0:0];
  _RAND_4140 = {1{`RANDOM}};
  T_47616 = _RAND_4140[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
