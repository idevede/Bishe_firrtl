module HwachaSequencer(
  input         clock,
  input         reset,
  output        io_op_ready,
  input         io_op_valid,
  input  [9:0]  io_op_bits_fn_union,
  input  [63:0] io_op_bits_sreg_ss1,
  input  [63:0] io_op_bits_sreg_ss2,
  input  [63:0] io_op_bits_sreg_ss3,
  input  [3:0]  io_op_bits_base_vp_id,
  input         io_op_bits_base_vp_valid,
  input         io_op_bits_base_vp_scalar,
  input         io_op_bits_base_vp_pred,
  input  [7:0]  io_op_bits_base_vs1_id,
  input         io_op_bits_base_vs1_valid,
  input         io_op_bits_base_vs1_scalar,
  input         io_op_bits_base_vs1_pred,
  input  [1:0]  io_op_bits_base_vs1_prec,
  input  [7:0]  io_op_bits_base_vs2_id,
  input         io_op_bits_base_vs2_valid,
  input         io_op_bits_base_vs2_scalar,
  input         io_op_bits_base_vs2_pred,
  input  [1:0]  io_op_bits_base_vs2_prec,
  input  [7:0]  io_op_bits_base_vs3_id,
  input         io_op_bits_base_vs3_valid,
  input         io_op_bits_base_vs3_scalar,
  input         io_op_bits_base_vs3_pred,
  input  [1:0]  io_op_bits_base_vs3_prec,
  input  [7:0]  io_op_bits_base_vd_id,
  input         io_op_bits_base_vd_valid,
  input         io_op_bits_base_vd_scalar,
  input         io_op_bits_base_vd_pred,
  input  [1:0]  io_op_bits_base_vd_prec,
  input  [7:0]  io_op_bits_reg_vp_id,
  input  [7:0]  io_op_bits_reg_vs1_id,
  input  [7:0]  io_op_bits_reg_vs2_id,
  input  [7:0]  io_op_bits_reg_vs3_id,
  input  [7:0]  io_op_bits_reg_vd_id,
  input         io_op_bits_active_vint,
  input         io_op_bits_active_vipred,
  input         io_op_bits_active_vimul,
  input         io_op_bits_active_vidiv,
  input         io_op_bits_active_vfma,
  input         io_op_bits_active_vfdiv,
  input         io_op_bits_active_vfcmp,
  input         io_op_bits_active_vfconv,
  input         io_op_bits_active_vrpred,
  input         io_op_bits_active_vrfirst,
  input         io_op_bits_active_vamo,
  input         io_op_bits_active_vldx,
  input         io_op_bits_active_vstx,
  input         io_op_bits_active_vld,
  input         io_op_bits_active_vst,
  output        io_master_state_valid_0,
  output        io_master_state_valid_1,
  output        io_master_state_valid_2,
  output        io_master_state_valid_3,
  output        io_master_state_valid_4,
  output        io_master_state_valid_5,
  output        io_master_state_valid_6,
  output        io_master_state_valid_7,
  output [9:0]  io_master_state_e_0_fn_union,
  output [63:0] io_master_state_e_0_sreg_ss1,
  output [63:0] io_master_state_e_0_sreg_ss2,
  output [63:0] io_master_state_e_0_sreg_ss3,
  output [3:0]  io_master_state_e_0_base_vp_id,
  output        io_master_state_e_0_base_vp_valid,
  output        io_master_state_e_0_base_vp_scalar,
  output        io_master_state_e_0_base_vp_pred,
  output [7:0]  io_master_state_e_0_base_vs1_id,
  output        io_master_state_e_0_base_vs1_valid,
  output        io_master_state_e_0_base_vs1_scalar,
  output        io_master_state_e_0_base_vs1_pred,
  output [1:0]  io_master_state_e_0_base_vs1_prec,
  output [7:0]  io_master_state_e_0_base_vs2_id,
  output        io_master_state_e_0_base_vs2_valid,
  output        io_master_state_e_0_base_vs2_scalar,
  output        io_master_state_e_0_base_vs2_pred,
  output [1:0]  io_master_state_e_0_base_vs2_prec,
  output [7:0]  io_master_state_e_0_base_vs3_id,
  output        io_master_state_e_0_base_vs3_valid,
  output        io_master_state_e_0_base_vs3_scalar,
  output        io_master_state_e_0_base_vs3_pred,
  output [1:0]  io_master_state_e_0_base_vs3_prec,
  output [7:0]  io_master_state_e_0_base_vd_id,
  output        io_master_state_e_0_base_vd_valid,
  output        io_master_state_e_0_base_vd_scalar,
  output        io_master_state_e_0_base_vd_pred,
  output [1:0]  io_master_state_e_0_base_vd_prec,
  output        io_master_state_e_0_rate,
  output        io_master_state_e_0_active_viu,
  output        io_master_state_e_0_active_vipu,
  output        io_master_state_e_0_active_vimu,
  output        io_master_state_e_0_active_vidu,
  output        io_master_state_e_0_active_vfmu,
  output        io_master_state_e_0_active_vfdu,
  output        io_master_state_e_0_active_vfcu,
  output        io_master_state_e_0_active_vfvu,
  output        io_master_state_e_0_active_vrpu,
  output        io_master_state_e_0_active_vrfu,
  output        io_master_state_e_0_active_vpu,
  output        io_master_state_e_0_active_vgu,
  output        io_master_state_e_0_active_vcu,
  output        io_master_state_e_0_active_vlu,
  output        io_master_state_e_0_active_vsu,
  output        io_master_state_e_0_active_vqu,
  output        io_master_state_e_0_raw_0,
  output        io_master_state_e_0_raw_1,
  output        io_master_state_e_0_raw_2,
  output        io_master_state_e_0_raw_3,
  output        io_master_state_e_0_raw_4,
  output        io_master_state_e_0_raw_5,
  output        io_master_state_e_0_raw_6,
  output        io_master_state_e_0_raw_7,
  output        io_master_state_e_0_war_0,
  output        io_master_state_e_0_war_1,
  output        io_master_state_e_0_war_2,
  output        io_master_state_e_0_war_3,
  output        io_master_state_e_0_war_4,
  output        io_master_state_e_0_war_5,
  output        io_master_state_e_0_war_6,
  output        io_master_state_e_0_war_7,
  output        io_master_state_e_0_waw_0,
  output        io_master_state_e_0_waw_1,
  output        io_master_state_e_0_waw_2,
  output        io_master_state_e_0_waw_3,
  output        io_master_state_e_0_waw_4,
  output        io_master_state_e_0_waw_5,
  output        io_master_state_e_0_waw_6,
  output        io_master_state_e_0_waw_7,
  output        io_master_state_e_0_last,
  output [1:0]  io_master_state_e_0_rports,
  output [3:0]  io_master_state_e_0_wport_sram,
  output [2:0]  io_master_state_e_0_wport_pred,
  output [9:0]  io_master_state_e_1_fn_union,
  output [63:0] io_master_state_e_1_sreg_ss1,
  output [63:0] io_master_state_e_1_sreg_ss2,
  output [63:0] io_master_state_e_1_sreg_ss3,
  output [3:0]  io_master_state_e_1_base_vp_id,
  output        io_master_state_e_1_base_vp_valid,
  output        io_master_state_e_1_base_vp_scalar,
  output        io_master_state_e_1_base_vp_pred,
  output [7:0]  io_master_state_e_1_base_vs1_id,
  output        io_master_state_e_1_base_vs1_valid,
  output        io_master_state_e_1_base_vs1_scalar,
  output        io_master_state_e_1_base_vs1_pred,
  output [1:0]  io_master_state_e_1_base_vs1_prec,
  output [7:0]  io_master_state_e_1_base_vs2_id,
  output        io_master_state_e_1_base_vs2_valid,
  output        io_master_state_e_1_base_vs2_scalar,
  output        io_master_state_e_1_base_vs2_pred,
  output [1:0]  io_master_state_e_1_base_vs2_prec,
  output [7:0]  io_master_state_e_1_base_vs3_id,
  output        io_master_state_e_1_base_vs3_valid,
  output        io_master_state_e_1_base_vs3_scalar,
  output        io_master_state_e_1_base_vs3_pred,
  output [1:0]  io_master_state_e_1_base_vs3_prec,
  output [7:0]  io_master_state_e_1_base_vd_id,
  output        io_master_state_e_1_base_vd_valid,
  output        io_master_state_e_1_base_vd_scalar,
  output        io_master_state_e_1_base_vd_pred,
  output [1:0]  io_master_state_e_1_base_vd_prec,
  output        io_master_state_e_1_rate,
  output        io_master_state_e_1_active_viu,
  output        io_master_state_e_1_active_vipu,
  output        io_master_state_e_1_active_vimu,
  output        io_master_state_e_1_active_vidu,
  output        io_master_state_e_1_active_vfmu,
  output        io_master_state_e_1_active_vfdu,
  output        io_master_state_e_1_active_vfcu,
  output        io_master_state_e_1_active_vfvu,
  output        io_master_state_e_1_active_vrpu,
  output        io_master_state_e_1_active_vrfu,
  output        io_master_state_e_1_active_vpu,
  output        io_master_state_e_1_active_vgu,
  output        io_master_state_e_1_active_vcu,
  output        io_master_state_e_1_active_vlu,
  output        io_master_state_e_1_active_vsu,
  output        io_master_state_e_1_active_vqu,
  output        io_master_state_e_1_raw_0,
  output        io_master_state_e_1_raw_1,
  output        io_master_state_e_1_raw_2,
  output        io_master_state_e_1_raw_3,
  output        io_master_state_e_1_raw_4,
  output        io_master_state_e_1_raw_5,
  output        io_master_state_e_1_raw_6,
  output        io_master_state_e_1_raw_7,
  output        io_master_state_e_1_war_0,
  output        io_master_state_e_1_war_1,
  output        io_master_state_e_1_war_2,
  output        io_master_state_e_1_war_3,
  output        io_master_state_e_1_war_4,
  output        io_master_state_e_1_war_5,
  output        io_master_state_e_1_war_6,
  output        io_master_state_e_1_war_7,
  output        io_master_state_e_1_waw_0,
  output        io_master_state_e_1_waw_1,
  output        io_master_state_e_1_waw_2,
  output        io_master_state_e_1_waw_3,
  output        io_master_state_e_1_waw_4,
  output        io_master_state_e_1_waw_5,
  output        io_master_state_e_1_waw_6,
  output        io_master_state_e_1_waw_7,
  output        io_master_state_e_1_last,
  output [1:0]  io_master_state_e_1_rports,
  output [3:0]  io_master_state_e_1_wport_sram,
  output [2:0]  io_master_state_e_1_wport_pred,
  output [9:0]  io_master_state_e_2_fn_union,
  output [63:0] io_master_state_e_2_sreg_ss1,
  output [63:0] io_master_state_e_2_sreg_ss2,
  output [63:0] io_master_state_e_2_sreg_ss3,
  output [3:0]  io_master_state_e_2_base_vp_id,
  output        io_master_state_e_2_base_vp_valid,
  output        io_master_state_e_2_base_vp_scalar,
  output        io_master_state_e_2_base_vp_pred,
  output [7:0]  io_master_state_e_2_base_vs1_id,
  output        io_master_state_e_2_base_vs1_valid,
  output        io_master_state_e_2_base_vs1_scalar,
  output        io_master_state_e_2_base_vs1_pred,
  output [1:0]  io_master_state_e_2_base_vs1_prec,
  output [7:0]  io_master_state_e_2_base_vs2_id,
  output        io_master_state_e_2_base_vs2_valid,
  output        io_master_state_e_2_base_vs2_scalar,
  output        io_master_state_e_2_base_vs2_pred,
  output [1:0]  io_master_state_e_2_base_vs2_prec,
  output [7:0]  io_master_state_e_2_base_vs3_id,
  output        io_master_state_e_2_base_vs3_valid,
  output        io_master_state_e_2_base_vs3_scalar,
  output        io_master_state_e_2_base_vs3_pred,
  output [1:0]  io_master_state_e_2_base_vs3_prec,
  output [7:0]  io_master_state_e_2_base_vd_id,
  output        io_master_state_e_2_base_vd_valid,
  output        io_master_state_e_2_base_vd_scalar,
  output        io_master_state_e_2_base_vd_pred,
  output [1:0]  io_master_state_e_2_base_vd_prec,
  output        io_master_state_e_2_rate,
  output        io_master_state_e_2_active_viu,
  output        io_master_state_e_2_active_vipu,
  output        io_master_state_e_2_active_vimu,
  output        io_master_state_e_2_active_vidu,
  output        io_master_state_e_2_active_vfmu,
  output        io_master_state_e_2_active_vfdu,
  output        io_master_state_e_2_active_vfcu,
  output        io_master_state_e_2_active_vfvu,
  output        io_master_state_e_2_active_vrpu,
  output        io_master_state_e_2_active_vrfu,
  output        io_master_state_e_2_active_vpu,
  output        io_master_state_e_2_active_vgu,
  output        io_master_state_e_2_active_vcu,
  output        io_master_state_e_2_active_vlu,
  output        io_master_state_e_2_active_vsu,
  output        io_master_state_e_2_active_vqu,
  output        io_master_state_e_2_raw_0,
  output        io_master_state_e_2_raw_1,
  output        io_master_state_e_2_raw_2,
  output        io_master_state_e_2_raw_3,
  output        io_master_state_e_2_raw_4,
  output        io_master_state_e_2_raw_5,
  output        io_master_state_e_2_raw_6,
  output        io_master_state_e_2_raw_7,
  output        io_master_state_e_2_war_0,
  output        io_master_state_e_2_war_1,
  output        io_master_state_e_2_war_2,
  output        io_master_state_e_2_war_3,
  output        io_master_state_e_2_war_4,
  output        io_master_state_e_2_war_5,
  output        io_master_state_e_2_war_6,
  output        io_master_state_e_2_war_7,
  output        io_master_state_e_2_waw_0,
  output        io_master_state_e_2_waw_1,
  output        io_master_state_e_2_waw_2,
  output        io_master_state_e_2_waw_3,
  output        io_master_state_e_2_waw_4,
  output        io_master_state_e_2_waw_5,
  output        io_master_state_e_2_waw_6,
  output        io_master_state_e_2_waw_7,
  output        io_master_state_e_2_last,
  output [1:0]  io_master_state_e_2_rports,
  output [3:0]  io_master_state_e_2_wport_sram,
  output [2:0]  io_master_state_e_2_wport_pred,
  output [9:0]  io_master_state_e_3_fn_union,
  output [63:0] io_master_state_e_3_sreg_ss1,
  output [63:0] io_master_state_e_3_sreg_ss2,
  output [63:0] io_master_state_e_3_sreg_ss3,
  output [3:0]  io_master_state_e_3_base_vp_id,
  output        io_master_state_e_3_base_vp_valid,
  output        io_master_state_e_3_base_vp_scalar,
  output        io_master_state_e_3_base_vp_pred,
  output [7:0]  io_master_state_e_3_base_vs1_id,
  output        io_master_state_e_3_base_vs1_valid,
  output        io_master_state_e_3_base_vs1_scalar,
  output        io_master_state_e_3_base_vs1_pred,
  output [1:0]  io_master_state_e_3_base_vs1_prec,
  output [7:0]  io_master_state_e_3_base_vs2_id,
  output        io_master_state_e_3_base_vs2_valid,
  output        io_master_state_e_3_base_vs2_scalar,
  output        io_master_state_e_3_base_vs2_pred,
  output [1:0]  io_master_state_e_3_base_vs2_prec,
  output [7:0]  io_master_state_e_3_base_vs3_id,
  output        io_master_state_e_3_base_vs3_valid,
  output        io_master_state_e_3_base_vs3_scalar,
  output        io_master_state_e_3_base_vs3_pred,
  output [1:0]  io_master_state_e_3_base_vs3_prec,
  output [7:0]  io_master_state_e_3_base_vd_id,
  output        io_master_state_e_3_base_vd_valid,
  output        io_master_state_e_3_base_vd_scalar,
  output        io_master_state_e_3_base_vd_pred,
  output [1:0]  io_master_state_e_3_base_vd_prec,
  output        io_master_state_e_3_rate,
  output        io_master_state_e_3_active_viu,
  output        io_master_state_e_3_active_vipu,
  output        io_master_state_e_3_active_vimu,
  output        io_master_state_e_3_active_vidu,
  output        io_master_state_e_3_active_vfmu,
  output        io_master_state_e_3_active_vfdu,
  output        io_master_state_e_3_active_vfcu,
  output        io_master_state_e_3_active_vfvu,
  output        io_master_state_e_3_active_vrpu,
  output        io_master_state_e_3_active_vrfu,
  output        io_master_state_e_3_active_vpu,
  output        io_master_state_e_3_active_vgu,
  output        io_master_state_e_3_active_vcu,
  output        io_master_state_e_3_active_vlu,
  output        io_master_state_e_3_active_vsu,
  output        io_master_state_e_3_active_vqu,
  output        io_master_state_e_3_raw_0,
  output        io_master_state_e_3_raw_1,
  output        io_master_state_e_3_raw_2,
  output        io_master_state_e_3_raw_3,
  output        io_master_state_e_3_raw_4,
  output        io_master_state_e_3_raw_5,
  output        io_master_state_e_3_raw_6,
  output        io_master_state_e_3_raw_7,
  output        io_master_state_e_3_war_0,
  output        io_master_state_e_3_war_1,
  output        io_master_state_e_3_war_2,
  output        io_master_state_e_3_war_3,
  output        io_master_state_e_3_war_4,
  output        io_master_state_e_3_war_5,
  output        io_master_state_e_3_war_6,
  output        io_master_state_e_3_war_7,
  output        io_master_state_e_3_waw_0,
  output        io_master_state_e_3_waw_1,
  output        io_master_state_e_3_waw_2,
  output        io_master_state_e_3_waw_3,
  output        io_master_state_e_3_waw_4,
  output        io_master_state_e_3_waw_5,
  output        io_master_state_e_3_waw_6,
  output        io_master_state_e_3_waw_7,
  output        io_master_state_e_3_last,
  output [1:0]  io_master_state_e_3_rports,
  output [3:0]  io_master_state_e_3_wport_sram,
  output [2:0]  io_master_state_e_3_wport_pred,
  output [9:0]  io_master_state_e_4_fn_union,
  output [63:0] io_master_state_e_4_sreg_ss1,
  output [63:0] io_master_state_e_4_sreg_ss2,
  output [63:0] io_master_state_e_4_sreg_ss3,
  output [3:0]  io_master_state_e_4_base_vp_id,
  output        io_master_state_e_4_base_vp_valid,
  output        io_master_state_e_4_base_vp_scalar,
  output        io_master_state_e_4_base_vp_pred,
  output [7:0]  io_master_state_e_4_base_vs1_id,
  output        io_master_state_e_4_base_vs1_valid,
  output        io_master_state_e_4_base_vs1_scalar,
  output        io_master_state_e_4_base_vs1_pred,
  output [1:0]  io_master_state_e_4_base_vs1_prec,
  output [7:0]  io_master_state_e_4_base_vs2_id,
  output        io_master_state_e_4_base_vs2_valid,
  output        io_master_state_e_4_base_vs2_scalar,
  output        io_master_state_e_4_base_vs2_pred,
  output [1:0]  io_master_state_e_4_base_vs2_prec,
  output [7:0]  io_master_state_e_4_base_vs3_id,
  output        io_master_state_e_4_base_vs3_valid,
  output        io_master_state_e_4_base_vs3_scalar,
  output        io_master_state_e_4_base_vs3_pred,
  output [1:0]  io_master_state_e_4_base_vs3_prec,
  output [7:0]  io_master_state_e_4_base_vd_id,
  output        io_master_state_e_4_base_vd_valid,
  output        io_master_state_e_4_base_vd_scalar,
  output        io_master_state_e_4_base_vd_pred,
  output [1:0]  io_master_state_e_4_base_vd_prec,
  output        io_master_state_e_4_rate,
  output        io_master_state_e_4_active_viu,
  output        io_master_state_e_4_active_vipu,
  output        io_master_state_e_4_active_vimu,
  output        io_master_state_e_4_active_vidu,
  output        io_master_state_e_4_active_vfmu,
  output        io_master_state_e_4_active_vfdu,
  output        io_master_state_e_4_active_vfcu,
  output        io_master_state_e_4_active_vfvu,
  output        io_master_state_e_4_active_vrpu,
  output        io_master_state_e_4_active_vrfu,
  output        io_master_state_e_4_active_vpu,
  output        io_master_state_e_4_active_vgu,
  output        io_master_state_e_4_active_vcu,
  output        io_master_state_e_4_active_vlu,
  output        io_master_state_e_4_active_vsu,
  output        io_master_state_e_4_active_vqu,
  output        io_master_state_e_4_raw_0,
  output        io_master_state_e_4_raw_1,
  output        io_master_state_e_4_raw_2,
  output        io_master_state_e_4_raw_3,
  output        io_master_state_e_4_raw_4,
  output        io_master_state_e_4_raw_5,
  output        io_master_state_e_4_raw_6,
  output        io_master_state_e_4_raw_7,
  output        io_master_state_e_4_war_0,
  output        io_master_state_e_4_war_1,
  output        io_master_state_e_4_war_2,
  output        io_master_state_e_4_war_3,
  output        io_master_state_e_4_war_4,
  output        io_master_state_e_4_war_5,
  output        io_master_state_e_4_war_6,
  output        io_master_state_e_4_war_7,
  output        io_master_state_e_4_waw_0,
  output        io_master_state_e_4_waw_1,
  output        io_master_state_e_4_waw_2,
  output        io_master_state_e_4_waw_3,
  output        io_master_state_e_4_waw_4,
  output        io_master_state_e_4_waw_5,
  output        io_master_state_e_4_waw_6,
  output        io_master_state_e_4_waw_7,
  output        io_master_state_e_4_last,
  output [1:0]  io_master_state_e_4_rports,
  output [3:0]  io_master_state_e_4_wport_sram,
  output [2:0]  io_master_state_e_4_wport_pred,
  output [9:0]  io_master_state_e_5_fn_union,
  output [63:0] io_master_state_e_5_sreg_ss1,
  output [63:0] io_master_state_e_5_sreg_ss2,
  output [63:0] io_master_state_e_5_sreg_ss3,
  output [3:0]  io_master_state_e_5_base_vp_id,
  output        io_master_state_e_5_base_vp_valid,
  output        io_master_state_e_5_base_vp_scalar,
  output        io_master_state_e_5_base_vp_pred,
  output [7:0]  io_master_state_e_5_base_vs1_id,
  output        io_master_state_e_5_base_vs1_valid,
  output        io_master_state_e_5_base_vs1_scalar,
  output        io_master_state_e_5_base_vs1_pred,
  output [1:0]  io_master_state_e_5_base_vs1_prec,
  output [7:0]  io_master_state_e_5_base_vs2_id,
  output        io_master_state_e_5_base_vs2_valid,
  output        io_master_state_e_5_base_vs2_scalar,
  output        io_master_state_e_5_base_vs2_pred,
  output [1:0]  io_master_state_e_5_base_vs2_prec,
  output [7:0]  io_master_state_e_5_base_vs3_id,
  output        io_master_state_e_5_base_vs3_valid,
  output        io_master_state_e_5_base_vs3_scalar,
  output        io_master_state_e_5_base_vs3_pred,
  output [1:0]  io_master_state_e_5_base_vs3_prec,
  output [7:0]  io_master_state_e_5_base_vd_id,
  output        io_master_state_e_5_base_vd_valid,
  output        io_master_state_e_5_base_vd_scalar,
  output        io_master_state_e_5_base_vd_pred,
  output [1:0]  io_master_state_e_5_base_vd_prec,
  output        io_master_state_e_5_rate,
  output        io_master_state_e_5_active_viu,
  output        io_master_state_e_5_active_vipu,
  output        io_master_state_e_5_active_vimu,
  output        io_master_state_e_5_active_vidu,
  output        io_master_state_e_5_active_vfmu,
  output        io_master_state_e_5_active_vfdu,
  output        io_master_state_e_5_active_vfcu,
  output        io_master_state_e_5_active_vfvu,
  output        io_master_state_e_5_active_vrpu,
  output        io_master_state_e_5_active_vrfu,
  output        io_master_state_e_5_active_vpu,
  output        io_master_state_e_5_active_vgu,
  output        io_master_state_e_5_active_vcu,
  output        io_master_state_e_5_active_vlu,
  output        io_master_state_e_5_active_vsu,
  output        io_master_state_e_5_active_vqu,
  output        io_master_state_e_5_raw_0,
  output        io_master_state_e_5_raw_1,
  output        io_master_state_e_5_raw_2,
  output        io_master_state_e_5_raw_3,
  output        io_master_state_e_5_raw_4,
  output        io_master_state_e_5_raw_5,
  output        io_master_state_e_5_raw_6,
  output        io_master_state_e_5_raw_7,
  output        io_master_state_e_5_war_0,
  output        io_master_state_e_5_war_1,
  output        io_master_state_e_5_war_2,
  output        io_master_state_e_5_war_3,
  output        io_master_state_e_5_war_4,
  output        io_master_state_e_5_war_5,
  output        io_master_state_e_5_war_6,
  output        io_master_state_e_5_war_7,
  output        io_master_state_e_5_waw_0,
  output        io_master_state_e_5_waw_1,
  output        io_master_state_e_5_waw_2,
  output        io_master_state_e_5_waw_3,
  output        io_master_state_e_5_waw_4,
  output        io_master_state_e_5_waw_5,
  output        io_master_state_e_5_waw_6,
  output        io_master_state_e_5_waw_7,
  output        io_master_state_e_5_last,
  output [1:0]  io_master_state_e_5_rports,
  output [3:0]  io_master_state_e_5_wport_sram,
  output [2:0]  io_master_state_e_5_wport_pred,
  output [9:0]  io_master_state_e_6_fn_union,
  output [63:0] io_master_state_e_6_sreg_ss1,
  output [63:0] io_master_state_e_6_sreg_ss2,
  output [63:0] io_master_state_e_6_sreg_ss3,
  output [3:0]  io_master_state_e_6_base_vp_id,
  output        io_master_state_e_6_base_vp_valid,
  output        io_master_state_e_6_base_vp_scalar,
  output        io_master_state_e_6_base_vp_pred,
  output [7:0]  io_master_state_e_6_base_vs1_id,
  output        io_master_state_e_6_base_vs1_valid,
  output        io_master_state_e_6_base_vs1_scalar,
  output        io_master_state_e_6_base_vs1_pred,
  output [1:0]  io_master_state_e_6_base_vs1_prec,
  output [7:0]  io_master_state_e_6_base_vs2_id,
  output        io_master_state_e_6_base_vs2_valid,
  output        io_master_state_e_6_base_vs2_scalar,
  output        io_master_state_e_6_base_vs2_pred,
  output [1:0]  io_master_state_e_6_base_vs2_prec,
  output [7:0]  io_master_state_e_6_base_vs3_id,
  output        io_master_state_e_6_base_vs3_valid,
  output        io_master_state_e_6_base_vs3_scalar,
  output        io_master_state_e_6_base_vs3_pred,
  output [1:0]  io_master_state_e_6_base_vs3_prec,
  output [7:0]  io_master_state_e_6_base_vd_id,
  output        io_master_state_e_6_base_vd_valid,
  output        io_master_state_e_6_base_vd_scalar,
  output        io_master_state_e_6_base_vd_pred,
  output [1:0]  io_master_state_e_6_base_vd_prec,
  output        io_master_state_e_6_rate,
  output        io_master_state_e_6_active_viu,
  output        io_master_state_e_6_active_vipu,
  output        io_master_state_e_6_active_vimu,
  output        io_master_state_e_6_active_vidu,
  output        io_master_state_e_6_active_vfmu,
  output        io_master_state_e_6_active_vfdu,
  output        io_master_state_e_6_active_vfcu,
  output        io_master_state_e_6_active_vfvu,
  output        io_master_state_e_6_active_vrpu,
  output        io_master_state_e_6_active_vrfu,
  output        io_master_state_e_6_active_vpu,
  output        io_master_state_e_6_active_vgu,
  output        io_master_state_e_6_active_vcu,
  output        io_master_state_e_6_active_vlu,
  output        io_master_state_e_6_active_vsu,
  output        io_master_state_e_6_active_vqu,
  output        io_master_state_e_6_raw_0,
  output        io_master_state_e_6_raw_1,
  output        io_master_state_e_6_raw_2,
  output        io_master_state_e_6_raw_3,
  output        io_master_state_e_6_raw_4,
  output        io_master_state_e_6_raw_5,
  output        io_master_state_e_6_raw_6,
  output        io_master_state_e_6_raw_7,
  output        io_master_state_e_6_war_0,
  output        io_master_state_e_6_war_1,
  output        io_master_state_e_6_war_2,
  output        io_master_state_e_6_war_3,
  output        io_master_state_e_6_war_4,
  output        io_master_state_e_6_war_5,
  output        io_master_state_e_6_war_6,
  output        io_master_state_e_6_war_7,
  output        io_master_state_e_6_waw_0,
  output        io_master_state_e_6_waw_1,
  output        io_master_state_e_6_waw_2,
  output        io_master_state_e_6_waw_3,
  output        io_master_state_e_6_waw_4,
  output        io_master_state_e_6_waw_5,
  output        io_master_state_e_6_waw_6,
  output        io_master_state_e_6_waw_7,
  output        io_master_state_e_6_last,
  output [1:0]  io_master_state_e_6_rports,
  output [3:0]  io_master_state_e_6_wport_sram,
  output [2:0]  io_master_state_e_6_wport_pred,
  output [9:0]  io_master_state_e_7_fn_union,
  output [63:0] io_master_state_e_7_sreg_ss1,
  output [63:0] io_master_state_e_7_sreg_ss2,
  output [63:0] io_master_state_e_7_sreg_ss3,
  output [3:0]  io_master_state_e_7_base_vp_id,
  output        io_master_state_e_7_base_vp_valid,
  output        io_master_state_e_7_base_vp_scalar,
  output        io_master_state_e_7_base_vp_pred,
  output [7:0]  io_master_state_e_7_base_vs1_id,
  output        io_master_state_e_7_base_vs1_valid,
  output        io_master_state_e_7_base_vs1_scalar,
  output        io_master_state_e_7_base_vs1_pred,
  output [1:0]  io_master_state_e_7_base_vs1_prec,
  output [7:0]  io_master_state_e_7_base_vs2_id,
  output        io_master_state_e_7_base_vs2_valid,
  output        io_master_state_e_7_base_vs2_scalar,
  output        io_master_state_e_7_base_vs2_pred,
  output [1:0]  io_master_state_e_7_base_vs2_prec,
  output [7:0]  io_master_state_e_7_base_vs3_id,
  output        io_master_state_e_7_base_vs3_valid,
  output        io_master_state_e_7_base_vs3_scalar,
  output        io_master_state_e_7_base_vs3_pred,
  output [1:0]  io_master_state_e_7_base_vs3_prec,
  output [7:0]  io_master_state_e_7_base_vd_id,
  output        io_master_state_e_7_base_vd_valid,
  output        io_master_state_e_7_base_vd_scalar,
  output        io_master_state_e_7_base_vd_pred,
  output [1:0]  io_master_state_e_7_base_vd_prec,
  output        io_master_state_e_7_rate,
  output        io_master_state_e_7_active_viu,
  output        io_master_state_e_7_active_vipu,
  output        io_master_state_e_7_active_vimu,
  output        io_master_state_e_7_active_vidu,
  output        io_master_state_e_7_active_vfmu,
  output        io_master_state_e_7_active_vfdu,
  output        io_master_state_e_7_active_vfcu,
  output        io_master_state_e_7_active_vfvu,
  output        io_master_state_e_7_active_vrpu,
  output        io_master_state_e_7_active_vrfu,
  output        io_master_state_e_7_active_vpu,
  output        io_master_state_e_7_active_vgu,
  output        io_master_state_e_7_active_vcu,
  output        io_master_state_e_7_active_vlu,
  output        io_master_state_e_7_active_vsu,
  output        io_master_state_e_7_active_vqu,
  output        io_master_state_e_7_raw_0,
  output        io_master_state_e_7_raw_1,
  output        io_master_state_e_7_raw_2,
  output        io_master_state_e_7_raw_3,
  output        io_master_state_e_7_raw_4,
  output        io_master_state_e_7_raw_5,
  output        io_master_state_e_7_raw_6,
  output        io_master_state_e_7_raw_7,
  output        io_master_state_e_7_war_0,
  output        io_master_state_e_7_war_1,
  output        io_master_state_e_7_war_2,
  output        io_master_state_e_7_war_3,
  output        io_master_state_e_7_war_4,
  output        io_master_state_e_7_war_5,
  output        io_master_state_e_7_war_6,
  output        io_master_state_e_7_war_7,
  output        io_master_state_e_7_waw_0,
  output        io_master_state_e_7_waw_1,
  output        io_master_state_e_7_waw_2,
  output        io_master_state_e_7_waw_3,
  output        io_master_state_e_7_waw_4,
  output        io_master_state_e_7_waw_5,
  output        io_master_state_e_7_waw_6,
  output        io_master_state_e_7_waw_7,
  output        io_master_state_e_7_last,
  output [1:0]  io_master_state_e_7_rports,
  output [3:0]  io_master_state_e_7_wport_sram,
  output [2:0]  io_master_state_e_7_wport_pred,
  output [2:0]  io_master_state_head,
  output        io_master_update_valid_0,
  output        io_master_update_valid_1,
  output        io_master_update_valid_2,
  output        io_master_update_valid_3,
  output        io_master_update_valid_4,
  output        io_master_update_valid_5,
  output        io_master_update_valid_6,
  output        io_master_update_valid_7,
  output [7:0]  io_master_update_reg_0_vp_id,
  output [7:0]  io_master_update_reg_0_vs1_id,
  output [7:0]  io_master_update_reg_0_vs2_id,
  output [7:0]  io_master_update_reg_0_vs3_id,
  output [7:0]  io_master_update_reg_0_vd_id,
  output [7:0]  io_master_update_reg_1_vp_id,
  output [7:0]  io_master_update_reg_1_vs1_id,
  output [7:0]  io_master_update_reg_1_vs2_id,
  output [7:0]  io_master_update_reg_1_vs3_id,
  output [7:0]  io_master_update_reg_1_vd_id,
  output [7:0]  io_master_update_reg_2_vp_id,
  output [7:0]  io_master_update_reg_2_vs1_id,
  output [7:0]  io_master_update_reg_2_vs2_id,
  output [7:0]  io_master_update_reg_2_vs3_id,
  output [7:0]  io_master_update_reg_2_vd_id,
  output [7:0]  io_master_update_reg_3_vp_id,
  output [7:0]  io_master_update_reg_3_vs1_id,
  output [7:0]  io_master_update_reg_3_vs2_id,
  output [7:0]  io_master_update_reg_3_vs3_id,
  output [7:0]  io_master_update_reg_3_vd_id,
  output [7:0]  io_master_update_reg_4_vp_id,
  output [7:0]  io_master_update_reg_4_vs1_id,
  output [7:0]  io_master_update_reg_4_vs2_id,
  output [7:0]  io_master_update_reg_4_vs3_id,
  output [7:0]  io_master_update_reg_4_vd_id,
  output [7:0]  io_master_update_reg_5_vp_id,
  output [7:0]  io_master_update_reg_5_vs1_id,
  output [7:0]  io_master_update_reg_5_vs2_id,
  output [7:0]  io_master_update_reg_5_vs3_id,
  output [7:0]  io_master_update_reg_5_vd_id,
  output [7:0]  io_master_update_reg_6_vp_id,
  output [7:0]  io_master_update_reg_6_vs1_id,
  output [7:0]  io_master_update_reg_6_vs2_id,
  output [7:0]  io_master_update_reg_6_vs3_id,
  output [7:0]  io_master_update_reg_6_vd_id,
  output [7:0]  io_master_update_reg_7_vp_id,
  output [7:0]  io_master_update_reg_7_vs1_id,
  output [7:0]  io_master_update_reg_7_vs2_id,
  output [7:0]  io_master_update_reg_7_vs3_id,
  output [7:0]  io_master_update_reg_7_vd_id,
  input         io_master_clear_0,
  input         io_master_clear_1,
  input         io_master_clear_2,
  input         io_master_clear_3,
  input         io_master_clear_4,
  input         io_master_clear_5,
  input         io_master_clear_6,
  input         io_master_clear_7,
  output        io_pending_mem,
  output        io_pending_all,
  input         io_vf_stop,
  output        io_vf_last,
  output [2:0]  io_counters_memoryUOps,
  output [2:0]  io_counters_arithUOps,
  output [2:0]  io_counters_predUOps,
  output [2:0]  io_debug_head,
  output [2:0]  io_debug_tail,
  output        io_debug_maybe_full,
  output [3:0]  io_debug_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [63:0] _RAND_289;
  reg [63:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [63:0] _RAND_359;
  reg [63:0] _RAND_360;
  reg [63:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [63:0] _RAND_429;
  reg [63:0] _RAND_430;
  reg [63:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [63:0] _RAND_499;
  reg [63:0] _RAND_500;
  reg [63:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
`endif // RANDOMIZE_REG_INIT
  reg  v_0; // @[sequencer-master.scala 107:14]
  reg  v_1; // @[sequencer-master.scala 107:14]
  reg  v_2; // @[sequencer-master.scala 107:14]
  reg  v_3; // @[sequencer-master.scala 107:14]
  reg  v_4; // @[sequencer-master.scala 107:14]
  reg  v_5; // @[sequencer-master.scala 107:14]
  reg  v_6; // @[sequencer-master.scala 107:14]
  reg  v_7; // @[sequencer-master.scala 107:14]
  reg [9:0] e_0_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_0_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_0_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_0_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_0_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_0_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_0_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_0_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_0_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_0_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_0_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_0_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_0_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_0_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_0_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_0_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_0_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_0_war_0; // @[sequencer-master.scala 109:14]
  reg  e_0_war_1; // @[sequencer-master.scala 109:14]
  reg  e_0_war_2; // @[sequencer-master.scala 109:14]
  reg  e_0_war_3; // @[sequencer-master.scala 109:14]
  reg  e_0_war_4; // @[sequencer-master.scala 109:14]
  reg  e_0_war_5; // @[sequencer-master.scala 109:14]
  reg  e_0_war_6; // @[sequencer-master.scala 109:14]
  reg  e_0_war_7; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_0_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_0_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_0_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_0_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_0_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_1_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_1_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_1_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_1_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_1_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_1_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_1_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_1_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_1_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_1_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_1_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_1_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_1_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_1_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_1_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_1_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_1_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_1_war_0; // @[sequencer-master.scala 109:14]
  reg  e_1_war_1; // @[sequencer-master.scala 109:14]
  reg  e_1_war_2; // @[sequencer-master.scala 109:14]
  reg  e_1_war_3; // @[sequencer-master.scala 109:14]
  reg  e_1_war_4; // @[sequencer-master.scala 109:14]
  reg  e_1_war_5; // @[sequencer-master.scala 109:14]
  reg  e_1_war_6; // @[sequencer-master.scala 109:14]
  reg  e_1_war_7; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_1_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_1_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_1_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_1_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_1_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_2_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_2_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_2_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_2_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_2_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_2_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_2_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_2_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_2_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_2_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_2_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_2_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_2_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_2_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_2_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_2_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_2_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_2_war_0; // @[sequencer-master.scala 109:14]
  reg  e_2_war_1; // @[sequencer-master.scala 109:14]
  reg  e_2_war_2; // @[sequencer-master.scala 109:14]
  reg  e_2_war_3; // @[sequencer-master.scala 109:14]
  reg  e_2_war_4; // @[sequencer-master.scala 109:14]
  reg  e_2_war_5; // @[sequencer-master.scala 109:14]
  reg  e_2_war_6; // @[sequencer-master.scala 109:14]
  reg  e_2_war_7; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_2_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_2_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_2_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_2_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_2_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_3_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_3_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_3_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_3_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_3_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_3_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_3_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_3_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_3_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_3_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_3_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_3_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_3_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_3_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_3_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_3_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_3_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_3_war_0; // @[sequencer-master.scala 109:14]
  reg  e_3_war_1; // @[sequencer-master.scala 109:14]
  reg  e_3_war_2; // @[sequencer-master.scala 109:14]
  reg  e_3_war_3; // @[sequencer-master.scala 109:14]
  reg  e_3_war_4; // @[sequencer-master.scala 109:14]
  reg  e_3_war_5; // @[sequencer-master.scala 109:14]
  reg  e_3_war_6; // @[sequencer-master.scala 109:14]
  reg  e_3_war_7; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_3_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_3_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_3_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_3_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_3_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_4_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_4_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_4_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_4_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_4_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_4_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_4_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_4_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_4_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_4_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_4_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_4_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_4_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_4_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_4_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_4_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_4_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_4_war_0; // @[sequencer-master.scala 109:14]
  reg  e_4_war_1; // @[sequencer-master.scala 109:14]
  reg  e_4_war_2; // @[sequencer-master.scala 109:14]
  reg  e_4_war_3; // @[sequencer-master.scala 109:14]
  reg  e_4_war_4; // @[sequencer-master.scala 109:14]
  reg  e_4_war_5; // @[sequencer-master.scala 109:14]
  reg  e_4_war_6; // @[sequencer-master.scala 109:14]
  reg  e_4_war_7; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_4_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_4_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_4_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_4_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_4_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_5_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_5_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_5_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_5_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_5_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_5_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_5_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_5_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_5_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_5_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_5_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_5_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_5_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_5_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_5_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_5_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_5_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_5_war_0; // @[sequencer-master.scala 109:14]
  reg  e_5_war_1; // @[sequencer-master.scala 109:14]
  reg  e_5_war_2; // @[sequencer-master.scala 109:14]
  reg  e_5_war_3; // @[sequencer-master.scala 109:14]
  reg  e_5_war_4; // @[sequencer-master.scala 109:14]
  reg  e_5_war_5; // @[sequencer-master.scala 109:14]
  reg  e_5_war_6; // @[sequencer-master.scala 109:14]
  reg  e_5_war_7; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_5_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_5_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_5_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_5_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_5_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_6_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_6_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_6_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_6_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_6_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_6_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_6_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_6_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_6_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_6_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_6_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_6_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_6_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_6_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_6_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_6_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_6_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_6_war_0; // @[sequencer-master.scala 109:14]
  reg  e_6_war_1; // @[sequencer-master.scala 109:14]
  reg  e_6_war_2; // @[sequencer-master.scala 109:14]
  reg  e_6_war_3; // @[sequencer-master.scala 109:14]
  reg  e_6_war_4; // @[sequencer-master.scala 109:14]
  reg  e_6_war_5; // @[sequencer-master.scala 109:14]
  reg  e_6_war_6; // @[sequencer-master.scala 109:14]
  reg  e_6_war_7; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_6_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_6_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_6_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_6_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_6_wport_pred; // @[sequencer-master.scala 109:14]
  reg [9:0] e_7_fn_union; // @[sequencer-master.scala 109:14]
  reg [63:0] e_7_sreg_ss1; // @[sequencer-master.scala 109:14]
  reg [63:0] e_7_sreg_ss2; // @[sequencer-master.scala 109:14]
  reg [63:0] e_7_sreg_ss3; // @[sequencer-master.scala 109:14]
  reg [3:0] e_7_base_vp_id; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vp_valid; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vp_scalar; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vp_pred; // @[sequencer-master.scala 109:14]
  reg [7:0] e_7_base_vs1_id; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs1_valid; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs1_scalar; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs1_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_7_base_vs1_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_7_base_vs2_id; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs2_valid; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs2_scalar; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs2_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_7_base_vs2_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_7_base_vs3_id; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs3_valid; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs3_scalar; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vs3_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_7_base_vs3_prec; // @[sequencer-master.scala 109:14]
  reg [7:0] e_7_base_vd_id; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vd_valid; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vd_scalar; // @[sequencer-master.scala 109:14]
  reg  e_7_base_vd_pred; // @[sequencer-master.scala 109:14]
  reg [1:0] e_7_base_vd_prec; // @[sequencer-master.scala 109:14]
  reg  e_7_active_viu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vipu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vimu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vidu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vfmu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vfdu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vfcu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vfvu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vpu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vgu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vcu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vlu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vsu; // @[sequencer-master.scala 109:14]
  reg  e_7_active_vqu; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_0; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_1; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_2; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_3; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_4; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_5; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_6; // @[sequencer-master.scala 109:14]
  reg  e_7_raw_7; // @[sequencer-master.scala 109:14]
  reg  e_7_war_0; // @[sequencer-master.scala 109:14]
  reg  e_7_war_1; // @[sequencer-master.scala 109:14]
  reg  e_7_war_2; // @[sequencer-master.scala 109:14]
  reg  e_7_war_3; // @[sequencer-master.scala 109:14]
  reg  e_7_war_4; // @[sequencer-master.scala 109:14]
  reg  e_7_war_5; // @[sequencer-master.scala 109:14]
  reg  e_7_war_6; // @[sequencer-master.scala 109:14]
  reg  e_7_war_7; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_0; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_1; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_2; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_3; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_4; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_5; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_6; // @[sequencer-master.scala 109:14]
  reg  e_7_waw_7; // @[sequencer-master.scala 109:14]
  reg  e_7_last; // @[sequencer-master.scala 109:14]
  reg [1:0] e_7_rports; // @[sequencer-master.scala 109:14]
  reg [3:0] e_7_wport_sram; // @[sequencer-master.scala 109:14]
  reg [2:0] e_7_wport_pred; // @[sequencer-master.scala 109:14]
  reg  maybe_full; // @[sequencer-master.scala 111:23]
  reg [2:0] head; // @[sequencer-master.scala 112:17]
  reg [2:0] tail; // @[sequencer-master.scala 113:17]
  wire  _T_5 = v_0 & e_0_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_8 = ~e_0_base_vd_pred & e_0_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_9 = ~_T_8; // @[sequencer-master.scala 138:11]
  wire  _T_10 = _T_5 & io_op_bits_base_vp_valid & _T_9; // @[sequencer-master.scala 137:62]
  wire  _T_12 = ~io_op_bits_base_vp_pred & io_op_bits_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_22 = e_0_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_23 = ~(e_0_base_vd_pred | e_0_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_22; // @[sequencer-master.scala 139:75]
  wire  _T_24 = _T_10 & ~_T_12 & _T_23; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32712 = {{4'd0}, io_op_bits_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_25 = e_0_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_26 = _T_24 & _T_25; // @[sequencer-master.scala 140:72]
  wire  _T_27 = v_1 & e_1_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_30 = ~e_1_base_vd_pred & e_1_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_31 = ~_T_30; // @[sequencer-master.scala 138:11]
  wire  _T_32 = _T_27 & io_op_bits_base_vp_valid & _T_31; // @[sequencer-master.scala 137:62]
  wire  _T_44 = e_1_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_45 = ~(e_1_base_vd_pred | e_1_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_44; // @[sequencer-master.scala 139:75]
  wire  _T_46 = _T_32 & ~_T_12 & _T_45; // @[sequencer-master.scala 138:76]
  wire  _T_47 = e_1_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_48 = _T_46 & _T_47; // @[sequencer-master.scala 140:72]
  wire  _T_49 = v_2 & e_2_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_52 = ~e_2_base_vd_pred & e_2_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_53 = ~_T_52; // @[sequencer-master.scala 138:11]
  wire  _T_54 = _T_49 & io_op_bits_base_vp_valid & _T_53; // @[sequencer-master.scala 137:62]
  wire  _T_66 = e_2_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_67 = ~(e_2_base_vd_pred | e_2_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_66; // @[sequencer-master.scala 139:75]
  wire  _T_68 = _T_54 & ~_T_12 & _T_67; // @[sequencer-master.scala 138:76]
  wire  _T_69 = e_2_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_70 = _T_68 & _T_69; // @[sequencer-master.scala 140:72]
  wire  _T_71 = v_3 & e_3_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_74 = ~e_3_base_vd_pred & e_3_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_75 = ~_T_74; // @[sequencer-master.scala 138:11]
  wire  _T_76 = _T_71 & io_op_bits_base_vp_valid & _T_75; // @[sequencer-master.scala 137:62]
  wire  _T_88 = e_3_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_89 = ~(e_3_base_vd_pred | e_3_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_88; // @[sequencer-master.scala 139:75]
  wire  _T_90 = _T_76 & ~_T_12 & _T_89; // @[sequencer-master.scala 138:76]
  wire  _T_91 = e_3_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_92 = _T_90 & _T_91; // @[sequencer-master.scala 140:72]
  wire  _T_93 = v_4 & e_4_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_96 = ~e_4_base_vd_pred & e_4_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_97 = ~_T_96; // @[sequencer-master.scala 138:11]
  wire  _T_98 = _T_93 & io_op_bits_base_vp_valid & _T_97; // @[sequencer-master.scala 137:62]
  wire  _T_110 = e_4_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_111 = ~(e_4_base_vd_pred | e_4_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_110; // @[sequencer-master.scala 139:75]
  wire  _T_112 = _T_98 & ~_T_12 & _T_111; // @[sequencer-master.scala 138:76]
  wire  _T_113 = e_4_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_114 = _T_112 & _T_113; // @[sequencer-master.scala 140:72]
  wire  _T_115 = v_5 & e_5_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_118 = ~e_5_base_vd_pred & e_5_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_119 = ~_T_118; // @[sequencer-master.scala 138:11]
  wire  _T_120 = _T_115 & io_op_bits_base_vp_valid & _T_119; // @[sequencer-master.scala 137:62]
  wire  _T_132 = e_5_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_133 = ~(e_5_base_vd_pred | e_5_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_132; // @[sequencer-master.scala 139:75]
  wire  _T_134 = _T_120 & ~_T_12 & _T_133; // @[sequencer-master.scala 138:76]
  wire  _T_135 = e_5_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_136 = _T_134 & _T_135; // @[sequencer-master.scala 140:72]
  wire  _T_137 = v_6 & e_6_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_140 = ~e_6_base_vd_pred & e_6_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_141 = ~_T_140; // @[sequencer-master.scala 138:11]
  wire  _T_142 = _T_137 & io_op_bits_base_vp_valid & _T_141; // @[sequencer-master.scala 137:62]
  wire  _T_154 = e_6_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_155 = ~(e_6_base_vd_pred | e_6_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_154; // @[sequencer-master.scala 139:75]
  wire  _T_156 = _T_142 & ~_T_12 & _T_155; // @[sequencer-master.scala 138:76]
  wire  _T_157 = e_6_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_158 = _T_156 & _T_157; // @[sequencer-master.scala 140:72]
  wire  _T_159 = v_7 & e_7_base_vd_valid; // @[sequencer-master.scala 136:44]
  wire  _T_162 = ~e_7_base_vd_pred & e_7_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_163 = ~_T_162; // @[sequencer-master.scala 138:11]
  wire  _T_164 = _T_159 & io_op_bits_base_vp_valid & _T_163; // @[sequencer-master.scala 137:62]
  wire  _T_176 = e_7_base_vd_pred & io_op_bits_base_vp_pred; // @[sequencer-master.scala 140:37]
  wire  _T_177 = ~(e_7_base_vd_pred | e_7_base_vd_scalar) & ~(io_op_bits_base_vp_pred | io_op_bits_base_vp_scalar) |
    _T_176; // @[sequencer-master.scala 139:75]
  wire  _T_178 = _T_164 & ~_T_12 & _T_177; // @[sequencer-master.scala 138:76]
  wire  _T_179 = e_7_base_vd_id == _GEN_32712; // @[sequencer-master.scala 141:29]
  wire  _T_180 = _T_178 & _T_179; // @[sequencer-master.scala 140:72]
  wire  _T_187 = _T_5 & io_op_bits_base_vs1_valid & _T_9; // @[sequencer-master.scala 137:62]
  wire  _T_189 = ~io_op_bits_base_vs1_pred & io_op_bits_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_199 = e_0_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_200 = ~(e_0_base_vd_pred | e_0_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_199; // @[sequencer-master.scala 139:75]
  wire  _T_201 = _T_187 & ~_T_189 & _T_200; // @[sequencer-master.scala 138:76]
  wire  _T_202 = e_0_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_203 = _T_201 & _T_202; // @[sequencer-master.scala 140:72]
  wire  _T_209 = _T_27 & io_op_bits_base_vs1_valid & _T_31; // @[sequencer-master.scala 137:62]
  wire  _T_221 = e_1_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_222 = ~(e_1_base_vd_pred | e_1_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_221; // @[sequencer-master.scala 139:75]
  wire  _T_223 = _T_209 & ~_T_189 & _T_222; // @[sequencer-master.scala 138:76]
  wire  _T_224 = e_1_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_225 = _T_223 & _T_224; // @[sequencer-master.scala 140:72]
  wire  _T_231 = _T_49 & io_op_bits_base_vs1_valid & _T_53; // @[sequencer-master.scala 137:62]
  wire  _T_243 = e_2_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_244 = ~(e_2_base_vd_pred | e_2_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_243; // @[sequencer-master.scala 139:75]
  wire  _T_245 = _T_231 & ~_T_189 & _T_244; // @[sequencer-master.scala 138:76]
  wire  _T_246 = e_2_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_247 = _T_245 & _T_246; // @[sequencer-master.scala 140:72]
  wire  _T_253 = _T_71 & io_op_bits_base_vs1_valid & _T_75; // @[sequencer-master.scala 137:62]
  wire  _T_265 = e_3_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_266 = ~(e_3_base_vd_pred | e_3_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_265; // @[sequencer-master.scala 139:75]
  wire  _T_267 = _T_253 & ~_T_189 & _T_266; // @[sequencer-master.scala 138:76]
  wire  _T_268 = e_3_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_269 = _T_267 & _T_268; // @[sequencer-master.scala 140:72]
  wire  _T_275 = _T_93 & io_op_bits_base_vs1_valid & _T_97; // @[sequencer-master.scala 137:62]
  wire  _T_287 = e_4_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_288 = ~(e_4_base_vd_pred | e_4_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_287; // @[sequencer-master.scala 139:75]
  wire  _T_289 = _T_275 & ~_T_189 & _T_288; // @[sequencer-master.scala 138:76]
  wire  _T_290 = e_4_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_291 = _T_289 & _T_290; // @[sequencer-master.scala 140:72]
  wire  _T_297 = _T_115 & io_op_bits_base_vs1_valid & _T_119; // @[sequencer-master.scala 137:62]
  wire  _T_309 = e_5_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_310 = ~(e_5_base_vd_pred | e_5_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_309; // @[sequencer-master.scala 139:75]
  wire  _T_311 = _T_297 & ~_T_189 & _T_310; // @[sequencer-master.scala 138:76]
  wire  _T_312 = e_5_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_313 = _T_311 & _T_312; // @[sequencer-master.scala 140:72]
  wire  _T_319 = _T_137 & io_op_bits_base_vs1_valid & _T_141; // @[sequencer-master.scala 137:62]
  wire  _T_331 = e_6_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_332 = ~(e_6_base_vd_pred | e_6_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_331; // @[sequencer-master.scala 139:75]
  wire  _T_333 = _T_319 & ~_T_189 & _T_332; // @[sequencer-master.scala 138:76]
  wire  _T_334 = e_6_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_335 = _T_333 & _T_334; // @[sequencer-master.scala 140:72]
  wire  _T_341 = _T_159 & io_op_bits_base_vs1_valid & _T_163; // @[sequencer-master.scala 137:62]
  wire  _T_353 = e_7_base_vd_pred & io_op_bits_base_vs1_pred; // @[sequencer-master.scala 140:37]
  wire  _T_354 = ~(e_7_base_vd_pred | e_7_base_vd_scalar) & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar) |
    _T_353; // @[sequencer-master.scala 139:75]
  wire  _T_355 = _T_341 & ~_T_189 & _T_354; // @[sequencer-master.scala 138:76]
  wire  _T_356 = e_7_base_vd_id == io_op_bits_base_vs1_id; // @[sequencer-master.scala 141:29]
  wire  _T_357 = _T_355 & _T_356; // @[sequencer-master.scala 140:72]
  wire  _T_364 = _T_5 & io_op_bits_base_vs2_valid & _T_9; // @[sequencer-master.scala 137:62]
  wire  _T_366 = ~io_op_bits_base_vs2_pred & io_op_bits_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_376 = e_0_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_377 = ~(e_0_base_vd_pred | e_0_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_376; // @[sequencer-master.scala 139:75]
  wire  _T_378 = _T_364 & ~_T_366 & _T_377; // @[sequencer-master.scala 138:76]
  wire  _T_379 = e_0_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_380 = _T_378 & _T_379; // @[sequencer-master.scala 140:72]
  wire  _T_386 = _T_27 & io_op_bits_base_vs2_valid & _T_31; // @[sequencer-master.scala 137:62]
  wire  _T_398 = e_1_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_399 = ~(e_1_base_vd_pred | e_1_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_398; // @[sequencer-master.scala 139:75]
  wire  _T_400 = _T_386 & ~_T_366 & _T_399; // @[sequencer-master.scala 138:76]
  wire  _T_401 = e_1_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_402 = _T_400 & _T_401; // @[sequencer-master.scala 140:72]
  wire  _T_408 = _T_49 & io_op_bits_base_vs2_valid & _T_53; // @[sequencer-master.scala 137:62]
  wire  _T_420 = e_2_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_421 = ~(e_2_base_vd_pred | e_2_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_420; // @[sequencer-master.scala 139:75]
  wire  _T_422 = _T_408 & ~_T_366 & _T_421; // @[sequencer-master.scala 138:76]
  wire  _T_423 = e_2_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_424 = _T_422 & _T_423; // @[sequencer-master.scala 140:72]
  wire  _T_430 = _T_71 & io_op_bits_base_vs2_valid & _T_75; // @[sequencer-master.scala 137:62]
  wire  _T_442 = e_3_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_443 = ~(e_3_base_vd_pred | e_3_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_442; // @[sequencer-master.scala 139:75]
  wire  _T_444 = _T_430 & ~_T_366 & _T_443; // @[sequencer-master.scala 138:76]
  wire  _T_445 = e_3_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_446 = _T_444 & _T_445; // @[sequencer-master.scala 140:72]
  wire  _T_452 = _T_93 & io_op_bits_base_vs2_valid & _T_97; // @[sequencer-master.scala 137:62]
  wire  _T_464 = e_4_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_465 = ~(e_4_base_vd_pred | e_4_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_464; // @[sequencer-master.scala 139:75]
  wire  _T_466 = _T_452 & ~_T_366 & _T_465; // @[sequencer-master.scala 138:76]
  wire  _T_467 = e_4_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_468 = _T_466 & _T_467; // @[sequencer-master.scala 140:72]
  wire  _T_474 = _T_115 & io_op_bits_base_vs2_valid & _T_119; // @[sequencer-master.scala 137:62]
  wire  _T_486 = e_5_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_487 = ~(e_5_base_vd_pred | e_5_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_486; // @[sequencer-master.scala 139:75]
  wire  _T_488 = _T_474 & ~_T_366 & _T_487; // @[sequencer-master.scala 138:76]
  wire  _T_489 = e_5_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_490 = _T_488 & _T_489; // @[sequencer-master.scala 140:72]
  wire  _T_496 = _T_137 & io_op_bits_base_vs2_valid & _T_141; // @[sequencer-master.scala 137:62]
  wire  _T_508 = e_6_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_509 = ~(e_6_base_vd_pred | e_6_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_508; // @[sequencer-master.scala 139:75]
  wire  _T_510 = _T_496 & ~_T_366 & _T_509; // @[sequencer-master.scala 138:76]
  wire  _T_511 = e_6_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_512 = _T_510 & _T_511; // @[sequencer-master.scala 140:72]
  wire  _T_518 = _T_159 & io_op_bits_base_vs2_valid & _T_163; // @[sequencer-master.scala 137:62]
  wire  _T_530 = e_7_base_vd_pred & io_op_bits_base_vs2_pred; // @[sequencer-master.scala 140:37]
  wire  _T_531 = ~(e_7_base_vd_pred | e_7_base_vd_scalar) & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar) |
    _T_530; // @[sequencer-master.scala 139:75]
  wire  _T_532 = _T_518 & ~_T_366 & _T_531; // @[sequencer-master.scala 138:76]
  wire  _T_533 = e_7_base_vd_id == io_op_bits_base_vs2_id; // @[sequencer-master.scala 141:29]
  wire  _T_534 = _T_532 & _T_533; // @[sequencer-master.scala 140:72]
  wire  _T_541 = _T_5 & io_op_bits_base_vs3_valid & _T_9; // @[sequencer-master.scala 137:62]
  wire  _T_543 = ~io_op_bits_base_vs3_pred & io_op_bits_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_553 = e_0_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_554 = ~(e_0_base_vd_pred | e_0_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_553; // @[sequencer-master.scala 139:75]
  wire  _T_555 = _T_541 & ~_T_543 & _T_554; // @[sequencer-master.scala 138:76]
  wire  _T_556 = e_0_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_557 = _T_555 & _T_556; // @[sequencer-master.scala 140:72]
  wire  _T_563 = _T_27 & io_op_bits_base_vs3_valid & _T_31; // @[sequencer-master.scala 137:62]
  wire  _T_575 = e_1_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_576 = ~(e_1_base_vd_pred | e_1_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_575; // @[sequencer-master.scala 139:75]
  wire  _T_577 = _T_563 & ~_T_543 & _T_576; // @[sequencer-master.scala 138:76]
  wire  _T_578 = e_1_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_579 = _T_577 & _T_578; // @[sequencer-master.scala 140:72]
  wire  _T_585 = _T_49 & io_op_bits_base_vs3_valid & _T_53; // @[sequencer-master.scala 137:62]
  wire  _T_597 = e_2_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_598 = ~(e_2_base_vd_pred | e_2_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_597; // @[sequencer-master.scala 139:75]
  wire  _T_599 = _T_585 & ~_T_543 & _T_598; // @[sequencer-master.scala 138:76]
  wire  _T_600 = e_2_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_601 = _T_599 & _T_600; // @[sequencer-master.scala 140:72]
  wire  _T_607 = _T_71 & io_op_bits_base_vs3_valid & _T_75; // @[sequencer-master.scala 137:62]
  wire  _T_619 = e_3_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_620 = ~(e_3_base_vd_pred | e_3_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_619; // @[sequencer-master.scala 139:75]
  wire  _T_621 = _T_607 & ~_T_543 & _T_620; // @[sequencer-master.scala 138:76]
  wire  _T_622 = e_3_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_623 = _T_621 & _T_622; // @[sequencer-master.scala 140:72]
  wire  _T_629 = _T_93 & io_op_bits_base_vs3_valid & _T_97; // @[sequencer-master.scala 137:62]
  wire  _T_641 = e_4_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_642 = ~(e_4_base_vd_pred | e_4_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_641; // @[sequencer-master.scala 139:75]
  wire  _T_643 = _T_629 & ~_T_543 & _T_642; // @[sequencer-master.scala 138:76]
  wire  _T_644 = e_4_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_645 = _T_643 & _T_644; // @[sequencer-master.scala 140:72]
  wire  _T_651 = _T_115 & io_op_bits_base_vs3_valid & _T_119; // @[sequencer-master.scala 137:62]
  wire  _T_663 = e_5_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_664 = ~(e_5_base_vd_pred | e_5_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_663; // @[sequencer-master.scala 139:75]
  wire  _T_665 = _T_651 & ~_T_543 & _T_664; // @[sequencer-master.scala 138:76]
  wire  _T_666 = e_5_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_667 = _T_665 & _T_666; // @[sequencer-master.scala 140:72]
  wire  _T_673 = _T_137 & io_op_bits_base_vs3_valid & _T_141; // @[sequencer-master.scala 137:62]
  wire  _T_685 = e_6_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_686 = ~(e_6_base_vd_pred | e_6_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_685; // @[sequencer-master.scala 139:75]
  wire  _T_687 = _T_673 & ~_T_543 & _T_686; // @[sequencer-master.scala 138:76]
  wire  _T_688 = e_6_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_689 = _T_687 & _T_688; // @[sequencer-master.scala 140:72]
  wire  _T_695 = _T_159 & io_op_bits_base_vs3_valid & _T_163; // @[sequencer-master.scala 137:62]
  wire  _T_707 = e_7_base_vd_pred & io_op_bits_base_vs3_pred; // @[sequencer-master.scala 140:37]
  wire  _T_708 = ~(e_7_base_vd_pred | e_7_base_vd_scalar) & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar) |
    _T_707; // @[sequencer-master.scala 139:75]
  wire  _T_709 = _T_695 & ~_T_543 & _T_708; // @[sequencer-master.scala 138:76]
  wire  _T_710 = e_7_base_vd_id == io_op_bits_base_vs3_id; // @[sequencer-master.scala 141:29]
  wire  _T_711 = _T_709 & _T_710; // @[sequencer-master.scala 140:72]
  wire  _T_713 = v_0 & e_0_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_716 = ~e_0_base_vp_pred & e_0_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_717 = ~_T_716; // @[sequencer-master.scala 138:11]
  wire  _T_718 = _T_713 & io_op_bits_base_vd_valid & _T_717; // @[sequencer-master.scala 137:62]
  wire  _T_720 = ~io_op_bits_base_vd_pred & io_op_bits_base_vd_scalar; // @[types-vxu.scala 119:37]
  wire  _T_721 = ~_T_720; // @[sequencer-master.scala 138:42]
  wire  _T_730 = e_0_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_731 = ~(e_0_base_vp_pred | e_0_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_730; // @[sequencer-master.scala 139:75]
  wire  _T_732 = _T_718 & ~_T_720 & _T_731; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32720 = {{4'd0}, e_0_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_733 = _GEN_32720 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_734 = _T_732 & _T_733; // @[sequencer-master.scala 140:72]
  wire  _T_735 = v_1 & e_1_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_738 = ~e_1_base_vp_pred & e_1_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_739 = ~_T_738; // @[sequencer-master.scala 138:11]
  wire  _T_740 = _T_735 & io_op_bits_base_vd_valid & _T_739; // @[sequencer-master.scala 137:62]
  wire  _T_752 = e_1_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_753 = ~(e_1_base_vp_pred | e_1_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_752; // @[sequencer-master.scala 139:75]
  wire  _T_754 = _T_740 & ~_T_720 & _T_753; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32721 = {{4'd0}, e_1_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_755 = _GEN_32721 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_756 = _T_754 & _T_755; // @[sequencer-master.scala 140:72]
  wire  _T_757 = v_2 & e_2_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_760 = ~e_2_base_vp_pred & e_2_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_761 = ~_T_760; // @[sequencer-master.scala 138:11]
  wire  _T_762 = _T_757 & io_op_bits_base_vd_valid & _T_761; // @[sequencer-master.scala 137:62]
  wire  _T_774 = e_2_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_775 = ~(e_2_base_vp_pred | e_2_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_774; // @[sequencer-master.scala 139:75]
  wire  _T_776 = _T_762 & ~_T_720 & _T_775; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32722 = {{4'd0}, e_2_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_777 = _GEN_32722 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_778 = _T_776 & _T_777; // @[sequencer-master.scala 140:72]
  wire  _T_779 = v_3 & e_3_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_782 = ~e_3_base_vp_pred & e_3_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_783 = ~_T_782; // @[sequencer-master.scala 138:11]
  wire  _T_784 = _T_779 & io_op_bits_base_vd_valid & _T_783; // @[sequencer-master.scala 137:62]
  wire  _T_796 = e_3_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_797 = ~(e_3_base_vp_pred | e_3_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_796; // @[sequencer-master.scala 139:75]
  wire  _T_798 = _T_784 & ~_T_720 & _T_797; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32723 = {{4'd0}, e_3_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_799 = _GEN_32723 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_800 = _T_798 & _T_799; // @[sequencer-master.scala 140:72]
  wire  _T_801 = v_4 & e_4_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_804 = ~e_4_base_vp_pred & e_4_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_805 = ~_T_804; // @[sequencer-master.scala 138:11]
  wire  _T_806 = _T_801 & io_op_bits_base_vd_valid & _T_805; // @[sequencer-master.scala 137:62]
  wire  _T_818 = e_4_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_819 = ~(e_4_base_vp_pred | e_4_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_818; // @[sequencer-master.scala 139:75]
  wire  _T_820 = _T_806 & ~_T_720 & _T_819; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32724 = {{4'd0}, e_4_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_821 = _GEN_32724 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_822 = _T_820 & _T_821; // @[sequencer-master.scala 140:72]
  wire  _T_823 = v_5 & e_5_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_826 = ~e_5_base_vp_pred & e_5_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_827 = ~_T_826; // @[sequencer-master.scala 138:11]
  wire  _T_828 = _T_823 & io_op_bits_base_vd_valid & _T_827; // @[sequencer-master.scala 137:62]
  wire  _T_840 = e_5_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_841 = ~(e_5_base_vp_pred | e_5_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_840; // @[sequencer-master.scala 139:75]
  wire  _T_842 = _T_828 & ~_T_720 & _T_841; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32725 = {{4'd0}, e_5_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_843 = _GEN_32725 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_844 = _T_842 & _T_843; // @[sequencer-master.scala 140:72]
  wire  _T_845 = v_6 & e_6_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_848 = ~e_6_base_vp_pred & e_6_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_849 = ~_T_848; // @[sequencer-master.scala 138:11]
  wire  _T_850 = _T_845 & io_op_bits_base_vd_valid & _T_849; // @[sequencer-master.scala 137:62]
  wire  _T_862 = e_6_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_863 = ~(e_6_base_vp_pred | e_6_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_862; // @[sequencer-master.scala 139:75]
  wire  _T_864 = _T_850 & ~_T_720 & _T_863; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32726 = {{4'd0}, e_6_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_865 = _GEN_32726 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_866 = _T_864 & _T_865; // @[sequencer-master.scala 140:72]
  wire  _T_867 = v_7 & e_7_base_vp_valid; // @[sequencer-master.scala 136:44]
  wire  _T_870 = ~e_7_base_vp_pred & e_7_base_vp_scalar; // @[types-vxu.scala 119:37]
  wire  _T_871 = ~_T_870; // @[sequencer-master.scala 138:11]
  wire  _T_872 = _T_867 & io_op_bits_base_vd_valid & _T_871; // @[sequencer-master.scala 137:62]
  wire  _T_884 = e_7_base_vp_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_885 = ~(e_7_base_vp_pred | e_7_base_vp_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_884; // @[sequencer-master.scala 139:75]
  wire  _T_886 = _T_872 & ~_T_720 & _T_885; // @[sequencer-master.scala 138:76]
  wire [7:0] _GEN_32727 = {{4'd0}, e_7_base_vp_id}; // @[sequencer-master.scala 141:29]
  wire  _T_887 = _GEN_32727 == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_888 = _T_886 & _T_887; // @[sequencer-master.scala 140:72]
  wire  _T_890 = v_0 & e_0_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_893 = ~e_0_base_vs1_pred & e_0_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_894 = ~_T_893; // @[sequencer-master.scala 138:11]
  wire  _T_895 = _T_890 & io_op_bits_base_vd_valid & _T_894; // @[sequencer-master.scala 137:62]
  wire  _T_907 = e_0_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_908 = ~(e_0_base_vs1_pred | e_0_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_907; // @[sequencer-master.scala 139:75]
  wire  _T_909 = _T_895 & ~_T_720 & _T_908; // @[sequencer-master.scala 138:76]
  wire  _T_910 = e_0_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_911 = _T_909 & _T_910; // @[sequencer-master.scala 140:72]
  wire  _T_912 = v_1 & e_1_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_915 = ~e_1_base_vs1_pred & e_1_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_916 = ~_T_915; // @[sequencer-master.scala 138:11]
  wire  _T_917 = _T_912 & io_op_bits_base_vd_valid & _T_916; // @[sequencer-master.scala 137:62]
  wire  _T_929 = e_1_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_930 = ~(e_1_base_vs1_pred | e_1_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_929; // @[sequencer-master.scala 139:75]
  wire  _T_931 = _T_917 & ~_T_720 & _T_930; // @[sequencer-master.scala 138:76]
  wire  _T_932 = e_1_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_933 = _T_931 & _T_932; // @[sequencer-master.scala 140:72]
  wire  _T_934 = v_2 & e_2_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_937 = ~e_2_base_vs1_pred & e_2_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_938 = ~_T_937; // @[sequencer-master.scala 138:11]
  wire  _T_939 = _T_934 & io_op_bits_base_vd_valid & _T_938; // @[sequencer-master.scala 137:62]
  wire  _T_951 = e_2_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_952 = ~(e_2_base_vs1_pred | e_2_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_951; // @[sequencer-master.scala 139:75]
  wire  _T_953 = _T_939 & ~_T_720 & _T_952; // @[sequencer-master.scala 138:76]
  wire  _T_954 = e_2_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_955 = _T_953 & _T_954; // @[sequencer-master.scala 140:72]
  wire  _T_956 = v_3 & e_3_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_959 = ~e_3_base_vs1_pred & e_3_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_960 = ~_T_959; // @[sequencer-master.scala 138:11]
  wire  _T_961 = _T_956 & io_op_bits_base_vd_valid & _T_960; // @[sequencer-master.scala 137:62]
  wire  _T_973 = e_3_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_974 = ~(e_3_base_vs1_pred | e_3_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_973; // @[sequencer-master.scala 139:75]
  wire  _T_975 = _T_961 & ~_T_720 & _T_974; // @[sequencer-master.scala 138:76]
  wire  _T_976 = e_3_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_977 = _T_975 & _T_976; // @[sequencer-master.scala 140:72]
  wire  _T_978 = v_4 & e_4_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_981 = ~e_4_base_vs1_pred & e_4_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_982 = ~_T_981; // @[sequencer-master.scala 138:11]
  wire  _T_983 = _T_978 & io_op_bits_base_vd_valid & _T_982; // @[sequencer-master.scala 137:62]
  wire  _T_995 = e_4_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_996 = ~(e_4_base_vs1_pred | e_4_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_995; // @[sequencer-master.scala 139:75]
  wire  _T_997 = _T_983 & ~_T_720 & _T_996; // @[sequencer-master.scala 138:76]
  wire  _T_998 = e_4_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_999 = _T_997 & _T_998; // @[sequencer-master.scala 140:72]
  wire  _T_1000 = v_5 & e_5_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1003 = ~e_5_base_vs1_pred & e_5_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1004 = ~_T_1003; // @[sequencer-master.scala 138:11]
  wire  _T_1005 = _T_1000 & io_op_bits_base_vd_valid & _T_1004; // @[sequencer-master.scala 137:62]
  wire  _T_1017 = e_5_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1018 = ~(e_5_base_vs1_pred | e_5_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1017; // @[sequencer-master.scala 139:75]
  wire  _T_1019 = _T_1005 & ~_T_720 & _T_1018; // @[sequencer-master.scala 138:76]
  wire  _T_1020 = e_5_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1021 = _T_1019 & _T_1020; // @[sequencer-master.scala 140:72]
  wire  _T_1022 = v_6 & e_6_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1025 = ~e_6_base_vs1_pred & e_6_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1026 = ~_T_1025; // @[sequencer-master.scala 138:11]
  wire  _T_1027 = _T_1022 & io_op_bits_base_vd_valid & _T_1026; // @[sequencer-master.scala 137:62]
  wire  _T_1039 = e_6_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1040 = ~(e_6_base_vs1_pred | e_6_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1039; // @[sequencer-master.scala 139:75]
  wire  _T_1041 = _T_1027 & ~_T_720 & _T_1040; // @[sequencer-master.scala 138:76]
  wire  _T_1042 = e_6_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1043 = _T_1041 & _T_1042; // @[sequencer-master.scala 140:72]
  wire  _T_1044 = v_7 & e_7_base_vs1_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1047 = ~e_7_base_vs1_pred & e_7_base_vs1_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1048 = ~_T_1047; // @[sequencer-master.scala 138:11]
  wire  _T_1049 = _T_1044 & io_op_bits_base_vd_valid & _T_1048; // @[sequencer-master.scala 137:62]
  wire  _T_1061 = e_7_base_vs1_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1062 = ~(e_7_base_vs1_pred | e_7_base_vs1_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1061; // @[sequencer-master.scala 139:75]
  wire  _T_1063 = _T_1049 & ~_T_720 & _T_1062; // @[sequencer-master.scala 138:76]
  wire  _T_1064 = e_7_base_vs1_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1065 = _T_1063 & _T_1064; // @[sequencer-master.scala 140:72]
  wire  _T_1067 = v_0 & e_0_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1070 = ~e_0_base_vs2_pred & e_0_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1071 = ~_T_1070; // @[sequencer-master.scala 138:11]
  wire  _T_1072 = _T_1067 & io_op_bits_base_vd_valid & _T_1071; // @[sequencer-master.scala 137:62]
  wire  _T_1084 = e_0_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1085 = ~(e_0_base_vs2_pred | e_0_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1084; // @[sequencer-master.scala 139:75]
  wire  _T_1086 = _T_1072 & ~_T_720 & _T_1085; // @[sequencer-master.scala 138:76]
  wire  _T_1087 = e_0_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1088 = _T_1086 & _T_1087; // @[sequencer-master.scala 140:72]
  wire  _T_1089 = v_1 & e_1_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1092 = ~e_1_base_vs2_pred & e_1_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1093 = ~_T_1092; // @[sequencer-master.scala 138:11]
  wire  _T_1094 = _T_1089 & io_op_bits_base_vd_valid & _T_1093; // @[sequencer-master.scala 137:62]
  wire  _T_1106 = e_1_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1107 = ~(e_1_base_vs2_pred | e_1_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1106; // @[sequencer-master.scala 139:75]
  wire  _T_1108 = _T_1094 & ~_T_720 & _T_1107; // @[sequencer-master.scala 138:76]
  wire  _T_1109 = e_1_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1110 = _T_1108 & _T_1109; // @[sequencer-master.scala 140:72]
  wire  _T_1111 = v_2 & e_2_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1114 = ~e_2_base_vs2_pred & e_2_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1115 = ~_T_1114; // @[sequencer-master.scala 138:11]
  wire  _T_1116 = _T_1111 & io_op_bits_base_vd_valid & _T_1115; // @[sequencer-master.scala 137:62]
  wire  _T_1128 = e_2_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1129 = ~(e_2_base_vs2_pred | e_2_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1128; // @[sequencer-master.scala 139:75]
  wire  _T_1130 = _T_1116 & ~_T_720 & _T_1129; // @[sequencer-master.scala 138:76]
  wire  _T_1131 = e_2_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1132 = _T_1130 & _T_1131; // @[sequencer-master.scala 140:72]
  wire  _T_1133 = v_3 & e_3_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1136 = ~e_3_base_vs2_pred & e_3_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1137 = ~_T_1136; // @[sequencer-master.scala 138:11]
  wire  _T_1138 = _T_1133 & io_op_bits_base_vd_valid & _T_1137; // @[sequencer-master.scala 137:62]
  wire  _T_1150 = e_3_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1151 = ~(e_3_base_vs2_pred | e_3_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1150; // @[sequencer-master.scala 139:75]
  wire  _T_1152 = _T_1138 & ~_T_720 & _T_1151; // @[sequencer-master.scala 138:76]
  wire  _T_1153 = e_3_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1154 = _T_1152 & _T_1153; // @[sequencer-master.scala 140:72]
  wire  _T_1155 = v_4 & e_4_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1158 = ~e_4_base_vs2_pred & e_4_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1159 = ~_T_1158; // @[sequencer-master.scala 138:11]
  wire  _T_1160 = _T_1155 & io_op_bits_base_vd_valid & _T_1159; // @[sequencer-master.scala 137:62]
  wire  _T_1172 = e_4_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1173 = ~(e_4_base_vs2_pred | e_4_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1172; // @[sequencer-master.scala 139:75]
  wire  _T_1174 = _T_1160 & ~_T_720 & _T_1173; // @[sequencer-master.scala 138:76]
  wire  _T_1175 = e_4_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1176 = _T_1174 & _T_1175; // @[sequencer-master.scala 140:72]
  wire  _T_1177 = v_5 & e_5_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1180 = ~e_5_base_vs2_pred & e_5_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1181 = ~_T_1180; // @[sequencer-master.scala 138:11]
  wire  _T_1182 = _T_1177 & io_op_bits_base_vd_valid & _T_1181; // @[sequencer-master.scala 137:62]
  wire  _T_1194 = e_5_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1195 = ~(e_5_base_vs2_pred | e_5_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1194; // @[sequencer-master.scala 139:75]
  wire  _T_1196 = _T_1182 & ~_T_720 & _T_1195; // @[sequencer-master.scala 138:76]
  wire  _T_1197 = e_5_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1198 = _T_1196 & _T_1197; // @[sequencer-master.scala 140:72]
  wire  _T_1199 = v_6 & e_6_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1202 = ~e_6_base_vs2_pred & e_6_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1203 = ~_T_1202; // @[sequencer-master.scala 138:11]
  wire  _T_1204 = _T_1199 & io_op_bits_base_vd_valid & _T_1203; // @[sequencer-master.scala 137:62]
  wire  _T_1216 = e_6_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1217 = ~(e_6_base_vs2_pred | e_6_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1216; // @[sequencer-master.scala 139:75]
  wire  _T_1218 = _T_1204 & ~_T_720 & _T_1217; // @[sequencer-master.scala 138:76]
  wire  _T_1219 = e_6_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1220 = _T_1218 & _T_1219; // @[sequencer-master.scala 140:72]
  wire  _T_1221 = v_7 & e_7_base_vs2_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1224 = ~e_7_base_vs2_pred & e_7_base_vs2_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1225 = ~_T_1224; // @[sequencer-master.scala 138:11]
  wire  _T_1226 = _T_1221 & io_op_bits_base_vd_valid & _T_1225; // @[sequencer-master.scala 137:62]
  wire  _T_1238 = e_7_base_vs2_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1239 = ~(e_7_base_vs2_pred | e_7_base_vs2_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1238; // @[sequencer-master.scala 139:75]
  wire  _T_1240 = _T_1226 & ~_T_720 & _T_1239; // @[sequencer-master.scala 138:76]
  wire  _T_1241 = e_7_base_vs2_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1242 = _T_1240 & _T_1241; // @[sequencer-master.scala 140:72]
  wire  _T_1244 = v_0 & e_0_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1247 = ~e_0_base_vs3_pred & e_0_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1248 = ~_T_1247; // @[sequencer-master.scala 138:11]
  wire  _T_1249 = _T_1244 & io_op_bits_base_vd_valid & _T_1248; // @[sequencer-master.scala 137:62]
  wire  _T_1261 = e_0_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1262 = ~(e_0_base_vs3_pred | e_0_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1261; // @[sequencer-master.scala 139:75]
  wire  _T_1263 = _T_1249 & ~_T_720 & _T_1262; // @[sequencer-master.scala 138:76]
  wire  _T_1264 = e_0_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1265 = _T_1263 & _T_1264; // @[sequencer-master.scala 140:72]
  wire  _T_1266 = v_1 & e_1_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1269 = ~e_1_base_vs3_pred & e_1_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1270 = ~_T_1269; // @[sequencer-master.scala 138:11]
  wire  _T_1271 = _T_1266 & io_op_bits_base_vd_valid & _T_1270; // @[sequencer-master.scala 137:62]
  wire  _T_1283 = e_1_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1284 = ~(e_1_base_vs3_pred | e_1_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1283; // @[sequencer-master.scala 139:75]
  wire  _T_1285 = _T_1271 & ~_T_720 & _T_1284; // @[sequencer-master.scala 138:76]
  wire  _T_1286 = e_1_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1287 = _T_1285 & _T_1286; // @[sequencer-master.scala 140:72]
  wire  _T_1288 = v_2 & e_2_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1291 = ~e_2_base_vs3_pred & e_2_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1292 = ~_T_1291; // @[sequencer-master.scala 138:11]
  wire  _T_1293 = _T_1288 & io_op_bits_base_vd_valid & _T_1292; // @[sequencer-master.scala 137:62]
  wire  _T_1305 = e_2_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1306 = ~(e_2_base_vs3_pred | e_2_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1305; // @[sequencer-master.scala 139:75]
  wire  _T_1307 = _T_1293 & ~_T_720 & _T_1306; // @[sequencer-master.scala 138:76]
  wire  _T_1308 = e_2_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1309 = _T_1307 & _T_1308; // @[sequencer-master.scala 140:72]
  wire  _T_1310 = v_3 & e_3_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1313 = ~e_3_base_vs3_pred & e_3_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1314 = ~_T_1313; // @[sequencer-master.scala 138:11]
  wire  _T_1315 = _T_1310 & io_op_bits_base_vd_valid & _T_1314; // @[sequencer-master.scala 137:62]
  wire  _T_1327 = e_3_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1328 = ~(e_3_base_vs3_pred | e_3_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1327; // @[sequencer-master.scala 139:75]
  wire  _T_1329 = _T_1315 & ~_T_720 & _T_1328; // @[sequencer-master.scala 138:76]
  wire  _T_1330 = e_3_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1331 = _T_1329 & _T_1330; // @[sequencer-master.scala 140:72]
  wire  _T_1332 = v_4 & e_4_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1335 = ~e_4_base_vs3_pred & e_4_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1336 = ~_T_1335; // @[sequencer-master.scala 138:11]
  wire  _T_1337 = _T_1332 & io_op_bits_base_vd_valid & _T_1336; // @[sequencer-master.scala 137:62]
  wire  _T_1349 = e_4_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1350 = ~(e_4_base_vs3_pred | e_4_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1349; // @[sequencer-master.scala 139:75]
  wire  _T_1351 = _T_1337 & ~_T_720 & _T_1350; // @[sequencer-master.scala 138:76]
  wire  _T_1352 = e_4_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1353 = _T_1351 & _T_1352; // @[sequencer-master.scala 140:72]
  wire  _T_1354 = v_5 & e_5_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1357 = ~e_5_base_vs3_pred & e_5_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1358 = ~_T_1357; // @[sequencer-master.scala 138:11]
  wire  _T_1359 = _T_1354 & io_op_bits_base_vd_valid & _T_1358; // @[sequencer-master.scala 137:62]
  wire  _T_1371 = e_5_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1372 = ~(e_5_base_vs3_pred | e_5_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1371; // @[sequencer-master.scala 139:75]
  wire  _T_1373 = _T_1359 & ~_T_720 & _T_1372; // @[sequencer-master.scala 138:76]
  wire  _T_1374 = e_5_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1375 = _T_1373 & _T_1374; // @[sequencer-master.scala 140:72]
  wire  _T_1376 = v_6 & e_6_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1379 = ~e_6_base_vs3_pred & e_6_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1380 = ~_T_1379; // @[sequencer-master.scala 138:11]
  wire  _T_1381 = _T_1376 & io_op_bits_base_vd_valid & _T_1380; // @[sequencer-master.scala 137:62]
  wire  _T_1393 = e_6_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1394 = ~(e_6_base_vs3_pred | e_6_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1393; // @[sequencer-master.scala 139:75]
  wire  _T_1395 = _T_1381 & ~_T_720 & _T_1394; // @[sequencer-master.scala 138:76]
  wire  _T_1396 = e_6_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1397 = _T_1395 & _T_1396; // @[sequencer-master.scala 140:72]
  wire  _T_1398 = v_7 & e_7_base_vs3_valid; // @[sequencer-master.scala 136:44]
  wire  _T_1401 = ~e_7_base_vs3_pred & e_7_base_vs3_scalar; // @[types-vxu.scala 119:37]
  wire  _T_1402 = ~_T_1401; // @[sequencer-master.scala 138:11]
  wire  _T_1403 = _T_1398 & io_op_bits_base_vd_valid & _T_1402; // @[sequencer-master.scala 137:62]
  wire  _T_1415 = e_7_base_vs3_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1416 = ~(e_7_base_vs3_pred | e_7_base_vs3_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1415; // @[sequencer-master.scala 139:75]
  wire  _T_1417 = _T_1403 & ~_T_720 & _T_1416; // @[sequencer-master.scala 138:76]
  wire  _T_1418 = e_7_base_vs3_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1419 = _T_1417 & _T_1418; // @[sequencer-master.scala 140:72]
  wire  _T_1426 = _T_5 & io_op_bits_base_vd_valid & _T_9; // @[sequencer-master.scala 137:62]
  wire  _T_1438 = e_0_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1439 = ~(e_0_base_vd_pred | e_0_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1438; // @[sequencer-master.scala 139:75]
  wire  _T_1440 = _T_1426 & ~_T_720 & _T_1439; // @[sequencer-master.scala 138:76]
  wire  _T_1441 = e_0_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1442 = _T_1440 & _T_1441; // @[sequencer-master.scala 140:72]
  wire  _T_1448 = _T_27 & io_op_bits_base_vd_valid & _T_31; // @[sequencer-master.scala 137:62]
  wire  _T_1460 = e_1_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1461 = ~(e_1_base_vd_pred | e_1_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1460; // @[sequencer-master.scala 139:75]
  wire  _T_1462 = _T_1448 & ~_T_720 & _T_1461; // @[sequencer-master.scala 138:76]
  wire  _T_1463 = e_1_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1464 = _T_1462 & _T_1463; // @[sequencer-master.scala 140:72]
  wire  _T_1470 = _T_49 & io_op_bits_base_vd_valid & _T_53; // @[sequencer-master.scala 137:62]
  wire  _T_1482 = e_2_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1483 = ~(e_2_base_vd_pred | e_2_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1482; // @[sequencer-master.scala 139:75]
  wire  _T_1484 = _T_1470 & ~_T_720 & _T_1483; // @[sequencer-master.scala 138:76]
  wire  _T_1485 = e_2_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1486 = _T_1484 & _T_1485; // @[sequencer-master.scala 140:72]
  wire  _T_1492 = _T_71 & io_op_bits_base_vd_valid & _T_75; // @[sequencer-master.scala 137:62]
  wire  _T_1504 = e_3_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1505 = ~(e_3_base_vd_pred | e_3_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1504; // @[sequencer-master.scala 139:75]
  wire  _T_1506 = _T_1492 & ~_T_720 & _T_1505; // @[sequencer-master.scala 138:76]
  wire  _T_1507 = e_3_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1508 = _T_1506 & _T_1507; // @[sequencer-master.scala 140:72]
  wire  _T_1514 = _T_93 & io_op_bits_base_vd_valid & _T_97; // @[sequencer-master.scala 137:62]
  wire  _T_1526 = e_4_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1527 = ~(e_4_base_vd_pred | e_4_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1526; // @[sequencer-master.scala 139:75]
  wire  _T_1528 = _T_1514 & ~_T_720 & _T_1527; // @[sequencer-master.scala 138:76]
  wire  _T_1529 = e_4_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1530 = _T_1528 & _T_1529; // @[sequencer-master.scala 140:72]
  wire  _T_1536 = _T_115 & io_op_bits_base_vd_valid & _T_119; // @[sequencer-master.scala 137:62]
  wire  _T_1548 = e_5_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1549 = ~(e_5_base_vd_pred | e_5_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1548; // @[sequencer-master.scala 139:75]
  wire  _T_1550 = _T_1536 & ~_T_720 & _T_1549; // @[sequencer-master.scala 138:76]
  wire  _T_1551 = e_5_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1552 = _T_1550 & _T_1551; // @[sequencer-master.scala 140:72]
  wire  _T_1558 = _T_137 & io_op_bits_base_vd_valid & _T_141; // @[sequencer-master.scala 137:62]
  wire  _T_1570 = e_6_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1571 = ~(e_6_base_vd_pred | e_6_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1570; // @[sequencer-master.scala 139:75]
  wire  _T_1572 = _T_1558 & ~_T_720 & _T_1571; // @[sequencer-master.scala 138:76]
  wire  _T_1573 = e_6_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1574 = _T_1572 & _T_1573; // @[sequencer-master.scala 140:72]
  wire  _T_1580 = _T_159 & io_op_bits_base_vd_valid & _T_163; // @[sequencer-master.scala 137:62]
  wire  _T_1592 = e_7_base_vd_pred & io_op_bits_base_vd_pred; // @[sequencer-master.scala 140:37]
  wire  _T_1593 = ~(e_7_base_vd_pred | e_7_base_vd_scalar) & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) |
    _T_1592; // @[sequencer-master.scala 139:75]
  wire  _T_1594 = _T_1580 & ~_T_720 & _T_1593; // @[sequencer-master.scala 138:76]
  wire  _T_1595 = e_7_base_vd_id == io_op_bits_base_vd_id; // @[sequencer-master.scala 141:29]
  wire  _T_1596 = _T_1594 & _T_1595; // @[sequencer-master.scala 140:72]
  wire  _T_1601 = io_op_bits_base_vs1_valid & ~(io_op_bits_base_vs1_pred | io_op_bits_base_vs1_scalar); // @[sequencer-master.scala 218:69]
  wire  _T_1605 = io_op_bits_base_vs2_valid & ~(io_op_bits_base_vs2_pred | io_op_bits_base_vs2_scalar); // @[sequencer-master.scala 218:69]
  wire  _T_1609 = io_op_bits_base_vs3_valid & ~(io_op_bits_base_vs3_pred | io_op_bits_base_vs3_scalar); // @[sequencer-master.scala 218:69]
  wire [1:0] _T_1610 = _T_1605 + _T_1609; // @[Bitwise.scala 48:55]
  wire [1:0] _GEN_32728 = {{1'd0}, _T_1601}; // @[Bitwise.scala 48:55]
  wire [2:0] _T_1611 = _GEN_32728 + _T_1610; // @[Bitwise.scala 48:55]
  wire  _T_1612 = ~io_op_bits_active_vipred; // @[sequencer-master.scala 220:21]
  wire [2:0] _T_1615 = _T_1611 > 3'h0 ? _T_1611 : {{2'd0}, _T_1612}; // @[sequencer-master.scala 222:12]
  wire  _T_1623 = _T_1601 > 1'h0 ? _T_1601 : _T_1612; // @[sequencer-master.scala 222:12]
  wire  _T_1631 = _T_1605 > 1'h0 ? _T_1605 : _T_1612; // @[sequencer-master.scala 222:12]
  wire  _T_1635 = io_op_bits_base_vd_valid & ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar); // @[sequencer-master.scala 218:69]
  wire  _T_1639 = _T_1635 > 1'h0 ? _T_1635 : _T_1612; // @[sequencer-master.scala 222:12]
  wire [2:0] _T_1645 = tail + 3'h1; // @[util.scala 94:11]
  wire [2:0] _T_1647 = tail + 3'h2; // @[util.scala 94:11]
  wire [2:0] _T_1649 = tail + 3'h3; // @[util.scala 94:11]
  wire [2:0] _T_1651 = tail + 3'h4; // @[util.scala 94:11]
  wire  _T_1752 = io_op_ready & io_op_valid; // @[Decoupled.scala 37:37]
  wire  _GEN_32729 = 3'h0 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_0 = 3'h0 == tail | v_0; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32730 = 3'h1 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_1 = 3'h1 == tail | v_1; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32731 = 3'h2 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_2 = 3'h2 == tail | v_2; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32732 = 3'h3 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_3 = 3'h3 == tail | v_3; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32733 = 3'h4 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_4 = 3'h4 == tail | v_4; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32734 = 3'h5 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_5 = 3'h5 == tail | v_5; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32735 = 3'h6 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_6 = 3'h6 == tail | v_6; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_32736 = 3'h7 == tail; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_7 = 3'h7 == tail | v_7; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35 sequencer-master.scala 107:14]
  wire  _GEN_16 = 3'h0 == tail ? 1'h0 : e_0_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_17 = 3'h1 == tail ? 1'h0 : e_1_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_18 = 3'h2 == tail ? 1'h0 : e_2_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_19 = 3'h3 == tail ? 1'h0 : e_3_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_20 = 3'h4 == tail ? 1'h0 : e_4_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_21 = 3'h5 == tail ? 1'h0 : e_5_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_22 = 3'h6 == tail ? 1'h0 : e_6_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_23 = 3'h7 == tail ? 1'h0 : e_7_base_vp_valid; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28 sequencer-master.scala 109:14]
  wire  _GEN_24 = 3'h0 == tail ? 1'h0 : e_0_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_25 = 3'h1 == tail ? 1'h0 : e_1_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_26 = 3'h2 == tail ? 1'h0 : e_2_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_27 = 3'h3 == tail ? 1'h0 : e_3_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_28 = 3'h4 == tail ? 1'h0 : e_4_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_29 = 3'h5 == tail ? 1'h0 : e_5_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_30 = 3'h6 == tail ? 1'h0 : e_6_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_31 = 3'h7 == tail ? 1'h0 : e_7_base_vs1_valid; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29 sequencer-master.scala 109:14]
  wire  _GEN_32 = 3'h0 == tail ? 1'h0 : e_0_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_33 = 3'h1 == tail ? 1'h0 : e_1_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_34 = 3'h2 == tail ? 1'h0 : e_2_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_35 = 3'h3 == tail ? 1'h0 : e_3_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_36 = 3'h4 == tail ? 1'h0 : e_4_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_37 = 3'h5 == tail ? 1'h0 : e_5_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_38 = 3'h6 == tail ? 1'h0 : e_6_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_39 = 3'h7 == tail ? 1'h0 : e_7_base_vs2_valid; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29 sequencer-master.scala 109:14]
  wire  _GEN_40 = 3'h0 == tail ? 1'h0 : e_0_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_41 = 3'h1 == tail ? 1'h0 : e_1_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_42 = 3'h2 == tail ? 1'h0 : e_2_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_43 = 3'h3 == tail ? 1'h0 : e_3_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_44 = 3'h4 == tail ? 1'h0 : e_4_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_45 = 3'h5 == tail ? 1'h0 : e_5_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_46 = 3'h6 == tail ? 1'h0 : e_6_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_47 = 3'h7 == tail ? 1'h0 : e_7_base_vs3_valid; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29 sequencer-master.scala 109:14]
  wire  _GEN_48 = 3'h0 == tail ? 1'h0 : e_0_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_49 = 3'h1 == tail ? 1'h0 : e_1_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_50 = 3'h2 == tail ? 1'h0 : e_2_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_51 = 3'h3 == tail ? 1'h0 : e_3_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_52 = 3'h4 == tail ? 1'h0 : e_4_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_53 = 3'h5 == tail ? 1'h0 : e_5_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_54 = 3'h6 == tail ? 1'h0 : e_6_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_55 = 3'h7 == tail ? 1'h0 : e_7_base_vd_valid; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28 sequencer-master.scala 109:14]
  wire  _GEN_64 = 3'h0 == tail ? 1'h0 : e_0_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_65 = 3'h1 == tail ? 1'h0 : e_1_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_66 = 3'h2 == tail ? 1'h0 : e_2_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_67 = 3'h3 == tail ? 1'h0 : e_3_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_68 = 3'h4 == tail ? 1'h0 : e_4_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_69 = 3'h5 == tail ? 1'h0 : e_5_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_70 = 3'h6 == tail ? 1'h0 : e_6_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_71 = 3'h7 == tail ? 1'h0 : e_7_raw_0; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_72 = 3'h0 == tail ? 1'h0 : e_0_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_73 = 3'h1 == tail ? 1'h0 : e_1_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_74 = 3'h2 == tail ? 1'h0 : e_2_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_75 = 3'h3 == tail ? 1'h0 : e_3_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_76 = 3'h4 == tail ? 1'h0 : e_4_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_77 = 3'h5 == tail ? 1'h0 : e_5_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_78 = 3'h6 == tail ? 1'h0 : e_6_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_79 = 3'h7 == tail ? 1'h0 : e_7_war_0; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_80 = 3'h0 == tail ? 1'h0 : e_0_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_81 = 3'h1 == tail ? 1'h0 : e_1_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_82 = 3'h2 == tail ? 1'h0 : e_2_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_83 = 3'h3 == tail ? 1'h0 : e_3_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_84 = 3'h4 == tail ? 1'h0 : e_4_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_85 = 3'h5 == tail ? 1'h0 : e_5_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_86 = 3'h6 == tail ? 1'h0 : e_6_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_87 = 3'h7 == tail ? 1'h0 : e_7_waw_0; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_88 = 3'h0 == tail ? 1'h0 : e_0_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_89 = 3'h1 == tail ? 1'h0 : e_1_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_90 = 3'h2 == tail ? 1'h0 : e_2_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_91 = 3'h3 == tail ? 1'h0 : e_3_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_92 = 3'h4 == tail ? 1'h0 : e_4_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_93 = 3'h5 == tail ? 1'h0 : e_5_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_94 = 3'h6 == tail ? 1'h0 : e_6_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_95 = 3'h7 == tail ? 1'h0 : e_7_raw_1; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_96 = 3'h0 == tail ? 1'h0 : e_0_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_97 = 3'h1 == tail ? 1'h0 : e_1_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_98 = 3'h2 == tail ? 1'h0 : e_2_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_99 = 3'h3 == tail ? 1'h0 : e_3_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_100 = 3'h4 == tail ? 1'h0 : e_4_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_101 = 3'h5 == tail ? 1'h0 : e_5_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_102 = 3'h6 == tail ? 1'h0 : e_6_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_103 = 3'h7 == tail ? 1'h0 : e_7_war_1; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_104 = 3'h0 == tail ? 1'h0 : e_0_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_105 = 3'h1 == tail ? 1'h0 : e_1_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_106 = 3'h2 == tail ? 1'h0 : e_2_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_107 = 3'h3 == tail ? 1'h0 : e_3_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_108 = 3'h4 == tail ? 1'h0 : e_4_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_109 = 3'h5 == tail ? 1'h0 : e_5_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_110 = 3'h6 == tail ? 1'h0 : e_6_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_111 = 3'h7 == tail ? 1'h0 : e_7_waw_1; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_112 = 3'h0 == tail ? 1'h0 : e_0_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_113 = 3'h1 == tail ? 1'h0 : e_1_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_114 = 3'h2 == tail ? 1'h0 : e_2_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_115 = 3'h3 == tail ? 1'h0 : e_3_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_116 = 3'h4 == tail ? 1'h0 : e_4_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_117 = 3'h5 == tail ? 1'h0 : e_5_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_118 = 3'h6 == tail ? 1'h0 : e_6_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_119 = 3'h7 == tail ? 1'h0 : e_7_raw_2; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_120 = 3'h0 == tail ? 1'h0 : e_0_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_121 = 3'h1 == tail ? 1'h0 : e_1_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_122 = 3'h2 == tail ? 1'h0 : e_2_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_123 = 3'h3 == tail ? 1'h0 : e_3_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_124 = 3'h4 == tail ? 1'h0 : e_4_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_125 = 3'h5 == tail ? 1'h0 : e_5_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_126 = 3'h6 == tail ? 1'h0 : e_6_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_127 = 3'h7 == tail ? 1'h0 : e_7_war_2; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_128 = 3'h0 == tail ? 1'h0 : e_0_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_129 = 3'h1 == tail ? 1'h0 : e_1_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_130 = 3'h2 == tail ? 1'h0 : e_2_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_131 = 3'h3 == tail ? 1'h0 : e_3_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_132 = 3'h4 == tail ? 1'h0 : e_4_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_133 = 3'h5 == tail ? 1'h0 : e_5_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_134 = 3'h6 == tail ? 1'h0 : e_6_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_135 = 3'h7 == tail ? 1'h0 : e_7_waw_2; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_136 = 3'h0 == tail ? 1'h0 : e_0_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_137 = 3'h1 == tail ? 1'h0 : e_1_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_138 = 3'h2 == tail ? 1'h0 : e_2_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_139 = 3'h3 == tail ? 1'h0 : e_3_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_140 = 3'h4 == tail ? 1'h0 : e_4_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_141 = 3'h5 == tail ? 1'h0 : e_5_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_142 = 3'h6 == tail ? 1'h0 : e_6_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_143 = 3'h7 == tail ? 1'h0 : e_7_raw_3; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_144 = 3'h0 == tail ? 1'h0 : e_0_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_145 = 3'h1 == tail ? 1'h0 : e_1_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_146 = 3'h2 == tail ? 1'h0 : e_2_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_147 = 3'h3 == tail ? 1'h0 : e_3_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_148 = 3'h4 == tail ? 1'h0 : e_4_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_149 = 3'h5 == tail ? 1'h0 : e_5_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_150 = 3'h6 == tail ? 1'h0 : e_6_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_151 = 3'h7 == tail ? 1'h0 : e_7_war_3; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_152 = 3'h0 == tail ? 1'h0 : e_0_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_153 = 3'h1 == tail ? 1'h0 : e_1_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_154 = 3'h2 == tail ? 1'h0 : e_2_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_155 = 3'h3 == tail ? 1'h0 : e_3_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_156 = 3'h4 == tail ? 1'h0 : e_4_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_157 = 3'h5 == tail ? 1'h0 : e_5_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_158 = 3'h6 == tail ? 1'h0 : e_6_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_159 = 3'h7 == tail ? 1'h0 : e_7_waw_3; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_160 = 3'h0 == tail ? 1'h0 : e_0_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_161 = 3'h1 == tail ? 1'h0 : e_1_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_162 = 3'h2 == tail ? 1'h0 : e_2_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_163 = 3'h3 == tail ? 1'h0 : e_3_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_164 = 3'h4 == tail ? 1'h0 : e_4_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_165 = 3'h5 == tail ? 1'h0 : e_5_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_166 = 3'h6 == tail ? 1'h0 : e_6_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_167 = 3'h7 == tail ? 1'h0 : e_7_raw_4; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_168 = 3'h0 == tail ? 1'h0 : e_0_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_169 = 3'h1 == tail ? 1'h0 : e_1_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_170 = 3'h2 == tail ? 1'h0 : e_2_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_171 = 3'h3 == tail ? 1'h0 : e_3_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_172 = 3'h4 == tail ? 1'h0 : e_4_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_173 = 3'h5 == tail ? 1'h0 : e_5_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_174 = 3'h6 == tail ? 1'h0 : e_6_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_175 = 3'h7 == tail ? 1'h0 : e_7_war_4; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_176 = 3'h0 == tail ? 1'h0 : e_0_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_177 = 3'h1 == tail ? 1'h0 : e_1_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_178 = 3'h2 == tail ? 1'h0 : e_2_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_179 = 3'h3 == tail ? 1'h0 : e_3_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_180 = 3'h4 == tail ? 1'h0 : e_4_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_181 = 3'h5 == tail ? 1'h0 : e_5_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_182 = 3'h6 == tail ? 1'h0 : e_6_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_183 = 3'h7 == tail ? 1'h0 : e_7_waw_4; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_184 = 3'h0 == tail ? 1'h0 : e_0_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_185 = 3'h1 == tail ? 1'h0 : e_1_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_186 = 3'h2 == tail ? 1'h0 : e_2_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_187 = 3'h3 == tail ? 1'h0 : e_3_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_188 = 3'h4 == tail ? 1'h0 : e_4_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_189 = 3'h5 == tail ? 1'h0 : e_5_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_190 = 3'h6 == tail ? 1'h0 : e_6_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_191 = 3'h7 == tail ? 1'h0 : e_7_raw_5; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_192 = 3'h0 == tail ? 1'h0 : e_0_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_193 = 3'h1 == tail ? 1'h0 : e_1_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_194 = 3'h2 == tail ? 1'h0 : e_2_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_195 = 3'h3 == tail ? 1'h0 : e_3_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_196 = 3'h4 == tail ? 1'h0 : e_4_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_197 = 3'h5 == tail ? 1'h0 : e_5_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_198 = 3'h6 == tail ? 1'h0 : e_6_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_199 = 3'h7 == tail ? 1'h0 : e_7_war_5; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_200 = 3'h0 == tail ? 1'h0 : e_0_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_201 = 3'h1 == tail ? 1'h0 : e_1_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_202 = 3'h2 == tail ? 1'h0 : e_2_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_203 = 3'h3 == tail ? 1'h0 : e_3_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_204 = 3'h4 == tail ? 1'h0 : e_4_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_205 = 3'h5 == tail ? 1'h0 : e_5_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_206 = 3'h6 == tail ? 1'h0 : e_6_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_207 = 3'h7 == tail ? 1'h0 : e_7_waw_5; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_208 = 3'h0 == tail ? 1'h0 : e_0_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_209 = 3'h1 == tail ? 1'h0 : e_1_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_210 = 3'h2 == tail ? 1'h0 : e_2_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_211 = 3'h3 == tail ? 1'h0 : e_3_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_212 = 3'h4 == tail ? 1'h0 : e_4_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_213 = 3'h5 == tail ? 1'h0 : e_5_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_214 = 3'h6 == tail ? 1'h0 : e_6_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_215 = 3'h7 == tail ? 1'h0 : e_7_raw_6; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_216 = 3'h0 == tail ? 1'h0 : e_0_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_217 = 3'h1 == tail ? 1'h0 : e_1_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_218 = 3'h2 == tail ? 1'h0 : e_2_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_219 = 3'h3 == tail ? 1'h0 : e_3_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_220 = 3'h4 == tail ? 1'h0 : e_4_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_221 = 3'h5 == tail ? 1'h0 : e_5_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_222 = 3'h6 == tail ? 1'h0 : e_6_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_223 = 3'h7 == tail ? 1'h0 : e_7_war_6; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_224 = 3'h0 == tail ? 1'h0 : e_0_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_225 = 3'h1 == tail ? 1'h0 : e_1_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_226 = 3'h2 == tail ? 1'h0 : e_2_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_227 = 3'h3 == tail ? 1'h0 : e_3_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_228 = 3'h4 == tail ? 1'h0 : e_4_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_229 = 3'h5 == tail ? 1'h0 : e_5_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_230 = 3'h6 == tail ? 1'h0 : e_6_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_231 = 3'h7 == tail ? 1'h0 : e_7_waw_6; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_232 = 3'h0 == tail ? 1'h0 : e_0_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_233 = 3'h1 == tail ? 1'h0 : e_1_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_234 = 3'h2 == tail ? 1'h0 : e_2_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_235 = 3'h3 == tail ? 1'h0 : e_3_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_236 = 3'h4 == tail ? 1'h0 : e_4_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_237 = 3'h5 == tail ? 1'h0 : e_5_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_238 = 3'h6 == tail ? 1'h0 : e_6_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_239 = 3'h7 == tail ? 1'h0 : e_7_raw_7; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52 sequencer-master.scala 194:26]
  wire  _GEN_240 = 3'h0 == tail ? 1'h0 : e_0_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_241 = 3'h1 == tail ? 1'h0 : e_1_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_242 = 3'h2 == tail ? 1'h0 : e_2_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_243 = 3'h3 == tail ? 1'h0 : e_3_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_244 = 3'h4 == tail ? 1'h0 : e_4_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_245 = 3'h5 == tail ? 1'h0 : e_5_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_246 = 3'h6 == tail ? 1'h0 : e_6_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_247 = 3'h7 == tail ? 1'h0 : e_7_war_7; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52 sequencer-master.scala 195:26]
  wire  _GEN_248 = 3'h0 == tail ? 1'h0 : e_0_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_249 = 3'h1 == tail ? 1'h0 : e_1_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_250 = 3'h2 == tail ? 1'h0 : e_2_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_251 = 3'h3 == tail ? 1'h0 : e_3_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_252 = 3'h4 == tail ? 1'h0 : e_4_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_253 = 3'h5 == tail ? 1'h0 : e_5_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_254 = 3'h6 == tail ? 1'h0 : e_6_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_255 = 3'h7 == tail ? 1'h0 : e_7_waw_7; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52 sequencer-master.scala 196:26]
  wire  _GEN_256 = 3'h0 == tail ? 1'h0 : e_0_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_257 = 3'h1 == tail ? 1'h0 : e_1_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_258 = 3'h2 == tail ? 1'h0 : e_2_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_259 = 3'h3 == tail ? 1'h0 : e_3_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_260 = 3'h4 == tail ? 1'h0 : e_4_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_261 = 3'h5 == tail ? 1'h0 : e_5_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_262 = 3'h6 == tail ? 1'h0 : e_6_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_263 = 3'h7 == tail ? 1'h0 : e_7_last; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19 sequencer-master.scala 109:14]
  wire  _GEN_272 = _GEN_32729 | e_0_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_273 = _GEN_32730 | e_1_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_274 = _GEN_32731 | e_2_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_275 = _GEN_32732 | e_3_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_276 = _GEN_32733 | e_4_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_277 = _GEN_32734 | e_5_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_278 = _GEN_32735 | e_6_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_279 = _GEN_32736 | e_7_active_viu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_280 = 3'h0 == tail ? io_op_bits_fn_union : e_0_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_281 = 3'h1 == tail ? io_op_bits_fn_union : e_1_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_282 = 3'h2 == tail ? io_op_bits_fn_union : e_2_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_283 = 3'h3 == tail ? io_op_bits_fn_union : e_3_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_284 = 3'h4 == tail ? io_op_bits_fn_union : e_4_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_285 = 3'h5 == tail ? io_op_bits_fn_union : e_5_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_286 = 3'h6 == tail ? io_op_bits_fn_union : e_6_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [9:0] _GEN_287 = 3'h7 == tail ? io_op_bits_fn_union : e_7_fn_union; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23 sequencer-master.scala 109:14]
  wire [3:0] _GEN_288 = 3'h0 == tail ? io_op_bits_base_vp_id : e_0_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_289 = 3'h1 == tail ? io_op_bits_base_vp_id : e_1_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_290 = 3'h2 == tail ? io_op_bits_base_vp_id : e_2_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_291 = 3'h3 == tail ? io_op_bits_base_vp_id : e_3_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_292 = 3'h4 == tail ? io_op_bits_base_vp_id : e_4_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_293 = 3'h5 == tail ? io_op_bits_base_vp_id : e_5_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_294 = 3'h6 == tail ? io_op_bits_base_vp_id : e_6_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [3:0] _GEN_295 = 3'h7 == tail ? io_op_bits_base_vp_id : e_7_base_vp_id; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_296 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_16; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_297 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_17; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_298 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_18; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_299 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_19; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_300 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_20; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_301 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_21; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_302 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_22; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_303 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_23; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_304 = 3'h0 == tail ? io_op_bits_base_vp_scalar : e_0_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_305 = 3'h1 == tail ? io_op_bits_base_vp_scalar : e_1_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_306 = 3'h2 == tail ? io_op_bits_base_vp_scalar : e_2_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_307 = 3'h3 == tail ? io_op_bits_base_vp_scalar : e_3_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_308 = 3'h4 == tail ? io_op_bits_base_vp_scalar : e_4_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_309 = 3'h5 == tail ? io_op_bits_base_vp_scalar : e_5_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_310 = 3'h6 == tail ? io_op_bits_base_vp_scalar : e_6_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_311 = 3'h7 == tail ? io_op_bits_base_vp_scalar : e_7_base_vp_scalar; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_312 = 3'h0 == tail ? io_op_bits_base_vp_pred : e_0_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_313 = 3'h1 == tail ? io_op_bits_base_vp_pred : e_1_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_314 = 3'h2 == tail ? io_op_bits_base_vp_pred : e_2_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_315 = 3'h3 == tail ? io_op_bits_base_vp_pred : e_3_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_316 = 3'h4 == tail ? io_op_bits_base_vp_pred : e_4_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_317 = 3'h5 == tail ? io_op_bits_base_vp_pred : e_5_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_318 = 3'h6 == tail ? io_op_bits_base_vp_pred : e_6_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire  _GEN_319 = 3'h7 == tail ? io_op_bits_base_vp_pred : e_7_base_vp_pred; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_320 = 3'h0 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_321 = 3'h1 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_322 = 3'h2 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_323 = 3'h3 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_324 = 3'h4 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_325 = 3'h5 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_326 = 3'h6 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_327 = 3'h7 == tail ? io_op_bits_reg_vp_id : 8'h0; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41 sequencer-master.scala 411:33]
  wire [3:0] _GEN_328 = io_op_bits_base_vp_valid ? _GEN_288 : e_0_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_329 = io_op_bits_base_vp_valid ? _GEN_289 : e_1_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_330 = io_op_bits_base_vp_valid ? _GEN_290 : e_2_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_331 = io_op_bits_base_vp_valid ? _GEN_291 : e_3_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_332 = io_op_bits_base_vp_valid ? _GEN_292 : e_4_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_333 = io_op_bits_base_vp_valid ? _GEN_293 : e_5_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_334 = io_op_bits_base_vp_valid ? _GEN_294 : e_6_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [3:0] _GEN_335 = io_op_bits_base_vp_valid ? _GEN_295 : e_7_base_vp_id; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_336 = io_op_bits_base_vp_valid ? _GEN_296 : _GEN_16; // @[sequencer-master.scala 320:41]
  wire  _GEN_337 = io_op_bits_base_vp_valid ? _GEN_297 : _GEN_17; // @[sequencer-master.scala 320:41]
  wire  _GEN_338 = io_op_bits_base_vp_valid ? _GEN_298 : _GEN_18; // @[sequencer-master.scala 320:41]
  wire  _GEN_339 = io_op_bits_base_vp_valid ? _GEN_299 : _GEN_19; // @[sequencer-master.scala 320:41]
  wire  _GEN_340 = io_op_bits_base_vp_valid ? _GEN_300 : _GEN_20; // @[sequencer-master.scala 320:41]
  wire  _GEN_341 = io_op_bits_base_vp_valid ? _GEN_301 : _GEN_21; // @[sequencer-master.scala 320:41]
  wire  _GEN_342 = io_op_bits_base_vp_valid ? _GEN_302 : _GEN_22; // @[sequencer-master.scala 320:41]
  wire  _GEN_343 = io_op_bits_base_vp_valid ? _GEN_303 : _GEN_23; // @[sequencer-master.scala 320:41]
  wire  _GEN_344 = io_op_bits_base_vp_valid ? _GEN_304 : e_0_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_345 = io_op_bits_base_vp_valid ? _GEN_305 : e_1_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_346 = io_op_bits_base_vp_valid ? _GEN_306 : e_2_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_347 = io_op_bits_base_vp_valid ? _GEN_307 : e_3_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_348 = io_op_bits_base_vp_valid ? _GEN_308 : e_4_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_349 = io_op_bits_base_vp_valid ? _GEN_309 : e_5_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_350 = io_op_bits_base_vp_valid ? _GEN_310 : e_6_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_351 = io_op_bits_base_vp_valid ? _GEN_311 : e_7_base_vp_scalar; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_352 = io_op_bits_base_vp_valid ? _GEN_312 : e_0_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_353 = io_op_bits_base_vp_valid ? _GEN_313 : e_1_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_354 = io_op_bits_base_vp_valid ? _GEN_314 : e_2_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_355 = io_op_bits_base_vp_valid ? _GEN_315 : e_3_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_356 = io_op_bits_base_vp_valid ? _GEN_316 : e_4_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_357 = io_op_bits_base_vp_valid ? _GEN_317 : e_5_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_358 = io_op_bits_base_vp_valid ? _GEN_318 : e_6_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire  _GEN_359 = io_op_bits_base_vp_valid ? _GEN_319 : e_7_base_vp_pred; // @[sequencer-master.scala 320:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_360 = io_op_bits_base_vp_valid ? _GEN_320 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_361 = io_op_bits_base_vp_valid ? _GEN_321 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_362 = io_op_bits_base_vp_valid ? _GEN_322 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_363 = io_op_bits_base_vp_valid ? _GEN_323 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_364 = io_op_bits_base_vp_valid ? _GEN_324 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_365 = io_op_bits_base_vp_valid ? _GEN_325 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_366 = io_op_bits_base_vp_valid ? _GEN_326 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_367 = io_op_bits_base_vp_valid ? _GEN_327 : 8'h0; // @[sequencer-master.scala 320:41 sequencer-master.scala 411:33]
  wire  _GEN_368 = _GEN_32729 | _GEN_64; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_369 = _GEN_32730 | _GEN_65; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_370 = _GEN_32731 | _GEN_66; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_371 = _GEN_32732 | _GEN_67; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_372 = _GEN_32733 | _GEN_68; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_373 = _GEN_32734 | _GEN_69; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_374 = _GEN_32735 | _GEN_70; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_375 = _GEN_32736 | _GEN_71; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_376 = _T_26 ? _GEN_368 : _GEN_64; // @[sequencer-master.scala 154:24]
  wire  _GEN_377 = _T_26 ? _GEN_369 : _GEN_65; // @[sequencer-master.scala 154:24]
  wire  _GEN_378 = _T_26 ? _GEN_370 : _GEN_66; // @[sequencer-master.scala 154:24]
  wire  _GEN_379 = _T_26 ? _GEN_371 : _GEN_67; // @[sequencer-master.scala 154:24]
  wire  _GEN_380 = _T_26 ? _GEN_372 : _GEN_68; // @[sequencer-master.scala 154:24]
  wire  _GEN_381 = _T_26 ? _GEN_373 : _GEN_69; // @[sequencer-master.scala 154:24]
  wire  _GEN_382 = _T_26 ? _GEN_374 : _GEN_70; // @[sequencer-master.scala 154:24]
  wire  _GEN_383 = _T_26 ? _GEN_375 : _GEN_71; // @[sequencer-master.scala 154:24]
  wire  _GEN_384 = _GEN_32729 | _GEN_88; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_385 = _GEN_32730 | _GEN_89; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_386 = _GEN_32731 | _GEN_90; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_387 = _GEN_32732 | _GEN_91; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_388 = _GEN_32733 | _GEN_92; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_389 = _GEN_32734 | _GEN_93; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_390 = _GEN_32735 | _GEN_94; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_391 = _GEN_32736 | _GEN_95; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_392 = _T_48 ? _GEN_384 : _GEN_88; // @[sequencer-master.scala 154:24]
  wire  _GEN_393 = _T_48 ? _GEN_385 : _GEN_89; // @[sequencer-master.scala 154:24]
  wire  _GEN_394 = _T_48 ? _GEN_386 : _GEN_90; // @[sequencer-master.scala 154:24]
  wire  _GEN_395 = _T_48 ? _GEN_387 : _GEN_91; // @[sequencer-master.scala 154:24]
  wire  _GEN_396 = _T_48 ? _GEN_388 : _GEN_92; // @[sequencer-master.scala 154:24]
  wire  _GEN_397 = _T_48 ? _GEN_389 : _GEN_93; // @[sequencer-master.scala 154:24]
  wire  _GEN_398 = _T_48 ? _GEN_390 : _GEN_94; // @[sequencer-master.scala 154:24]
  wire  _GEN_399 = _T_48 ? _GEN_391 : _GEN_95; // @[sequencer-master.scala 154:24]
  wire  _GEN_400 = _GEN_32729 | _GEN_112; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_401 = _GEN_32730 | _GEN_113; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_402 = _GEN_32731 | _GEN_114; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_403 = _GEN_32732 | _GEN_115; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_404 = _GEN_32733 | _GEN_116; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_405 = _GEN_32734 | _GEN_117; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_406 = _GEN_32735 | _GEN_118; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_407 = _GEN_32736 | _GEN_119; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_408 = _T_70 ? _GEN_400 : _GEN_112; // @[sequencer-master.scala 154:24]
  wire  _GEN_409 = _T_70 ? _GEN_401 : _GEN_113; // @[sequencer-master.scala 154:24]
  wire  _GEN_410 = _T_70 ? _GEN_402 : _GEN_114; // @[sequencer-master.scala 154:24]
  wire  _GEN_411 = _T_70 ? _GEN_403 : _GEN_115; // @[sequencer-master.scala 154:24]
  wire  _GEN_412 = _T_70 ? _GEN_404 : _GEN_116; // @[sequencer-master.scala 154:24]
  wire  _GEN_413 = _T_70 ? _GEN_405 : _GEN_117; // @[sequencer-master.scala 154:24]
  wire  _GEN_414 = _T_70 ? _GEN_406 : _GEN_118; // @[sequencer-master.scala 154:24]
  wire  _GEN_415 = _T_70 ? _GEN_407 : _GEN_119; // @[sequencer-master.scala 154:24]
  wire  _GEN_416 = _GEN_32729 | _GEN_136; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_417 = _GEN_32730 | _GEN_137; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_418 = _GEN_32731 | _GEN_138; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_419 = _GEN_32732 | _GEN_139; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_420 = _GEN_32733 | _GEN_140; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_421 = _GEN_32734 | _GEN_141; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_422 = _GEN_32735 | _GEN_142; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_423 = _GEN_32736 | _GEN_143; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_424 = _T_92 ? _GEN_416 : _GEN_136; // @[sequencer-master.scala 154:24]
  wire  _GEN_425 = _T_92 ? _GEN_417 : _GEN_137; // @[sequencer-master.scala 154:24]
  wire  _GEN_426 = _T_92 ? _GEN_418 : _GEN_138; // @[sequencer-master.scala 154:24]
  wire  _GEN_427 = _T_92 ? _GEN_419 : _GEN_139; // @[sequencer-master.scala 154:24]
  wire  _GEN_428 = _T_92 ? _GEN_420 : _GEN_140; // @[sequencer-master.scala 154:24]
  wire  _GEN_429 = _T_92 ? _GEN_421 : _GEN_141; // @[sequencer-master.scala 154:24]
  wire  _GEN_430 = _T_92 ? _GEN_422 : _GEN_142; // @[sequencer-master.scala 154:24]
  wire  _GEN_431 = _T_92 ? _GEN_423 : _GEN_143; // @[sequencer-master.scala 154:24]
  wire  _GEN_432 = _GEN_32729 | _GEN_160; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_433 = _GEN_32730 | _GEN_161; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_434 = _GEN_32731 | _GEN_162; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_435 = _GEN_32732 | _GEN_163; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_436 = _GEN_32733 | _GEN_164; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_437 = _GEN_32734 | _GEN_165; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_438 = _GEN_32735 | _GEN_166; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_439 = _GEN_32736 | _GEN_167; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_440 = _T_114 ? _GEN_432 : _GEN_160; // @[sequencer-master.scala 154:24]
  wire  _GEN_441 = _T_114 ? _GEN_433 : _GEN_161; // @[sequencer-master.scala 154:24]
  wire  _GEN_442 = _T_114 ? _GEN_434 : _GEN_162; // @[sequencer-master.scala 154:24]
  wire  _GEN_443 = _T_114 ? _GEN_435 : _GEN_163; // @[sequencer-master.scala 154:24]
  wire  _GEN_444 = _T_114 ? _GEN_436 : _GEN_164; // @[sequencer-master.scala 154:24]
  wire  _GEN_445 = _T_114 ? _GEN_437 : _GEN_165; // @[sequencer-master.scala 154:24]
  wire  _GEN_446 = _T_114 ? _GEN_438 : _GEN_166; // @[sequencer-master.scala 154:24]
  wire  _GEN_447 = _T_114 ? _GEN_439 : _GEN_167; // @[sequencer-master.scala 154:24]
  wire  _GEN_448 = _GEN_32729 | _GEN_184; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_449 = _GEN_32730 | _GEN_185; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_450 = _GEN_32731 | _GEN_186; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_451 = _GEN_32732 | _GEN_187; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_452 = _GEN_32733 | _GEN_188; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_453 = _GEN_32734 | _GEN_189; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_454 = _GEN_32735 | _GEN_190; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_455 = _GEN_32736 | _GEN_191; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_456 = _T_136 ? _GEN_448 : _GEN_184; // @[sequencer-master.scala 154:24]
  wire  _GEN_457 = _T_136 ? _GEN_449 : _GEN_185; // @[sequencer-master.scala 154:24]
  wire  _GEN_458 = _T_136 ? _GEN_450 : _GEN_186; // @[sequencer-master.scala 154:24]
  wire  _GEN_459 = _T_136 ? _GEN_451 : _GEN_187; // @[sequencer-master.scala 154:24]
  wire  _GEN_460 = _T_136 ? _GEN_452 : _GEN_188; // @[sequencer-master.scala 154:24]
  wire  _GEN_461 = _T_136 ? _GEN_453 : _GEN_189; // @[sequencer-master.scala 154:24]
  wire  _GEN_462 = _T_136 ? _GEN_454 : _GEN_190; // @[sequencer-master.scala 154:24]
  wire  _GEN_463 = _T_136 ? _GEN_455 : _GEN_191; // @[sequencer-master.scala 154:24]
  wire  _GEN_464 = _GEN_32729 | _GEN_208; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_465 = _GEN_32730 | _GEN_209; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_466 = _GEN_32731 | _GEN_210; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_467 = _GEN_32732 | _GEN_211; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_468 = _GEN_32733 | _GEN_212; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_469 = _GEN_32734 | _GEN_213; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_470 = _GEN_32735 | _GEN_214; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_471 = _GEN_32736 | _GEN_215; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_472 = _T_158 ? _GEN_464 : _GEN_208; // @[sequencer-master.scala 154:24]
  wire  _GEN_473 = _T_158 ? _GEN_465 : _GEN_209; // @[sequencer-master.scala 154:24]
  wire  _GEN_474 = _T_158 ? _GEN_466 : _GEN_210; // @[sequencer-master.scala 154:24]
  wire  _GEN_475 = _T_158 ? _GEN_467 : _GEN_211; // @[sequencer-master.scala 154:24]
  wire  _GEN_476 = _T_158 ? _GEN_468 : _GEN_212; // @[sequencer-master.scala 154:24]
  wire  _GEN_477 = _T_158 ? _GEN_469 : _GEN_213; // @[sequencer-master.scala 154:24]
  wire  _GEN_478 = _T_158 ? _GEN_470 : _GEN_214; // @[sequencer-master.scala 154:24]
  wire  _GEN_479 = _T_158 ? _GEN_471 : _GEN_215; // @[sequencer-master.scala 154:24]
  wire  _GEN_480 = _GEN_32729 | _GEN_232; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_481 = _GEN_32730 | _GEN_233; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_482 = _GEN_32731 | _GEN_234; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_483 = _GEN_32732 | _GEN_235; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_484 = _GEN_32733 | _GEN_236; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_485 = _GEN_32734 | _GEN_237; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_486 = _GEN_32735 | _GEN_238; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_487 = _GEN_32736 | _GEN_239; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_488 = _T_180 ? _GEN_480 : _GEN_232; // @[sequencer-master.scala 154:24]
  wire  _GEN_489 = _T_180 ? _GEN_481 : _GEN_233; // @[sequencer-master.scala 154:24]
  wire  _GEN_490 = _T_180 ? _GEN_482 : _GEN_234; // @[sequencer-master.scala 154:24]
  wire  _GEN_491 = _T_180 ? _GEN_483 : _GEN_235; // @[sequencer-master.scala 154:24]
  wire  _GEN_492 = _T_180 ? _GEN_484 : _GEN_236; // @[sequencer-master.scala 154:24]
  wire  _GEN_493 = _T_180 ? _GEN_485 : _GEN_237; // @[sequencer-master.scala 154:24]
  wire  _GEN_494 = _T_180 ? _GEN_486 : _GEN_238; // @[sequencer-master.scala 154:24]
  wire  _GEN_495 = _T_180 ? _GEN_487 : _GEN_239; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_496 = 3'h0 == tail ? io_op_bits_base_vs1_id : e_0_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_497 = 3'h1 == tail ? io_op_bits_base_vs1_id : e_1_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_498 = 3'h2 == tail ? io_op_bits_base_vs1_id : e_2_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_499 = 3'h3 == tail ? io_op_bits_base_vs1_id : e_3_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_500 = 3'h4 == tail ? io_op_bits_base_vs1_id : e_4_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_501 = 3'h5 == tail ? io_op_bits_base_vs1_id : e_5_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_502 = 3'h6 == tail ? io_op_bits_base_vs1_id : e_6_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_503 = 3'h7 == tail ? io_op_bits_base_vs1_id : e_7_base_vs1_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_504 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_24; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_505 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_25; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_506 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_26; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_507 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_27; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_508 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_28; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_509 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_29; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_510 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_30; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_511 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_31; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_512 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : e_0_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_513 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : e_1_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_514 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : e_2_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_515 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : e_3_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_516 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : e_4_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_517 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : e_5_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_518 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : e_6_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_519 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : e_7_base_vs1_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_520 = 3'h0 == tail ? io_op_bits_base_vs1_pred : e_0_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_521 = 3'h1 == tail ? io_op_bits_base_vs1_pred : e_1_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_522 = 3'h2 == tail ? io_op_bits_base_vs1_pred : e_2_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_523 = 3'h3 == tail ? io_op_bits_base_vs1_pred : e_3_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_524 = 3'h4 == tail ? io_op_bits_base_vs1_pred : e_4_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_525 = 3'h5 == tail ? io_op_bits_base_vs1_pred : e_5_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_526 = 3'h6 == tail ? io_op_bits_base_vs1_pred : e_6_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_527 = 3'h7 == tail ? io_op_bits_base_vs1_pred : e_7_base_vs1_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_528 = 3'h0 == tail ? io_op_bits_base_vs1_prec : e_0_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_529 = 3'h1 == tail ? io_op_bits_base_vs1_prec : e_1_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_530 = 3'h2 == tail ? io_op_bits_base_vs1_prec : e_2_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_531 = 3'h3 == tail ? io_op_bits_base_vs1_prec : e_3_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_532 = 3'h4 == tail ? io_op_bits_base_vs1_prec : e_4_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_533 = 3'h5 == tail ? io_op_bits_base_vs1_prec : e_5_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_534 = 3'h6 == tail ? io_op_bits_base_vs1_prec : e_6_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_535 = 3'h7 == tail ? io_op_bits_base_vs1_prec : e_7_base_vs1_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_536 = 3'h0 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_537 = 3'h1 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_538 = 3'h2 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_539 = 3'h3 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_540 = 3'h4 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_541 = 3'h5 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_542 = 3'h6 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_543 = 3'h7 == tail ? io_op_bits_reg_vs1_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [63:0] _GEN_544 = 3'h0 == tail ? io_op_bits_sreg_ss1 : e_0_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_545 = 3'h1 == tail ? io_op_bits_sreg_ss1 : e_1_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_546 = 3'h2 == tail ? io_op_bits_sreg_ss1 : e_2_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_547 = 3'h3 == tail ? io_op_bits_sreg_ss1 : e_3_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_548 = 3'h4 == tail ? io_op_bits_sreg_ss1 : e_4_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_549 = 3'h5 == tail ? io_op_bits_sreg_ss1 : e_5_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_550 = 3'h6 == tail ? io_op_bits_sreg_ss1 : e_6_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_551 = 3'h7 == tail ? io_op_bits_sreg_ss1 : e_7_sreg_ss1; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_552 = _T_189 ? _GEN_544 : e_0_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_553 = _T_189 ? _GEN_545 : e_1_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_554 = _T_189 ? _GEN_546 : e_2_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_555 = _T_189 ? _GEN_547 : e_3_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_556 = _T_189 ? _GEN_548 : e_4_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_557 = _T_189 ? _GEN_549 : e_5_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_558 = _T_189 ? _GEN_550 : e_6_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_559 = _T_189 ? _GEN_551 : e_7_sreg_ss1; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [7:0] _GEN_560 = io_op_bits_base_vs1_valid ? _GEN_496 : e_0_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_561 = io_op_bits_base_vs1_valid ? _GEN_497 : e_1_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_562 = io_op_bits_base_vs1_valid ? _GEN_498 : e_2_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_563 = io_op_bits_base_vs1_valid ? _GEN_499 : e_3_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_564 = io_op_bits_base_vs1_valid ? _GEN_500 : e_4_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_565 = io_op_bits_base_vs1_valid ? _GEN_501 : e_5_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_566 = io_op_bits_base_vs1_valid ? _GEN_502 : e_6_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_567 = io_op_bits_base_vs1_valid ? _GEN_503 : e_7_base_vs1_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_568 = io_op_bits_base_vs1_valid ? _GEN_504 : _GEN_24; // @[sequencer-master.scala 328:47]
  wire  _GEN_569 = io_op_bits_base_vs1_valid ? _GEN_505 : _GEN_25; // @[sequencer-master.scala 328:47]
  wire  _GEN_570 = io_op_bits_base_vs1_valid ? _GEN_506 : _GEN_26; // @[sequencer-master.scala 328:47]
  wire  _GEN_571 = io_op_bits_base_vs1_valid ? _GEN_507 : _GEN_27; // @[sequencer-master.scala 328:47]
  wire  _GEN_572 = io_op_bits_base_vs1_valid ? _GEN_508 : _GEN_28; // @[sequencer-master.scala 328:47]
  wire  _GEN_573 = io_op_bits_base_vs1_valid ? _GEN_509 : _GEN_29; // @[sequencer-master.scala 328:47]
  wire  _GEN_574 = io_op_bits_base_vs1_valid ? _GEN_510 : _GEN_30; // @[sequencer-master.scala 328:47]
  wire  _GEN_575 = io_op_bits_base_vs1_valid ? _GEN_511 : _GEN_31; // @[sequencer-master.scala 328:47]
  wire  _GEN_576 = io_op_bits_base_vs1_valid ? _GEN_512 : e_0_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_577 = io_op_bits_base_vs1_valid ? _GEN_513 : e_1_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_578 = io_op_bits_base_vs1_valid ? _GEN_514 : e_2_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_579 = io_op_bits_base_vs1_valid ? _GEN_515 : e_3_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_580 = io_op_bits_base_vs1_valid ? _GEN_516 : e_4_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_581 = io_op_bits_base_vs1_valid ? _GEN_517 : e_5_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_582 = io_op_bits_base_vs1_valid ? _GEN_518 : e_6_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_583 = io_op_bits_base_vs1_valid ? _GEN_519 : e_7_base_vs1_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_584 = io_op_bits_base_vs1_valid ? _GEN_520 : e_0_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_585 = io_op_bits_base_vs1_valid ? _GEN_521 : e_1_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_586 = io_op_bits_base_vs1_valid ? _GEN_522 : e_2_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_587 = io_op_bits_base_vs1_valid ? _GEN_523 : e_3_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_588 = io_op_bits_base_vs1_valid ? _GEN_524 : e_4_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_589 = io_op_bits_base_vs1_valid ? _GEN_525 : e_5_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_590 = io_op_bits_base_vs1_valid ? _GEN_526 : e_6_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_591 = io_op_bits_base_vs1_valid ? _GEN_527 : e_7_base_vs1_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_592 = io_op_bits_base_vs1_valid ? _GEN_528 : e_0_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_593 = io_op_bits_base_vs1_valid ? _GEN_529 : e_1_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_594 = io_op_bits_base_vs1_valid ? _GEN_530 : e_2_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_595 = io_op_bits_base_vs1_valid ? _GEN_531 : e_3_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_596 = io_op_bits_base_vs1_valid ? _GEN_532 : e_4_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_597 = io_op_bits_base_vs1_valid ? _GEN_533 : e_5_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_598 = io_op_bits_base_vs1_valid ? _GEN_534 : e_6_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_599 = io_op_bits_base_vs1_valid ? _GEN_535 : e_7_base_vs1_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_600 = io_op_bits_base_vs1_valid ? _GEN_536 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_601 = io_op_bits_base_vs1_valid ? _GEN_537 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_602 = io_op_bits_base_vs1_valid ? _GEN_538 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_603 = io_op_bits_base_vs1_valid ? _GEN_539 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_604 = io_op_bits_base_vs1_valid ? _GEN_540 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_605 = io_op_bits_base_vs1_valid ? _GEN_541 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_606 = io_op_bits_base_vs1_valid ? _GEN_542 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_607 = io_op_bits_base_vs1_valid ? _GEN_543 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [63:0] _GEN_608 = io_op_bits_base_vs1_valid ? _GEN_552 : e_0_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_609 = io_op_bits_base_vs1_valid ? _GEN_553 : e_1_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_610 = io_op_bits_base_vs1_valid ? _GEN_554 : e_2_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_611 = io_op_bits_base_vs1_valid ? _GEN_555 : e_3_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_612 = io_op_bits_base_vs1_valid ? _GEN_556 : e_4_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_613 = io_op_bits_base_vs1_valid ? _GEN_557 : e_5_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_614 = io_op_bits_base_vs1_valid ? _GEN_558 : e_6_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_615 = io_op_bits_base_vs1_valid ? _GEN_559 : e_7_sreg_ss1; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_616 = _GEN_32729 | _GEN_376; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_617 = _GEN_32730 | _GEN_377; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_618 = _GEN_32731 | _GEN_378; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_619 = _GEN_32732 | _GEN_379; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_620 = _GEN_32733 | _GEN_380; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_621 = _GEN_32734 | _GEN_381; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_622 = _GEN_32735 | _GEN_382; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_623 = _GEN_32736 | _GEN_383; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_624 = _T_203 ? _GEN_616 : _GEN_376; // @[sequencer-master.scala 154:24]
  wire  _GEN_625 = _T_203 ? _GEN_617 : _GEN_377; // @[sequencer-master.scala 154:24]
  wire  _GEN_626 = _T_203 ? _GEN_618 : _GEN_378; // @[sequencer-master.scala 154:24]
  wire  _GEN_627 = _T_203 ? _GEN_619 : _GEN_379; // @[sequencer-master.scala 154:24]
  wire  _GEN_628 = _T_203 ? _GEN_620 : _GEN_380; // @[sequencer-master.scala 154:24]
  wire  _GEN_629 = _T_203 ? _GEN_621 : _GEN_381; // @[sequencer-master.scala 154:24]
  wire  _GEN_630 = _T_203 ? _GEN_622 : _GEN_382; // @[sequencer-master.scala 154:24]
  wire  _GEN_631 = _T_203 ? _GEN_623 : _GEN_383; // @[sequencer-master.scala 154:24]
  wire  _GEN_632 = _GEN_32729 | _GEN_392; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_633 = _GEN_32730 | _GEN_393; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_634 = _GEN_32731 | _GEN_394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_635 = _GEN_32732 | _GEN_395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_636 = _GEN_32733 | _GEN_396; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_637 = _GEN_32734 | _GEN_397; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_638 = _GEN_32735 | _GEN_398; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_639 = _GEN_32736 | _GEN_399; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_640 = _T_225 ? _GEN_632 : _GEN_392; // @[sequencer-master.scala 154:24]
  wire  _GEN_641 = _T_225 ? _GEN_633 : _GEN_393; // @[sequencer-master.scala 154:24]
  wire  _GEN_642 = _T_225 ? _GEN_634 : _GEN_394; // @[sequencer-master.scala 154:24]
  wire  _GEN_643 = _T_225 ? _GEN_635 : _GEN_395; // @[sequencer-master.scala 154:24]
  wire  _GEN_644 = _T_225 ? _GEN_636 : _GEN_396; // @[sequencer-master.scala 154:24]
  wire  _GEN_645 = _T_225 ? _GEN_637 : _GEN_397; // @[sequencer-master.scala 154:24]
  wire  _GEN_646 = _T_225 ? _GEN_638 : _GEN_398; // @[sequencer-master.scala 154:24]
  wire  _GEN_647 = _T_225 ? _GEN_639 : _GEN_399; // @[sequencer-master.scala 154:24]
  wire  _GEN_648 = _GEN_32729 | _GEN_408; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_649 = _GEN_32730 | _GEN_409; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_650 = _GEN_32731 | _GEN_410; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_651 = _GEN_32732 | _GEN_411; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_652 = _GEN_32733 | _GEN_412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_653 = _GEN_32734 | _GEN_413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_654 = _GEN_32735 | _GEN_414; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_655 = _GEN_32736 | _GEN_415; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_656 = _T_247 ? _GEN_648 : _GEN_408; // @[sequencer-master.scala 154:24]
  wire  _GEN_657 = _T_247 ? _GEN_649 : _GEN_409; // @[sequencer-master.scala 154:24]
  wire  _GEN_658 = _T_247 ? _GEN_650 : _GEN_410; // @[sequencer-master.scala 154:24]
  wire  _GEN_659 = _T_247 ? _GEN_651 : _GEN_411; // @[sequencer-master.scala 154:24]
  wire  _GEN_660 = _T_247 ? _GEN_652 : _GEN_412; // @[sequencer-master.scala 154:24]
  wire  _GEN_661 = _T_247 ? _GEN_653 : _GEN_413; // @[sequencer-master.scala 154:24]
  wire  _GEN_662 = _T_247 ? _GEN_654 : _GEN_414; // @[sequencer-master.scala 154:24]
  wire  _GEN_663 = _T_247 ? _GEN_655 : _GEN_415; // @[sequencer-master.scala 154:24]
  wire  _GEN_664 = _GEN_32729 | _GEN_424; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_665 = _GEN_32730 | _GEN_425; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_666 = _GEN_32731 | _GEN_426; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_667 = _GEN_32732 | _GEN_427; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_668 = _GEN_32733 | _GEN_428; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_669 = _GEN_32734 | _GEN_429; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_670 = _GEN_32735 | _GEN_430; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_671 = _GEN_32736 | _GEN_431; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_672 = _T_269 ? _GEN_664 : _GEN_424; // @[sequencer-master.scala 154:24]
  wire  _GEN_673 = _T_269 ? _GEN_665 : _GEN_425; // @[sequencer-master.scala 154:24]
  wire  _GEN_674 = _T_269 ? _GEN_666 : _GEN_426; // @[sequencer-master.scala 154:24]
  wire  _GEN_675 = _T_269 ? _GEN_667 : _GEN_427; // @[sequencer-master.scala 154:24]
  wire  _GEN_676 = _T_269 ? _GEN_668 : _GEN_428; // @[sequencer-master.scala 154:24]
  wire  _GEN_677 = _T_269 ? _GEN_669 : _GEN_429; // @[sequencer-master.scala 154:24]
  wire  _GEN_678 = _T_269 ? _GEN_670 : _GEN_430; // @[sequencer-master.scala 154:24]
  wire  _GEN_679 = _T_269 ? _GEN_671 : _GEN_431; // @[sequencer-master.scala 154:24]
  wire  _GEN_680 = _GEN_32729 | _GEN_440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_681 = _GEN_32730 | _GEN_441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_682 = _GEN_32731 | _GEN_442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_683 = _GEN_32732 | _GEN_443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_684 = _GEN_32733 | _GEN_444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_685 = _GEN_32734 | _GEN_445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_686 = _GEN_32735 | _GEN_446; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_687 = _GEN_32736 | _GEN_447; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_688 = _T_291 ? _GEN_680 : _GEN_440; // @[sequencer-master.scala 154:24]
  wire  _GEN_689 = _T_291 ? _GEN_681 : _GEN_441; // @[sequencer-master.scala 154:24]
  wire  _GEN_690 = _T_291 ? _GEN_682 : _GEN_442; // @[sequencer-master.scala 154:24]
  wire  _GEN_691 = _T_291 ? _GEN_683 : _GEN_443; // @[sequencer-master.scala 154:24]
  wire  _GEN_692 = _T_291 ? _GEN_684 : _GEN_444; // @[sequencer-master.scala 154:24]
  wire  _GEN_693 = _T_291 ? _GEN_685 : _GEN_445; // @[sequencer-master.scala 154:24]
  wire  _GEN_694 = _T_291 ? _GEN_686 : _GEN_446; // @[sequencer-master.scala 154:24]
  wire  _GEN_695 = _T_291 ? _GEN_687 : _GEN_447; // @[sequencer-master.scala 154:24]
  wire  _GEN_696 = _GEN_32729 | _GEN_456; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_697 = _GEN_32730 | _GEN_457; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_698 = _GEN_32731 | _GEN_458; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_699 = _GEN_32732 | _GEN_459; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_700 = _GEN_32733 | _GEN_460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_701 = _GEN_32734 | _GEN_461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_702 = _GEN_32735 | _GEN_462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_703 = _GEN_32736 | _GEN_463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_704 = _T_313 ? _GEN_696 : _GEN_456; // @[sequencer-master.scala 154:24]
  wire  _GEN_705 = _T_313 ? _GEN_697 : _GEN_457; // @[sequencer-master.scala 154:24]
  wire  _GEN_706 = _T_313 ? _GEN_698 : _GEN_458; // @[sequencer-master.scala 154:24]
  wire  _GEN_707 = _T_313 ? _GEN_699 : _GEN_459; // @[sequencer-master.scala 154:24]
  wire  _GEN_708 = _T_313 ? _GEN_700 : _GEN_460; // @[sequencer-master.scala 154:24]
  wire  _GEN_709 = _T_313 ? _GEN_701 : _GEN_461; // @[sequencer-master.scala 154:24]
  wire  _GEN_710 = _T_313 ? _GEN_702 : _GEN_462; // @[sequencer-master.scala 154:24]
  wire  _GEN_711 = _T_313 ? _GEN_703 : _GEN_463; // @[sequencer-master.scala 154:24]
  wire  _GEN_712 = _GEN_32729 | _GEN_472; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_713 = _GEN_32730 | _GEN_473; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_714 = _GEN_32731 | _GEN_474; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_715 = _GEN_32732 | _GEN_475; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_716 = _GEN_32733 | _GEN_476; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_717 = _GEN_32734 | _GEN_477; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_718 = _GEN_32735 | _GEN_478; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_719 = _GEN_32736 | _GEN_479; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_720 = _T_335 ? _GEN_712 : _GEN_472; // @[sequencer-master.scala 154:24]
  wire  _GEN_721 = _T_335 ? _GEN_713 : _GEN_473; // @[sequencer-master.scala 154:24]
  wire  _GEN_722 = _T_335 ? _GEN_714 : _GEN_474; // @[sequencer-master.scala 154:24]
  wire  _GEN_723 = _T_335 ? _GEN_715 : _GEN_475; // @[sequencer-master.scala 154:24]
  wire  _GEN_724 = _T_335 ? _GEN_716 : _GEN_476; // @[sequencer-master.scala 154:24]
  wire  _GEN_725 = _T_335 ? _GEN_717 : _GEN_477; // @[sequencer-master.scala 154:24]
  wire  _GEN_726 = _T_335 ? _GEN_718 : _GEN_478; // @[sequencer-master.scala 154:24]
  wire  _GEN_727 = _T_335 ? _GEN_719 : _GEN_479; // @[sequencer-master.scala 154:24]
  wire  _GEN_728 = _GEN_32729 | _GEN_488; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_729 = _GEN_32730 | _GEN_489; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_730 = _GEN_32731 | _GEN_490; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_731 = _GEN_32732 | _GEN_491; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_732 = _GEN_32733 | _GEN_492; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_733 = _GEN_32734 | _GEN_493; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_734 = _GEN_32735 | _GEN_494; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_735 = _GEN_32736 | _GEN_495; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_736 = _T_357 ? _GEN_728 : _GEN_488; // @[sequencer-master.scala 154:24]
  wire  _GEN_737 = _T_357 ? _GEN_729 : _GEN_489; // @[sequencer-master.scala 154:24]
  wire  _GEN_738 = _T_357 ? _GEN_730 : _GEN_490; // @[sequencer-master.scala 154:24]
  wire  _GEN_739 = _T_357 ? _GEN_731 : _GEN_491; // @[sequencer-master.scala 154:24]
  wire  _GEN_740 = _T_357 ? _GEN_732 : _GEN_492; // @[sequencer-master.scala 154:24]
  wire  _GEN_741 = _T_357 ? _GEN_733 : _GEN_493; // @[sequencer-master.scala 154:24]
  wire  _GEN_742 = _T_357 ? _GEN_734 : _GEN_494; // @[sequencer-master.scala 154:24]
  wire  _GEN_743 = _T_357 ? _GEN_735 : _GEN_495; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_744 = 3'h0 == tail ? io_op_bits_base_vs2_id : e_0_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_745 = 3'h1 == tail ? io_op_bits_base_vs2_id : e_1_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_746 = 3'h2 == tail ? io_op_bits_base_vs2_id : e_2_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_747 = 3'h3 == tail ? io_op_bits_base_vs2_id : e_3_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_748 = 3'h4 == tail ? io_op_bits_base_vs2_id : e_4_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_749 = 3'h5 == tail ? io_op_bits_base_vs2_id : e_5_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_750 = 3'h6 == tail ? io_op_bits_base_vs2_id : e_6_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_751 = 3'h7 == tail ? io_op_bits_base_vs2_id : e_7_base_vs2_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_752 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_32; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_753 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_33; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_754 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_34; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_755 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_35; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_756 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_36; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_757 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_37; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_758 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_38; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_759 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_39; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_760 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : e_0_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_761 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : e_1_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_762 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : e_2_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_763 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : e_3_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_764 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : e_4_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_765 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : e_5_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_766 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : e_6_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_767 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : e_7_base_vs2_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_768 = 3'h0 == tail ? io_op_bits_base_vs2_pred : e_0_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_769 = 3'h1 == tail ? io_op_bits_base_vs2_pred : e_1_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_770 = 3'h2 == tail ? io_op_bits_base_vs2_pred : e_2_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_771 = 3'h3 == tail ? io_op_bits_base_vs2_pred : e_3_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_772 = 3'h4 == tail ? io_op_bits_base_vs2_pred : e_4_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_773 = 3'h5 == tail ? io_op_bits_base_vs2_pred : e_5_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_774 = 3'h6 == tail ? io_op_bits_base_vs2_pred : e_6_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_775 = 3'h7 == tail ? io_op_bits_base_vs2_pred : e_7_base_vs2_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_776 = 3'h0 == tail ? io_op_bits_base_vs2_prec : e_0_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_777 = 3'h1 == tail ? io_op_bits_base_vs2_prec : e_1_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_778 = 3'h2 == tail ? io_op_bits_base_vs2_prec : e_2_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_779 = 3'h3 == tail ? io_op_bits_base_vs2_prec : e_3_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_780 = 3'h4 == tail ? io_op_bits_base_vs2_prec : e_4_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_781 = 3'h5 == tail ? io_op_bits_base_vs2_prec : e_5_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_782 = 3'h6 == tail ? io_op_bits_base_vs2_prec : e_6_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_783 = 3'h7 == tail ? io_op_bits_base_vs2_prec : e_7_base_vs2_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_784 = 3'h0 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_785 = 3'h1 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_786 = 3'h2 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_787 = 3'h3 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_788 = 3'h4 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_789 = 3'h5 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_790 = 3'h6 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_791 = 3'h7 == tail ? io_op_bits_reg_vs2_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [63:0] _GEN_792 = 3'h0 == tail ? io_op_bits_sreg_ss2 : e_0_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_793 = 3'h1 == tail ? io_op_bits_sreg_ss2 : e_1_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_794 = 3'h2 == tail ? io_op_bits_sreg_ss2 : e_2_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_795 = 3'h3 == tail ? io_op_bits_sreg_ss2 : e_3_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_796 = 3'h4 == tail ? io_op_bits_sreg_ss2 : e_4_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_797 = 3'h5 == tail ? io_op_bits_sreg_ss2 : e_5_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_798 = 3'h6 == tail ? io_op_bits_sreg_ss2 : e_6_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_799 = 3'h7 == tail ? io_op_bits_sreg_ss2 : e_7_sreg_ss2; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_800 = _T_366 ? _GEN_792 : e_0_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_801 = _T_366 ? _GEN_793 : e_1_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_802 = _T_366 ? _GEN_794 : e_2_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_803 = _T_366 ? _GEN_795 : e_3_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_804 = _T_366 ? _GEN_796 : e_4_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_805 = _T_366 ? _GEN_797 : e_5_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_806 = _T_366 ? _GEN_798 : e_6_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_807 = _T_366 ? _GEN_799 : e_7_sreg_ss2; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [7:0] _GEN_808 = io_op_bits_base_vs2_valid ? _GEN_744 : e_0_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_809 = io_op_bits_base_vs2_valid ? _GEN_745 : e_1_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_810 = io_op_bits_base_vs2_valid ? _GEN_746 : e_2_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_811 = io_op_bits_base_vs2_valid ? _GEN_747 : e_3_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_812 = io_op_bits_base_vs2_valid ? _GEN_748 : e_4_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_813 = io_op_bits_base_vs2_valid ? _GEN_749 : e_5_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_814 = io_op_bits_base_vs2_valid ? _GEN_750 : e_6_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_815 = io_op_bits_base_vs2_valid ? _GEN_751 : e_7_base_vs2_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_816 = io_op_bits_base_vs2_valid ? _GEN_752 : _GEN_32; // @[sequencer-master.scala 328:47]
  wire  _GEN_817 = io_op_bits_base_vs2_valid ? _GEN_753 : _GEN_33; // @[sequencer-master.scala 328:47]
  wire  _GEN_818 = io_op_bits_base_vs2_valid ? _GEN_754 : _GEN_34; // @[sequencer-master.scala 328:47]
  wire  _GEN_819 = io_op_bits_base_vs2_valid ? _GEN_755 : _GEN_35; // @[sequencer-master.scala 328:47]
  wire  _GEN_820 = io_op_bits_base_vs2_valid ? _GEN_756 : _GEN_36; // @[sequencer-master.scala 328:47]
  wire  _GEN_821 = io_op_bits_base_vs2_valid ? _GEN_757 : _GEN_37; // @[sequencer-master.scala 328:47]
  wire  _GEN_822 = io_op_bits_base_vs2_valid ? _GEN_758 : _GEN_38; // @[sequencer-master.scala 328:47]
  wire  _GEN_823 = io_op_bits_base_vs2_valid ? _GEN_759 : _GEN_39; // @[sequencer-master.scala 328:47]
  wire  _GEN_824 = io_op_bits_base_vs2_valid ? _GEN_760 : e_0_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_825 = io_op_bits_base_vs2_valid ? _GEN_761 : e_1_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_826 = io_op_bits_base_vs2_valid ? _GEN_762 : e_2_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_827 = io_op_bits_base_vs2_valid ? _GEN_763 : e_3_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_828 = io_op_bits_base_vs2_valid ? _GEN_764 : e_4_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_829 = io_op_bits_base_vs2_valid ? _GEN_765 : e_5_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_830 = io_op_bits_base_vs2_valid ? _GEN_766 : e_6_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_831 = io_op_bits_base_vs2_valid ? _GEN_767 : e_7_base_vs2_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_832 = io_op_bits_base_vs2_valid ? _GEN_768 : e_0_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_833 = io_op_bits_base_vs2_valid ? _GEN_769 : e_1_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_834 = io_op_bits_base_vs2_valid ? _GEN_770 : e_2_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_835 = io_op_bits_base_vs2_valid ? _GEN_771 : e_3_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_836 = io_op_bits_base_vs2_valid ? _GEN_772 : e_4_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_837 = io_op_bits_base_vs2_valid ? _GEN_773 : e_5_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_838 = io_op_bits_base_vs2_valid ? _GEN_774 : e_6_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_839 = io_op_bits_base_vs2_valid ? _GEN_775 : e_7_base_vs2_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_840 = io_op_bits_base_vs2_valid ? _GEN_776 : e_0_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_841 = io_op_bits_base_vs2_valid ? _GEN_777 : e_1_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_842 = io_op_bits_base_vs2_valid ? _GEN_778 : e_2_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_843 = io_op_bits_base_vs2_valid ? _GEN_779 : e_3_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_844 = io_op_bits_base_vs2_valid ? _GEN_780 : e_4_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_845 = io_op_bits_base_vs2_valid ? _GEN_781 : e_5_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_846 = io_op_bits_base_vs2_valid ? _GEN_782 : e_6_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_847 = io_op_bits_base_vs2_valid ? _GEN_783 : e_7_base_vs2_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_848 = io_op_bits_base_vs2_valid ? _GEN_784 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_849 = io_op_bits_base_vs2_valid ? _GEN_785 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_850 = io_op_bits_base_vs2_valid ? _GEN_786 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_851 = io_op_bits_base_vs2_valid ? _GEN_787 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_852 = io_op_bits_base_vs2_valid ? _GEN_788 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_853 = io_op_bits_base_vs2_valid ? _GEN_789 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_854 = io_op_bits_base_vs2_valid ? _GEN_790 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_855 = io_op_bits_base_vs2_valid ? _GEN_791 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [63:0] _GEN_856 = io_op_bits_base_vs2_valid ? _GEN_800 : e_0_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_857 = io_op_bits_base_vs2_valid ? _GEN_801 : e_1_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_858 = io_op_bits_base_vs2_valid ? _GEN_802 : e_2_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_859 = io_op_bits_base_vs2_valid ? _GEN_803 : e_3_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_860 = io_op_bits_base_vs2_valid ? _GEN_804 : e_4_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_861 = io_op_bits_base_vs2_valid ? _GEN_805 : e_5_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_862 = io_op_bits_base_vs2_valid ? _GEN_806 : e_6_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_863 = io_op_bits_base_vs2_valid ? _GEN_807 : e_7_sreg_ss2; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_864 = _GEN_32729 | _GEN_624; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_865 = _GEN_32730 | _GEN_625; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_866 = _GEN_32731 | _GEN_626; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_867 = _GEN_32732 | _GEN_627; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_868 = _GEN_32733 | _GEN_628; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_869 = _GEN_32734 | _GEN_629; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_870 = _GEN_32735 | _GEN_630; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_871 = _GEN_32736 | _GEN_631; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_872 = _T_380 ? _GEN_864 : _GEN_624; // @[sequencer-master.scala 154:24]
  wire  _GEN_873 = _T_380 ? _GEN_865 : _GEN_625; // @[sequencer-master.scala 154:24]
  wire  _GEN_874 = _T_380 ? _GEN_866 : _GEN_626; // @[sequencer-master.scala 154:24]
  wire  _GEN_875 = _T_380 ? _GEN_867 : _GEN_627; // @[sequencer-master.scala 154:24]
  wire  _GEN_876 = _T_380 ? _GEN_868 : _GEN_628; // @[sequencer-master.scala 154:24]
  wire  _GEN_877 = _T_380 ? _GEN_869 : _GEN_629; // @[sequencer-master.scala 154:24]
  wire  _GEN_878 = _T_380 ? _GEN_870 : _GEN_630; // @[sequencer-master.scala 154:24]
  wire  _GEN_879 = _T_380 ? _GEN_871 : _GEN_631; // @[sequencer-master.scala 154:24]
  wire  _GEN_880 = _GEN_32729 | _GEN_640; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_881 = _GEN_32730 | _GEN_641; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_882 = _GEN_32731 | _GEN_642; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_883 = _GEN_32732 | _GEN_643; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_884 = _GEN_32733 | _GEN_644; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_885 = _GEN_32734 | _GEN_645; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_886 = _GEN_32735 | _GEN_646; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_887 = _GEN_32736 | _GEN_647; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_888 = _T_402 ? _GEN_880 : _GEN_640; // @[sequencer-master.scala 154:24]
  wire  _GEN_889 = _T_402 ? _GEN_881 : _GEN_641; // @[sequencer-master.scala 154:24]
  wire  _GEN_890 = _T_402 ? _GEN_882 : _GEN_642; // @[sequencer-master.scala 154:24]
  wire  _GEN_891 = _T_402 ? _GEN_883 : _GEN_643; // @[sequencer-master.scala 154:24]
  wire  _GEN_892 = _T_402 ? _GEN_884 : _GEN_644; // @[sequencer-master.scala 154:24]
  wire  _GEN_893 = _T_402 ? _GEN_885 : _GEN_645; // @[sequencer-master.scala 154:24]
  wire  _GEN_894 = _T_402 ? _GEN_886 : _GEN_646; // @[sequencer-master.scala 154:24]
  wire  _GEN_895 = _T_402 ? _GEN_887 : _GEN_647; // @[sequencer-master.scala 154:24]
  wire  _GEN_896 = _GEN_32729 | _GEN_656; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_897 = _GEN_32730 | _GEN_657; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_898 = _GEN_32731 | _GEN_658; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_899 = _GEN_32732 | _GEN_659; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_900 = _GEN_32733 | _GEN_660; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_901 = _GEN_32734 | _GEN_661; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_902 = _GEN_32735 | _GEN_662; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_903 = _GEN_32736 | _GEN_663; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_904 = _T_424 ? _GEN_896 : _GEN_656; // @[sequencer-master.scala 154:24]
  wire  _GEN_905 = _T_424 ? _GEN_897 : _GEN_657; // @[sequencer-master.scala 154:24]
  wire  _GEN_906 = _T_424 ? _GEN_898 : _GEN_658; // @[sequencer-master.scala 154:24]
  wire  _GEN_907 = _T_424 ? _GEN_899 : _GEN_659; // @[sequencer-master.scala 154:24]
  wire  _GEN_908 = _T_424 ? _GEN_900 : _GEN_660; // @[sequencer-master.scala 154:24]
  wire  _GEN_909 = _T_424 ? _GEN_901 : _GEN_661; // @[sequencer-master.scala 154:24]
  wire  _GEN_910 = _T_424 ? _GEN_902 : _GEN_662; // @[sequencer-master.scala 154:24]
  wire  _GEN_911 = _T_424 ? _GEN_903 : _GEN_663; // @[sequencer-master.scala 154:24]
  wire  _GEN_912 = _GEN_32729 | _GEN_672; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_913 = _GEN_32730 | _GEN_673; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_914 = _GEN_32731 | _GEN_674; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_915 = _GEN_32732 | _GEN_675; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_916 = _GEN_32733 | _GEN_676; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_917 = _GEN_32734 | _GEN_677; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_918 = _GEN_32735 | _GEN_678; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_919 = _GEN_32736 | _GEN_679; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_920 = _T_446 ? _GEN_912 : _GEN_672; // @[sequencer-master.scala 154:24]
  wire  _GEN_921 = _T_446 ? _GEN_913 : _GEN_673; // @[sequencer-master.scala 154:24]
  wire  _GEN_922 = _T_446 ? _GEN_914 : _GEN_674; // @[sequencer-master.scala 154:24]
  wire  _GEN_923 = _T_446 ? _GEN_915 : _GEN_675; // @[sequencer-master.scala 154:24]
  wire  _GEN_924 = _T_446 ? _GEN_916 : _GEN_676; // @[sequencer-master.scala 154:24]
  wire  _GEN_925 = _T_446 ? _GEN_917 : _GEN_677; // @[sequencer-master.scala 154:24]
  wire  _GEN_926 = _T_446 ? _GEN_918 : _GEN_678; // @[sequencer-master.scala 154:24]
  wire  _GEN_927 = _T_446 ? _GEN_919 : _GEN_679; // @[sequencer-master.scala 154:24]
  wire  _GEN_928 = _GEN_32729 | _GEN_688; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_929 = _GEN_32730 | _GEN_689; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_930 = _GEN_32731 | _GEN_690; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_931 = _GEN_32732 | _GEN_691; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_932 = _GEN_32733 | _GEN_692; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_933 = _GEN_32734 | _GEN_693; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_934 = _GEN_32735 | _GEN_694; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_935 = _GEN_32736 | _GEN_695; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_936 = _T_468 ? _GEN_928 : _GEN_688; // @[sequencer-master.scala 154:24]
  wire  _GEN_937 = _T_468 ? _GEN_929 : _GEN_689; // @[sequencer-master.scala 154:24]
  wire  _GEN_938 = _T_468 ? _GEN_930 : _GEN_690; // @[sequencer-master.scala 154:24]
  wire  _GEN_939 = _T_468 ? _GEN_931 : _GEN_691; // @[sequencer-master.scala 154:24]
  wire  _GEN_940 = _T_468 ? _GEN_932 : _GEN_692; // @[sequencer-master.scala 154:24]
  wire  _GEN_941 = _T_468 ? _GEN_933 : _GEN_693; // @[sequencer-master.scala 154:24]
  wire  _GEN_942 = _T_468 ? _GEN_934 : _GEN_694; // @[sequencer-master.scala 154:24]
  wire  _GEN_943 = _T_468 ? _GEN_935 : _GEN_695; // @[sequencer-master.scala 154:24]
  wire  _GEN_944 = _GEN_32729 | _GEN_704; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_945 = _GEN_32730 | _GEN_705; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_946 = _GEN_32731 | _GEN_706; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_947 = _GEN_32732 | _GEN_707; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_948 = _GEN_32733 | _GEN_708; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_949 = _GEN_32734 | _GEN_709; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_950 = _GEN_32735 | _GEN_710; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_951 = _GEN_32736 | _GEN_711; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_952 = _T_490 ? _GEN_944 : _GEN_704; // @[sequencer-master.scala 154:24]
  wire  _GEN_953 = _T_490 ? _GEN_945 : _GEN_705; // @[sequencer-master.scala 154:24]
  wire  _GEN_954 = _T_490 ? _GEN_946 : _GEN_706; // @[sequencer-master.scala 154:24]
  wire  _GEN_955 = _T_490 ? _GEN_947 : _GEN_707; // @[sequencer-master.scala 154:24]
  wire  _GEN_956 = _T_490 ? _GEN_948 : _GEN_708; // @[sequencer-master.scala 154:24]
  wire  _GEN_957 = _T_490 ? _GEN_949 : _GEN_709; // @[sequencer-master.scala 154:24]
  wire  _GEN_958 = _T_490 ? _GEN_950 : _GEN_710; // @[sequencer-master.scala 154:24]
  wire  _GEN_959 = _T_490 ? _GEN_951 : _GEN_711; // @[sequencer-master.scala 154:24]
  wire  _GEN_960 = _GEN_32729 | _GEN_720; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_961 = _GEN_32730 | _GEN_721; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_962 = _GEN_32731 | _GEN_722; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_963 = _GEN_32732 | _GEN_723; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_964 = _GEN_32733 | _GEN_724; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_965 = _GEN_32734 | _GEN_725; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_966 = _GEN_32735 | _GEN_726; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_967 = _GEN_32736 | _GEN_727; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_968 = _T_512 ? _GEN_960 : _GEN_720; // @[sequencer-master.scala 154:24]
  wire  _GEN_969 = _T_512 ? _GEN_961 : _GEN_721; // @[sequencer-master.scala 154:24]
  wire  _GEN_970 = _T_512 ? _GEN_962 : _GEN_722; // @[sequencer-master.scala 154:24]
  wire  _GEN_971 = _T_512 ? _GEN_963 : _GEN_723; // @[sequencer-master.scala 154:24]
  wire  _GEN_972 = _T_512 ? _GEN_964 : _GEN_724; // @[sequencer-master.scala 154:24]
  wire  _GEN_973 = _T_512 ? _GEN_965 : _GEN_725; // @[sequencer-master.scala 154:24]
  wire  _GEN_974 = _T_512 ? _GEN_966 : _GEN_726; // @[sequencer-master.scala 154:24]
  wire  _GEN_975 = _T_512 ? _GEN_967 : _GEN_727; // @[sequencer-master.scala 154:24]
  wire  _GEN_976 = _GEN_32729 | _GEN_736; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_977 = _GEN_32730 | _GEN_737; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_978 = _GEN_32731 | _GEN_738; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_979 = _GEN_32732 | _GEN_739; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_980 = _GEN_32733 | _GEN_740; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_981 = _GEN_32734 | _GEN_741; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_982 = _GEN_32735 | _GEN_742; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_983 = _GEN_32736 | _GEN_743; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_984 = _T_534 ? _GEN_976 : _GEN_736; // @[sequencer-master.scala 154:24]
  wire  _GEN_985 = _T_534 ? _GEN_977 : _GEN_737; // @[sequencer-master.scala 154:24]
  wire  _GEN_986 = _T_534 ? _GEN_978 : _GEN_738; // @[sequencer-master.scala 154:24]
  wire  _GEN_987 = _T_534 ? _GEN_979 : _GEN_739; // @[sequencer-master.scala 154:24]
  wire  _GEN_988 = _T_534 ? _GEN_980 : _GEN_740; // @[sequencer-master.scala 154:24]
  wire  _GEN_989 = _T_534 ? _GEN_981 : _GEN_741; // @[sequencer-master.scala 154:24]
  wire  _GEN_990 = _T_534 ? _GEN_982 : _GEN_742; // @[sequencer-master.scala 154:24]
  wire  _GEN_991 = _T_534 ? _GEN_983 : _GEN_743; // @[sequencer-master.scala 154:24]
  wire  _T_1764 = ~(~io_op_bits_base_vd_valid | _T_721 | reset); // @[sequencer-master.scala 361:15]
  wire [7:0] _GEN_992 = 3'h0 == tail ? io_op_bits_base_vd_id : e_0_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_993 = 3'h1 == tail ? io_op_bits_base_vd_id : e_1_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_994 = 3'h2 == tail ? io_op_bits_base_vd_id : e_2_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_995 = 3'h3 == tail ? io_op_bits_base_vd_id : e_3_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_996 = 3'h4 == tail ? io_op_bits_base_vd_id : e_4_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_997 = 3'h5 == tail ? io_op_bits_base_vd_id : e_5_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_998 = 3'h6 == tail ? io_op_bits_base_vd_id : e_6_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_999 = 3'h7 == tail ? io_op_bits_base_vd_id : e_7_base_vd_id; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1000 = 3'h0 == tail ? io_op_bits_base_vd_valid : _GEN_48; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1001 = 3'h1 == tail ? io_op_bits_base_vd_valid : _GEN_49; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1002 = 3'h2 == tail ? io_op_bits_base_vd_valid : _GEN_50; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1003 = 3'h3 == tail ? io_op_bits_base_vd_valid : _GEN_51; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1004 = 3'h4 == tail ? io_op_bits_base_vd_valid : _GEN_52; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1005 = 3'h5 == tail ? io_op_bits_base_vd_valid : _GEN_53; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1006 = 3'h6 == tail ? io_op_bits_base_vd_valid : _GEN_54; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1007 = 3'h7 == tail ? io_op_bits_base_vd_valid : _GEN_55; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_1008 = 3'h0 == tail ? io_op_bits_base_vd_scalar : e_0_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1009 = 3'h1 == tail ? io_op_bits_base_vd_scalar : e_1_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1010 = 3'h2 == tail ? io_op_bits_base_vd_scalar : e_2_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1011 = 3'h3 == tail ? io_op_bits_base_vd_scalar : e_3_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1012 = 3'h4 == tail ? io_op_bits_base_vd_scalar : e_4_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1013 = 3'h5 == tail ? io_op_bits_base_vd_scalar : e_5_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1014 = 3'h6 == tail ? io_op_bits_base_vd_scalar : e_6_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1015 = 3'h7 == tail ? io_op_bits_base_vd_scalar : e_7_base_vd_scalar; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1016 = 3'h0 == tail ? io_op_bits_base_vd_pred : e_0_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1017 = 3'h1 == tail ? io_op_bits_base_vd_pred : e_1_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1018 = 3'h2 == tail ? io_op_bits_base_vd_pred : e_2_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1019 = 3'h3 == tail ? io_op_bits_base_vd_pred : e_3_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1020 = 3'h4 == tail ? io_op_bits_base_vd_pred : e_4_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1021 = 3'h5 == tail ? io_op_bits_base_vd_pred : e_5_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1022 = 3'h6 == tail ? io_op_bits_base_vd_pred : e_6_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire  _GEN_1023 = 3'h7 == tail ? io_op_bits_base_vd_pred : e_7_base_vd_pred; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1024 = 3'h0 == tail ? io_op_bits_base_vd_prec : e_0_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1025 = 3'h1 == tail ? io_op_bits_base_vd_prec : e_1_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1026 = 3'h2 == tail ? io_op_bits_base_vd_prec : e_2_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1027 = 3'h3 == tail ? io_op_bits_base_vd_prec : e_3_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1028 = 3'h4 == tail ? io_op_bits_base_vd_prec : e_4_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1029 = 3'h5 == tail ? io_op_bits_base_vd_prec : e_5_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1030 = 3'h6 == tail ? io_op_bits_base_vd_prec : e_6_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1031 = 3'h7 == tail ? io_op_bits_base_vd_prec : e_7_base_vd_prec; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1032 = 3'h0 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1033 = 3'h1 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1034 = 3'h2 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1035 = 3'h3 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1036 = 3'h4 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1037 = 3'h5 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1038 = 3'h6 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1039 = 3'h7 == tail ? io_op_bits_reg_vd_id : 8'h0; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1040 = io_op_bits_base_vd_valid ? _GEN_992 : e_0_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1041 = io_op_bits_base_vd_valid ? _GEN_993 : e_1_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1042 = io_op_bits_base_vd_valid ? _GEN_994 : e_2_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1043 = io_op_bits_base_vd_valid ? _GEN_995 : e_3_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1044 = io_op_bits_base_vd_valid ? _GEN_996 : e_4_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1045 = io_op_bits_base_vd_valid ? _GEN_997 : e_5_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1046 = io_op_bits_base_vd_valid ? _GEN_998 : e_6_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1047 = io_op_bits_base_vd_valid ? _GEN_999 : e_7_base_vd_id; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1048 = io_op_bits_base_vd_valid ? _GEN_1000 : _GEN_48; // @[sequencer-master.scala 362:41]
  wire  _GEN_1049 = io_op_bits_base_vd_valid ? _GEN_1001 : _GEN_49; // @[sequencer-master.scala 362:41]
  wire  _GEN_1050 = io_op_bits_base_vd_valid ? _GEN_1002 : _GEN_50; // @[sequencer-master.scala 362:41]
  wire  _GEN_1051 = io_op_bits_base_vd_valid ? _GEN_1003 : _GEN_51; // @[sequencer-master.scala 362:41]
  wire  _GEN_1052 = io_op_bits_base_vd_valid ? _GEN_1004 : _GEN_52; // @[sequencer-master.scala 362:41]
  wire  _GEN_1053 = io_op_bits_base_vd_valid ? _GEN_1005 : _GEN_53; // @[sequencer-master.scala 362:41]
  wire  _GEN_1054 = io_op_bits_base_vd_valid ? _GEN_1006 : _GEN_54; // @[sequencer-master.scala 362:41]
  wire  _GEN_1055 = io_op_bits_base_vd_valid ? _GEN_1007 : _GEN_55; // @[sequencer-master.scala 362:41]
  wire  _GEN_1056 = io_op_bits_base_vd_valid ? _GEN_1008 : e_0_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1057 = io_op_bits_base_vd_valid ? _GEN_1009 : e_1_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1058 = io_op_bits_base_vd_valid ? _GEN_1010 : e_2_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1059 = io_op_bits_base_vd_valid ? _GEN_1011 : e_3_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1060 = io_op_bits_base_vd_valid ? _GEN_1012 : e_4_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1061 = io_op_bits_base_vd_valid ? _GEN_1013 : e_5_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1062 = io_op_bits_base_vd_valid ? _GEN_1014 : e_6_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1063 = io_op_bits_base_vd_valid ? _GEN_1015 : e_7_base_vd_scalar; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1064 = io_op_bits_base_vd_valid ? _GEN_1016 : e_0_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1065 = io_op_bits_base_vd_valid ? _GEN_1017 : e_1_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1066 = io_op_bits_base_vd_valid ? _GEN_1018 : e_2_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1067 = io_op_bits_base_vd_valid ? _GEN_1019 : e_3_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1068 = io_op_bits_base_vd_valid ? _GEN_1020 : e_4_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1069 = io_op_bits_base_vd_valid ? _GEN_1021 : e_5_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1070 = io_op_bits_base_vd_valid ? _GEN_1022 : e_6_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire  _GEN_1071 = io_op_bits_base_vd_valid ? _GEN_1023 : e_7_base_vd_pred; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1072 = io_op_bits_base_vd_valid ? _GEN_1024 : e_0_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1073 = io_op_bits_base_vd_valid ? _GEN_1025 : e_1_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1074 = io_op_bits_base_vd_valid ? _GEN_1026 : e_2_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1075 = io_op_bits_base_vd_valid ? _GEN_1027 : e_3_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1076 = io_op_bits_base_vd_valid ? _GEN_1028 : e_4_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1077 = io_op_bits_base_vd_valid ? _GEN_1029 : e_5_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1078 = io_op_bits_base_vd_valid ? _GEN_1030 : e_6_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1079 = io_op_bits_base_vd_valid ? _GEN_1031 : e_7_base_vd_prec; // @[sequencer-master.scala 362:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1080 = io_op_bits_base_vd_valid ? _GEN_1032 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1081 = io_op_bits_base_vd_valid ? _GEN_1033 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1082 = io_op_bits_base_vd_valid ? _GEN_1034 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1083 = io_op_bits_base_vd_valid ? _GEN_1035 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1084 = io_op_bits_base_vd_valid ? _GEN_1036 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1085 = io_op_bits_base_vd_valid ? _GEN_1037 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1086 = io_op_bits_base_vd_valid ? _GEN_1038 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1087 = io_op_bits_base_vd_valid ? _GEN_1039 : 8'h0; // @[sequencer-master.scala 362:41 sequencer-master.scala 411:33]
  wire  _GEN_1088 = _GEN_32729 | _GEN_72; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1089 = _GEN_32730 | _GEN_73; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1090 = _GEN_32731 | _GEN_74; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1091 = _GEN_32732 | _GEN_75; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1092 = _GEN_32733 | _GEN_76; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1093 = _GEN_32734 | _GEN_77; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1094 = _GEN_32735 | _GEN_78; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1095 = _GEN_32736 | _GEN_79; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1096 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1088 : _GEN_72; // @[sequencer-master.scala 161:86]
  wire  _GEN_1097 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1089 : _GEN_73; // @[sequencer-master.scala 161:86]
  wire  _GEN_1098 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1090 : _GEN_74; // @[sequencer-master.scala 161:86]
  wire  _GEN_1099 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1091 : _GEN_75; // @[sequencer-master.scala 161:86]
  wire  _GEN_1100 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1092 : _GEN_76; // @[sequencer-master.scala 161:86]
  wire  _GEN_1101 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1093 : _GEN_77; // @[sequencer-master.scala 161:86]
  wire  _GEN_1102 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1094 : _GEN_78; // @[sequencer-master.scala 161:86]
  wire  _GEN_1103 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_1095 : _GEN_79; // @[sequencer-master.scala 161:86]
  wire  _GEN_1104 = _GEN_32729 | _GEN_96; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1105 = _GEN_32730 | _GEN_97; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1106 = _GEN_32731 | _GEN_98; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1107 = _GEN_32732 | _GEN_99; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1108 = _GEN_32733 | _GEN_100; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1109 = _GEN_32734 | _GEN_101; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1110 = _GEN_32735 | _GEN_102; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1111 = _GEN_32736 | _GEN_103; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1112 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1104 : _GEN_96; // @[sequencer-master.scala 161:86]
  wire  _GEN_1113 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1105 : _GEN_97; // @[sequencer-master.scala 161:86]
  wire  _GEN_1114 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1106 : _GEN_98; // @[sequencer-master.scala 161:86]
  wire  _GEN_1115 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1107 : _GEN_99; // @[sequencer-master.scala 161:86]
  wire  _GEN_1116 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1108 : _GEN_100; // @[sequencer-master.scala 161:86]
  wire  _GEN_1117 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1109 : _GEN_101; // @[sequencer-master.scala 161:86]
  wire  _GEN_1118 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1110 : _GEN_102; // @[sequencer-master.scala 161:86]
  wire  _GEN_1119 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_1111 : _GEN_103; // @[sequencer-master.scala 161:86]
  wire  _GEN_1120 = _GEN_32729 | _GEN_120; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1121 = _GEN_32730 | _GEN_121; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1122 = _GEN_32731 | _GEN_122; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1123 = _GEN_32732 | _GEN_123; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1124 = _GEN_32733 | _GEN_124; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1125 = _GEN_32734 | _GEN_125; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1126 = _GEN_32735 | _GEN_126; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1127 = _GEN_32736 | _GEN_127; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1128 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1120 : _GEN_120; // @[sequencer-master.scala 161:86]
  wire  _GEN_1129 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1121 : _GEN_121; // @[sequencer-master.scala 161:86]
  wire  _GEN_1130 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1122 : _GEN_122; // @[sequencer-master.scala 161:86]
  wire  _GEN_1131 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1123 : _GEN_123; // @[sequencer-master.scala 161:86]
  wire  _GEN_1132 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1124 : _GEN_124; // @[sequencer-master.scala 161:86]
  wire  _GEN_1133 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1125 : _GEN_125; // @[sequencer-master.scala 161:86]
  wire  _GEN_1134 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1126 : _GEN_126; // @[sequencer-master.scala 161:86]
  wire  _GEN_1135 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_1127 : _GEN_127; // @[sequencer-master.scala 161:86]
  wire  _GEN_1136 = _GEN_32729 | _GEN_144; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1137 = _GEN_32730 | _GEN_145; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1138 = _GEN_32731 | _GEN_146; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1139 = _GEN_32732 | _GEN_147; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1140 = _GEN_32733 | _GEN_148; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1141 = _GEN_32734 | _GEN_149; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1142 = _GEN_32735 | _GEN_150; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1143 = _GEN_32736 | _GEN_151; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1144 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1136 : _GEN_144; // @[sequencer-master.scala 161:86]
  wire  _GEN_1145 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1137 : _GEN_145; // @[sequencer-master.scala 161:86]
  wire  _GEN_1146 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1138 : _GEN_146; // @[sequencer-master.scala 161:86]
  wire  _GEN_1147 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1139 : _GEN_147; // @[sequencer-master.scala 161:86]
  wire  _GEN_1148 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1140 : _GEN_148; // @[sequencer-master.scala 161:86]
  wire  _GEN_1149 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1141 : _GEN_149; // @[sequencer-master.scala 161:86]
  wire  _GEN_1150 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1142 : _GEN_150; // @[sequencer-master.scala 161:86]
  wire  _GEN_1151 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_1143 : _GEN_151; // @[sequencer-master.scala 161:86]
  wire  _GEN_1152 = _GEN_32729 | _GEN_168; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1153 = _GEN_32730 | _GEN_169; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1154 = _GEN_32731 | _GEN_170; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1155 = _GEN_32732 | _GEN_171; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1156 = _GEN_32733 | _GEN_172; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1157 = _GEN_32734 | _GEN_173; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1158 = _GEN_32735 | _GEN_174; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1159 = _GEN_32736 | _GEN_175; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1160 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1152 : _GEN_168; // @[sequencer-master.scala 161:86]
  wire  _GEN_1161 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1153 : _GEN_169; // @[sequencer-master.scala 161:86]
  wire  _GEN_1162 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1154 : _GEN_170; // @[sequencer-master.scala 161:86]
  wire  _GEN_1163 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1155 : _GEN_171; // @[sequencer-master.scala 161:86]
  wire  _GEN_1164 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1156 : _GEN_172; // @[sequencer-master.scala 161:86]
  wire  _GEN_1165 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1157 : _GEN_173; // @[sequencer-master.scala 161:86]
  wire  _GEN_1166 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1158 : _GEN_174; // @[sequencer-master.scala 161:86]
  wire  _GEN_1167 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_1159 : _GEN_175; // @[sequencer-master.scala 161:86]
  wire  _GEN_1168 = _GEN_32729 | _GEN_192; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1169 = _GEN_32730 | _GEN_193; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1170 = _GEN_32731 | _GEN_194; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1171 = _GEN_32732 | _GEN_195; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1172 = _GEN_32733 | _GEN_196; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1173 = _GEN_32734 | _GEN_197; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1174 = _GEN_32735 | _GEN_198; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1175 = _GEN_32736 | _GEN_199; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1176 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1168 : _GEN_192; // @[sequencer-master.scala 161:86]
  wire  _GEN_1177 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1169 : _GEN_193; // @[sequencer-master.scala 161:86]
  wire  _GEN_1178 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1170 : _GEN_194; // @[sequencer-master.scala 161:86]
  wire  _GEN_1179 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1171 : _GEN_195; // @[sequencer-master.scala 161:86]
  wire  _GEN_1180 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1172 : _GEN_196; // @[sequencer-master.scala 161:86]
  wire  _GEN_1181 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1173 : _GEN_197; // @[sequencer-master.scala 161:86]
  wire  _GEN_1182 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1174 : _GEN_198; // @[sequencer-master.scala 161:86]
  wire  _GEN_1183 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_1175 : _GEN_199; // @[sequencer-master.scala 161:86]
  wire  _GEN_1184 = _GEN_32729 | _GEN_216; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1185 = _GEN_32730 | _GEN_217; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1186 = _GEN_32731 | _GEN_218; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1187 = _GEN_32732 | _GEN_219; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1188 = _GEN_32733 | _GEN_220; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1189 = _GEN_32734 | _GEN_221; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1190 = _GEN_32735 | _GEN_222; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1191 = _GEN_32736 | _GEN_223; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1192 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1184 : _GEN_216; // @[sequencer-master.scala 161:86]
  wire  _GEN_1193 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1185 : _GEN_217; // @[sequencer-master.scala 161:86]
  wire  _GEN_1194 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1186 : _GEN_218; // @[sequencer-master.scala 161:86]
  wire  _GEN_1195 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1187 : _GEN_219; // @[sequencer-master.scala 161:86]
  wire  _GEN_1196 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1188 : _GEN_220; // @[sequencer-master.scala 161:86]
  wire  _GEN_1197 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1189 : _GEN_221; // @[sequencer-master.scala 161:86]
  wire  _GEN_1198 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1190 : _GEN_222; // @[sequencer-master.scala 161:86]
  wire  _GEN_1199 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_1191 : _GEN_223; // @[sequencer-master.scala 161:86]
  wire  _GEN_1200 = _GEN_32729 | _GEN_240; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1201 = _GEN_32730 | _GEN_241; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1202 = _GEN_32731 | _GEN_242; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1203 = _GEN_32732 | _GEN_243; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1204 = _GEN_32733 | _GEN_244; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1205 = _GEN_32734 | _GEN_245; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1206 = _GEN_32735 | _GEN_246; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1207 = _GEN_32736 | _GEN_247; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_1208 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1200 : _GEN_240; // @[sequencer-master.scala 161:86]
  wire  _GEN_1209 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1201 : _GEN_241; // @[sequencer-master.scala 161:86]
  wire  _GEN_1210 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1202 : _GEN_242; // @[sequencer-master.scala 161:86]
  wire  _GEN_1211 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1203 : _GEN_243; // @[sequencer-master.scala 161:86]
  wire  _GEN_1212 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1204 : _GEN_244; // @[sequencer-master.scala 161:86]
  wire  _GEN_1213 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1205 : _GEN_245; // @[sequencer-master.scala 161:86]
  wire  _GEN_1214 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1206 : _GEN_246; // @[sequencer-master.scala 161:86]
  wire  _GEN_1215 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_1207 : _GEN_247; // @[sequencer-master.scala 161:86]
  wire  _GEN_1216 = _GEN_32729 | _GEN_80; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1217 = _GEN_32730 | _GEN_81; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1218 = _GEN_32731 | _GEN_82; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1219 = _GEN_32732 | _GEN_83; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1220 = _GEN_32733 | _GEN_84; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1221 = _GEN_32734 | _GEN_85; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1222 = _GEN_32735 | _GEN_86; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1223 = _GEN_32736 | _GEN_87; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1224 = _T_1442 ? _GEN_1216 : _GEN_80; // @[sequencer-master.scala 168:32]
  wire  _GEN_1225 = _T_1442 ? _GEN_1217 : _GEN_81; // @[sequencer-master.scala 168:32]
  wire  _GEN_1226 = _T_1442 ? _GEN_1218 : _GEN_82; // @[sequencer-master.scala 168:32]
  wire  _GEN_1227 = _T_1442 ? _GEN_1219 : _GEN_83; // @[sequencer-master.scala 168:32]
  wire  _GEN_1228 = _T_1442 ? _GEN_1220 : _GEN_84; // @[sequencer-master.scala 168:32]
  wire  _GEN_1229 = _T_1442 ? _GEN_1221 : _GEN_85; // @[sequencer-master.scala 168:32]
  wire  _GEN_1230 = _T_1442 ? _GEN_1222 : _GEN_86; // @[sequencer-master.scala 168:32]
  wire  _GEN_1231 = _T_1442 ? _GEN_1223 : _GEN_87; // @[sequencer-master.scala 168:32]
  wire  _GEN_1232 = _GEN_32729 | _GEN_104; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1233 = _GEN_32730 | _GEN_105; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1234 = _GEN_32731 | _GEN_106; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1235 = _GEN_32732 | _GEN_107; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1236 = _GEN_32733 | _GEN_108; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1237 = _GEN_32734 | _GEN_109; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1238 = _GEN_32735 | _GEN_110; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1239 = _GEN_32736 | _GEN_111; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1240 = _T_1464 ? _GEN_1232 : _GEN_104; // @[sequencer-master.scala 168:32]
  wire  _GEN_1241 = _T_1464 ? _GEN_1233 : _GEN_105; // @[sequencer-master.scala 168:32]
  wire  _GEN_1242 = _T_1464 ? _GEN_1234 : _GEN_106; // @[sequencer-master.scala 168:32]
  wire  _GEN_1243 = _T_1464 ? _GEN_1235 : _GEN_107; // @[sequencer-master.scala 168:32]
  wire  _GEN_1244 = _T_1464 ? _GEN_1236 : _GEN_108; // @[sequencer-master.scala 168:32]
  wire  _GEN_1245 = _T_1464 ? _GEN_1237 : _GEN_109; // @[sequencer-master.scala 168:32]
  wire  _GEN_1246 = _T_1464 ? _GEN_1238 : _GEN_110; // @[sequencer-master.scala 168:32]
  wire  _GEN_1247 = _T_1464 ? _GEN_1239 : _GEN_111; // @[sequencer-master.scala 168:32]
  wire  _GEN_1248 = _GEN_32729 | _GEN_128; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1249 = _GEN_32730 | _GEN_129; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1250 = _GEN_32731 | _GEN_130; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1251 = _GEN_32732 | _GEN_131; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1252 = _GEN_32733 | _GEN_132; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1253 = _GEN_32734 | _GEN_133; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1254 = _GEN_32735 | _GEN_134; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1255 = _GEN_32736 | _GEN_135; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1256 = _T_1486 ? _GEN_1248 : _GEN_128; // @[sequencer-master.scala 168:32]
  wire  _GEN_1257 = _T_1486 ? _GEN_1249 : _GEN_129; // @[sequencer-master.scala 168:32]
  wire  _GEN_1258 = _T_1486 ? _GEN_1250 : _GEN_130; // @[sequencer-master.scala 168:32]
  wire  _GEN_1259 = _T_1486 ? _GEN_1251 : _GEN_131; // @[sequencer-master.scala 168:32]
  wire  _GEN_1260 = _T_1486 ? _GEN_1252 : _GEN_132; // @[sequencer-master.scala 168:32]
  wire  _GEN_1261 = _T_1486 ? _GEN_1253 : _GEN_133; // @[sequencer-master.scala 168:32]
  wire  _GEN_1262 = _T_1486 ? _GEN_1254 : _GEN_134; // @[sequencer-master.scala 168:32]
  wire  _GEN_1263 = _T_1486 ? _GEN_1255 : _GEN_135; // @[sequencer-master.scala 168:32]
  wire  _GEN_1264 = _GEN_32729 | _GEN_152; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1265 = _GEN_32730 | _GEN_153; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1266 = _GEN_32731 | _GEN_154; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1267 = _GEN_32732 | _GEN_155; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1268 = _GEN_32733 | _GEN_156; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1269 = _GEN_32734 | _GEN_157; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1270 = _GEN_32735 | _GEN_158; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1271 = _GEN_32736 | _GEN_159; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1272 = _T_1508 ? _GEN_1264 : _GEN_152; // @[sequencer-master.scala 168:32]
  wire  _GEN_1273 = _T_1508 ? _GEN_1265 : _GEN_153; // @[sequencer-master.scala 168:32]
  wire  _GEN_1274 = _T_1508 ? _GEN_1266 : _GEN_154; // @[sequencer-master.scala 168:32]
  wire  _GEN_1275 = _T_1508 ? _GEN_1267 : _GEN_155; // @[sequencer-master.scala 168:32]
  wire  _GEN_1276 = _T_1508 ? _GEN_1268 : _GEN_156; // @[sequencer-master.scala 168:32]
  wire  _GEN_1277 = _T_1508 ? _GEN_1269 : _GEN_157; // @[sequencer-master.scala 168:32]
  wire  _GEN_1278 = _T_1508 ? _GEN_1270 : _GEN_158; // @[sequencer-master.scala 168:32]
  wire  _GEN_1279 = _T_1508 ? _GEN_1271 : _GEN_159; // @[sequencer-master.scala 168:32]
  wire  _GEN_1280 = _GEN_32729 | _GEN_176; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1281 = _GEN_32730 | _GEN_177; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1282 = _GEN_32731 | _GEN_178; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1283 = _GEN_32732 | _GEN_179; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1284 = _GEN_32733 | _GEN_180; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1285 = _GEN_32734 | _GEN_181; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1286 = _GEN_32735 | _GEN_182; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1287 = _GEN_32736 | _GEN_183; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1288 = _T_1530 ? _GEN_1280 : _GEN_176; // @[sequencer-master.scala 168:32]
  wire  _GEN_1289 = _T_1530 ? _GEN_1281 : _GEN_177; // @[sequencer-master.scala 168:32]
  wire  _GEN_1290 = _T_1530 ? _GEN_1282 : _GEN_178; // @[sequencer-master.scala 168:32]
  wire  _GEN_1291 = _T_1530 ? _GEN_1283 : _GEN_179; // @[sequencer-master.scala 168:32]
  wire  _GEN_1292 = _T_1530 ? _GEN_1284 : _GEN_180; // @[sequencer-master.scala 168:32]
  wire  _GEN_1293 = _T_1530 ? _GEN_1285 : _GEN_181; // @[sequencer-master.scala 168:32]
  wire  _GEN_1294 = _T_1530 ? _GEN_1286 : _GEN_182; // @[sequencer-master.scala 168:32]
  wire  _GEN_1295 = _T_1530 ? _GEN_1287 : _GEN_183; // @[sequencer-master.scala 168:32]
  wire  _GEN_1296 = _GEN_32729 | _GEN_200; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1297 = _GEN_32730 | _GEN_201; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1298 = _GEN_32731 | _GEN_202; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1299 = _GEN_32732 | _GEN_203; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1300 = _GEN_32733 | _GEN_204; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1301 = _GEN_32734 | _GEN_205; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1302 = _GEN_32735 | _GEN_206; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1303 = _GEN_32736 | _GEN_207; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1304 = _T_1552 ? _GEN_1296 : _GEN_200; // @[sequencer-master.scala 168:32]
  wire  _GEN_1305 = _T_1552 ? _GEN_1297 : _GEN_201; // @[sequencer-master.scala 168:32]
  wire  _GEN_1306 = _T_1552 ? _GEN_1298 : _GEN_202; // @[sequencer-master.scala 168:32]
  wire  _GEN_1307 = _T_1552 ? _GEN_1299 : _GEN_203; // @[sequencer-master.scala 168:32]
  wire  _GEN_1308 = _T_1552 ? _GEN_1300 : _GEN_204; // @[sequencer-master.scala 168:32]
  wire  _GEN_1309 = _T_1552 ? _GEN_1301 : _GEN_205; // @[sequencer-master.scala 168:32]
  wire  _GEN_1310 = _T_1552 ? _GEN_1302 : _GEN_206; // @[sequencer-master.scala 168:32]
  wire  _GEN_1311 = _T_1552 ? _GEN_1303 : _GEN_207; // @[sequencer-master.scala 168:32]
  wire  _GEN_1312 = _GEN_32729 | _GEN_224; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1313 = _GEN_32730 | _GEN_225; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1314 = _GEN_32731 | _GEN_226; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1315 = _GEN_32732 | _GEN_227; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1316 = _GEN_32733 | _GEN_228; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1317 = _GEN_32734 | _GEN_229; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1318 = _GEN_32735 | _GEN_230; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1319 = _GEN_32736 | _GEN_231; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1320 = _T_1574 ? _GEN_1312 : _GEN_224; // @[sequencer-master.scala 168:32]
  wire  _GEN_1321 = _T_1574 ? _GEN_1313 : _GEN_225; // @[sequencer-master.scala 168:32]
  wire  _GEN_1322 = _T_1574 ? _GEN_1314 : _GEN_226; // @[sequencer-master.scala 168:32]
  wire  _GEN_1323 = _T_1574 ? _GEN_1315 : _GEN_227; // @[sequencer-master.scala 168:32]
  wire  _GEN_1324 = _T_1574 ? _GEN_1316 : _GEN_228; // @[sequencer-master.scala 168:32]
  wire  _GEN_1325 = _T_1574 ? _GEN_1317 : _GEN_229; // @[sequencer-master.scala 168:32]
  wire  _GEN_1326 = _T_1574 ? _GEN_1318 : _GEN_230; // @[sequencer-master.scala 168:32]
  wire  _GEN_1327 = _T_1574 ? _GEN_1319 : _GEN_231; // @[sequencer-master.scala 168:32]
  wire  _GEN_1328 = _GEN_32729 | _GEN_248; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1329 = _GEN_32730 | _GEN_249; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1330 = _GEN_32731 | _GEN_250; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1331 = _GEN_32732 | _GEN_251; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1332 = _GEN_32733 | _GEN_252; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1333 = _GEN_32734 | _GEN_253; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1334 = _GEN_32735 | _GEN_254; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1335 = _GEN_32736 | _GEN_255; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_1336 = _T_1596 ? _GEN_1328 : _GEN_248; // @[sequencer-master.scala 168:32]
  wire  _GEN_1337 = _T_1596 ? _GEN_1329 : _GEN_249; // @[sequencer-master.scala 168:32]
  wire  _GEN_1338 = _T_1596 ? _GEN_1330 : _GEN_250; // @[sequencer-master.scala 168:32]
  wire  _GEN_1339 = _T_1596 ? _GEN_1331 : _GEN_251; // @[sequencer-master.scala 168:32]
  wire  _GEN_1340 = _T_1596 ? _GEN_1332 : _GEN_252; // @[sequencer-master.scala 168:32]
  wire  _GEN_1341 = _T_1596 ? _GEN_1333 : _GEN_253; // @[sequencer-master.scala 168:32]
  wire  _GEN_1342 = _T_1596 ? _GEN_1334 : _GEN_254; // @[sequencer-master.scala 168:32]
  wire  _GEN_1343 = _T_1596 ? _GEN_1335 : _GEN_255; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_1344 = 3'h0 == tail ? _T_1615[1:0] : e_0_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1345 = 3'h1 == tail ? _T_1615[1:0] : e_1_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1346 = 3'h2 == tail ? _T_1615[1:0] : e_2_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1347 = 3'h3 == tail ? _T_1615[1:0] : e_3_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1348 = 3'h4 == tail ? _T_1615[1:0] : e_4_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1349 = 3'h5 == tail ? _T_1615[1:0] : e_5_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1350 = 3'h6 == tail ? _T_1615[1:0] : e_6_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1351 = 3'h7 == tail ? _T_1615[1:0] : e_7_rports; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1352 = 3'h0 == tail ? 4'h0 : e_0_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1353 = 3'h1 == tail ? 4'h0 : e_1_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1354 = 3'h2 == tail ? 4'h0 : e_2_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1355 = 3'h3 == tail ? 4'h0 : e_3_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1356 = 3'h4 == tail ? 4'h0 : e_4_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1357 = 3'h5 == tail ? 4'h0 : e_5_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1358 = 3'h6 == tail ? 4'h0 : e_6_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1359 = 3'h7 == tail ? 4'h0 : e_7_wport_sram; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1360 = 3'h0 == tail ? 3'h0 : e_0_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1361 = 3'h1 == tail ? 3'h0 : e_1_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1362 = 3'h2 == tail ? 3'h0 : e_2_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1363 = 3'h3 == tail ? 3'h0 : e_3_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1364 = 3'h4 == tail ? 3'h0 : e_4_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1365 = 3'h5 == tail ? 3'h0 : e_5_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1366 = 3'h6 == tail ? 3'h0 : e_6_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1367 = 3'h7 == tail ? 3'h0 : e_7_wport_pred; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25 sequencer-master.scala 109:14]
  wire [4:0] _T_1789 = {{2'd0}, _T_1615}; // @[sequencer-master.scala 247:46]
  wire [3:0] _T_1792 = _T_1789[3:0] + 4'h2; // @[sequencer-master.scala 247:56]
  wire [3:0] _GEN_1368 = 3'h0 == tail ? _T_1792 : _GEN_1352; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1369 = 3'h1 == tail ? _T_1792 : _GEN_1353; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1370 = 3'h2 == tail ? _T_1792 : _GEN_1354; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1371 = 3'h3 == tail ? _T_1792 : _GEN_1355; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1372 = 3'h4 == tail ? _T_1792 : _GEN_1356; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1373 = 3'h5 == tail ? _T_1792 : _GEN_1357; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1374 = 3'h6 == tail ? _T_1792 : _GEN_1358; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1375 = 3'h7 == tail ? _T_1792 : _GEN_1359; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_1376 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1368 : _GEN_1352; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1377 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1369 : _GEN_1353; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1378 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1370 : _GEN_1354; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1379 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1371 : _GEN_1355; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1380 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1372 : _GEN_1356; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1381 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1373 : _GEN_1357; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1382 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1374 : _GEN_1358; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_1383 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_1375 : _GEN_1359; // @[sequencer-master.scala 235:47]
  wire [2:0] _GEN_1384 = 3'h0 == tail ? _T_1792[2:0] : _GEN_1360; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1385 = 3'h1 == tail ? _T_1792[2:0] : _GEN_1361; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1386 = 3'h2 == tail ? _T_1792[2:0] : _GEN_1362; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1387 = 3'h3 == tail ? _T_1792[2:0] : _GEN_1363; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1388 = 3'h4 == tail ? _T_1792[2:0] : _GEN_1364; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1389 = 3'h5 == tail ? _T_1792[2:0] : _GEN_1365; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1390 = 3'h6 == tail ? _T_1792[2:0] : _GEN_1366; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1391 = 3'h7 == tail ? _T_1792[2:0] : _GEN_1367; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_1392 = io_op_bits_base_vd_pred ? _GEN_1384 : _GEN_1360; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1393 = io_op_bits_base_vd_pred ? _GEN_1385 : _GEN_1361; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1394 = io_op_bits_base_vd_pred ? _GEN_1386 : _GEN_1362; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1395 = io_op_bits_base_vd_pred ? _GEN_1387 : _GEN_1363; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1396 = io_op_bits_base_vd_pred ? _GEN_1388 : _GEN_1364; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1397 = io_op_bits_base_vd_pred ? _GEN_1389 : _GEN_1365; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1398 = io_op_bits_base_vd_pred ? _GEN_1390 : _GEN_1366; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_1399 = io_op_bits_base_vd_pred ? _GEN_1391 : _GEN_1367; // @[sequencer-master.scala 236:45]
  wire  _GEN_1400 = io_op_bits_active_vint ? _GEN_0 : v_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1401 = io_op_bits_active_vint ? _GEN_1 : v_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1402 = io_op_bits_active_vint ? _GEN_2 : v_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1403 = io_op_bits_active_vint ? _GEN_3 : v_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1404 = io_op_bits_active_vint ? _GEN_4 : v_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1405 = io_op_bits_active_vint ? _GEN_5 : v_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1406 = io_op_bits_active_vint ? _GEN_6 : v_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1407 = io_op_bits_active_vint ? _GEN_7 : v_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 107:14]
  wire  _GEN_1416 = io_op_bits_active_vint ? _GEN_336 : e_0_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1417 = io_op_bits_active_vint ? _GEN_337 : e_1_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1418 = io_op_bits_active_vint ? _GEN_338 : e_2_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1419 = io_op_bits_active_vint ? _GEN_339 : e_3_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1420 = io_op_bits_active_vint ? _GEN_340 : e_4_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1421 = io_op_bits_active_vint ? _GEN_341 : e_5_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1422 = io_op_bits_active_vint ? _GEN_342 : e_6_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1423 = io_op_bits_active_vint ? _GEN_343 : e_7_base_vp_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1424 = io_op_bits_active_vint ? _GEN_568 : e_0_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1425 = io_op_bits_active_vint ? _GEN_569 : e_1_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1426 = io_op_bits_active_vint ? _GEN_570 : e_2_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1427 = io_op_bits_active_vint ? _GEN_571 : e_3_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1428 = io_op_bits_active_vint ? _GEN_572 : e_4_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1429 = io_op_bits_active_vint ? _GEN_573 : e_5_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1430 = io_op_bits_active_vint ? _GEN_574 : e_6_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1431 = io_op_bits_active_vint ? _GEN_575 : e_7_base_vs1_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1432 = io_op_bits_active_vint ? _GEN_816 : e_0_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1433 = io_op_bits_active_vint ? _GEN_817 : e_1_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1434 = io_op_bits_active_vint ? _GEN_818 : e_2_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1435 = io_op_bits_active_vint ? _GEN_819 : e_3_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1436 = io_op_bits_active_vint ? _GEN_820 : e_4_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1437 = io_op_bits_active_vint ? _GEN_821 : e_5_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1438 = io_op_bits_active_vint ? _GEN_822 : e_6_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1439 = io_op_bits_active_vint ? _GEN_823 : e_7_base_vs2_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1440 = io_op_bits_active_vint ? _GEN_40 : e_0_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1441 = io_op_bits_active_vint ? _GEN_41 : e_1_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1442 = io_op_bits_active_vint ? _GEN_42 : e_2_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1443 = io_op_bits_active_vint ? _GEN_43 : e_3_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1444 = io_op_bits_active_vint ? _GEN_44 : e_4_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1445 = io_op_bits_active_vint ? _GEN_45 : e_5_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1446 = io_op_bits_active_vint ? _GEN_46 : e_6_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1447 = io_op_bits_active_vint ? _GEN_47 : e_7_base_vs3_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1448 = io_op_bits_active_vint ? _GEN_1048 : e_0_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1449 = io_op_bits_active_vint ? _GEN_1049 : e_1_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1450 = io_op_bits_active_vint ? _GEN_1050 : e_2_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1451 = io_op_bits_active_vint ? _GEN_1051 : e_3_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1452 = io_op_bits_active_vint ? _GEN_1052 : e_4_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1453 = io_op_bits_active_vint ? _GEN_1053 : e_5_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1454 = io_op_bits_active_vint ? _GEN_1054 : e_6_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1455 = io_op_bits_active_vint ? _GEN_1055 : e_7_base_vd_valid; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1456 = io_op_bits_active_vint & _GEN_32729; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1457 = io_op_bits_active_vint & _GEN_32730; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1458 = io_op_bits_active_vint & _GEN_32731; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1459 = io_op_bits_active_vint & _GEN_32732; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1460 = io_op_bits_active_vint & _GEN_32733; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1461 = io_op_bits_active_vint & _GEN_32734; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1462 = io_op_bits_active_vint & _GEN_32735; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1463 = io_op_bits_active_vint & _GEN_32736; // @[sequencer-master.scala 640:39 sequencer-master.scala 192:24]
  wire  _GEN_1464 = io_op_bits_active_vint ? _GEN_872 : e_0_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1465 = io_op_bits_active_vint ? _GEN_873 : e_1_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1466 = io_op_bits_active_vint ? _GEN_874 : e_2_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1467 = io_op_bits_active_vint ? _GEN_875 : e_3_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1468 = io_op_bits_active_vint ? _GEN_876 : e_4_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1469 = io_op_bits_active_vint ? _GEN_877 : e_5_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1470 = io_op_bits_active_vint ? _GEN_878 : e_6_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1471 = io_op_bits_active_vint ? _GEN_879 : e_7_raw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1472 = io_op_bits_active_vint ? _GEN_1096 : e_0_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1473 = io_op_bits_active_vint ? _GEN_1097 : e_1_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1474 = io_op_bits_active_vint ? _GEN_1098 : e_2_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1475 = io_op_bits_active_vint ? _GEN_1099 : e_3_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1476 = io_op_bits_active_vint ? _GEN_1100 : e_4_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1477 = io_op_bits_active_vint ? _GEN_1101 : e_5_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1478 = io_op_bits_active_vint ? _GEN_1102 : e_6_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1479 = io_op_bits_active_vint ? _GEN_1103 : e_7_war_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1480 = io_op_bits_active_vint ? _GEN_1224 : e_0_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1481 = io_op_bits_active_vint ? _GEN_1225 : e_1_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1482 = io_op_bits_active_vint ? _GEN_1226 : e_2_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1483 = io_op_bits_active_vint ? _GEN_1227 : e_3_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1484 = io_op_bits_active_vint ? _GEN_1228 : e_4_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1485 = io_op_bits_active_vint ? _GEN_1229 : e_5_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1486 = io_op_bits_active_vint ? _GEN_1230 : e_6_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1487 = io_op_bits_active_vint ? _GEN_1231 : e_7_waw_0; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1488 = io_op_bits_active_vint ? _GEN_888 : e_0_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1489 = io_op_bits_active_vint ? _GEN_889 : e_1_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1490 = io_op_bits_active_vint ? _GEN_890 : e_2_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1491 = io_op_bits_active_vint ? _GEN_891 : e_3_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1492 = io_op_bits_active_vint ? _GEN_892 : e_4_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1493 = io_op_bits_active_vint ? _GEN_893 : e_5_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1494 = io_op_bits_active_vint ? _GEN_894 : e_6_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1495 = io_op_bits_active_vint ? _GEN_895 : e_7_raw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1496 = io_op_bits_active_vint ? _GEN_1112 : e_0_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1497 = io_op_bits_active_vint ? _GEN_1113 : e_1_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1498 = io_op_bits_active_vint ? _GEN_1114 : e_2_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1499 = io_op_bits_active_vint ? _GEN_1115 : e_3_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1500 = io_op_bits_active_vint ? _GEN_1116 : e_4_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1501 = io_op_bits_active_vint ? _GEN_1117 : e_5_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1502 = io_op_bits_active_vint ? _GEN_1118 : e_6_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1503 = io_op_bits_active_vint ? _GEN_1119 : e_7_war_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1504 = io_op_bits_active_vint ? _GEN_1240 : e_0_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1505 = io_op_bits_active_vint ? _GEN_1241 : e_1_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1506 = io_op_bits_active_vint ? _GEN_1242 : e_2_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1507 = io_op_bits_active_vint ? _GEN_1243 : e_3_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1508 = io_op_bits_active_vint ? _GEN_1244 : e_4_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1509 = io_op_bits_active_vint ? _GEN_1245 : e_5_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1510 = io_op_bits_active_vint ? _GEN_1246 : e_6_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1511 = io_op_bits_active_vint ? _GEN_1247 : e_7_waw_1; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1512 = io_op_bits_active_vint ? _GEN_904 : e_0_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1513 = io_op_bits_active_vint ? _GEN_905 : e_1_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1514 = io_op_bits_active_vint ? _GEN_906 : e_2_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1515 = io_op_bits_active_vint ? _GEN_907 : e_3_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1516 = io_op_bits_active_vint ? _GEN_908 : e_4_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1517 = io_op_bits_active_vint ? _GEN_909 : e_5_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1518 = io_op_bits_active_vint ? _GEN_910 : e_6_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1519 = io_op_bits_active_vint ? _GEN_911 : e_7_raw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1520 = io_op_bits_active_vint ? _GEN_1128 : e_0_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1521 = io_op_bits_active_vint ? _GEN_1129 : e_1_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1522 = io_op_bits_active_vint ? _GEN_1130 : e_2_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1523 = io_op_bits_active_vint ? _GEN_1131 : e_3_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1524 = io_op_bits_active_vint ? _GEN_1132 : e_4_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1525 = io_op_bits_active_vint ? _GEN_1133 : e_5_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1526 = io_op_bits_active_vint ? _GEN_1134 : e_6_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1527 = io_op_bits_active_vint ? _GEN_1135 : e_7_war_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1528 = io_op_bits_active_vint ? _GEN_1256 : e_0_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1529 = io_op_bits_active_vint ? _GEN_1257 : e_1_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1530 = io_op_bits_active_vint ? _GEN_1258 : e_2_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1531 = io_op_bits_active_vint ? _GEN_1259 : e_3_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1532 = io_op_bits_active_vint ? _GEN_1260 : e_4_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1533 = io_op_bits_active_vint ? _GEN_1261 : e_5_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1534 = io_op_bits_active_vint ? _GEN_1262 : e_6_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1535 = io_op_bits_active_vint ? _GEN_1263 : e_7_waw_2; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1536 = io_op_bits_active_vint ? _GEN_920 : e_0_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1537 = io_op_bits_active_vint ? _GEN_921 : e_1_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1538 = io_op_bits_active_vint ? _GEN_922 : e_2_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1539 = io_op_bits_active_vint ? _GEN_923 : e_3_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1540 = io_op_bits_active_vint ? _GEN_924 : e_4_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1541 = io_op_bits_active_vint ? _GEN_925 : e_5_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1542 = io_op_bits_active_vint ? _GEN_926 : e_6_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1543 = io_op_bits_active_vint ? _GEN_927 : e_7_raw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1544 = io_op_bits_active_vint ? _GEN_1144 : e_0_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1545 = io_op_bits_active_vint ? _GEN_1145 : e_1_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1546 = io_op_bits_active_vint ? _GEN_1146 : e_2_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1547 = io_op_bits_active_vint ? _GEN_1147 : e_3_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1548 = io_op_bits_active_vint ? _GEN_1148 : e_4_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1549 = io_op_bits_active_vint ? _GEN_1149 : e_5_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1550 = io_op_bits_active_vint ? _GEN_1150 : e_6_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1551 = io_op_bits_active_vint ? _GEN_1151 : e_7_war_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1552 = io_op_bits_active_vint ? _GEN_1272 : e_0_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1553 = io_op_bits_active_vint ? _GEN_1273 : e_1_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1554 = io_op_bits_active_vint ? _GEN_1274 : e_2_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1555 = io_op_bits_active_vint ? _GEN_1275 : e_3_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1556 = io_op_bits_active_vint ? _GEN_1276 : e_4_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1557 = io_op_bits_active_vint ? _GEN_1277 : e_5_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1558 = io_op_bits_active_vint ? _GEN_1278 : e_6_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1559 = io_op_bits_active_vint ? _GEN_1279 : e_7_waw_3; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1560 = io_op_bits_active_vint ? _GEN_936 : e_0_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1561 = io_op_bits_active_vint ? _GEN_937 : e_1_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1562 = io_op_bits_active_vint ? _GEN_938 : e_2_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1563 = io_op_bits_active_vint ? _GEN_939 : e_3_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1564 = io_op_bits_active_vint ? _GEN_940 : e_4_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1565 = io_op_bits_active_vint ? _GEN_941 : e_5_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1566 = io_op_bits_active_vint ? _GEN_942 : e_6_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1567 = io_op_bits_active_vint ? _GEN_943 : e_7_raw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1568 = io_op_bits_active_vint ? _GEN_1160 : e_0_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1569 = io_op_bits_active_vint ? _GEN_1161 : e_1_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1570 = io_op_bits_active_vint ? _GEN_1162 : e_2_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1571 = io_op_bits_active_vint ? _GEN_1163 : e_3_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1572 = io_op_bits_active_vint ? _GEN_1164 : e_4_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1573 = io_op_bits_active_vint ? _GEN_1165 : e_5_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1574 = io_op_bits_active_vint ? _GEN_1166 : e_6_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1575 = io_op_bits_active_vint ? _GEN_1167 : e_7_war_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1576 = io_op_bits_active_vint ? _GEN_1288 : e_0_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1577 = io_op_bits_active_vint ? _GEN_1289 : e_1_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1578 = io_op_bits_active_vint ? _GEN_1290 : e_2_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1579 = io_op_bits_active_vint ? _GEN_1291 : e_3_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1580 = io_op_bits_active_vint ? _GEN_1292 : e_4_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1581 = io_op_bits_active_vint ? _GEN_1293 : e_5_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1582 = io_op_bits_active_vint ? _GEN_1294 : e_6_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1583 = io_op_bits_active_vint ? _GEN_1295 : e_7_waw_4; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1584 = io_op_bits_active_vint ? _GEN_952 : e_0_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1585 = io_op_bits_active_vint ? _GEN_953 : e_1_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1586 = io_op_bits_active_vint ? _GEN_954 : e_2_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1587 = io_op_bits_active_vint ? _GEN_955 : e_3_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1588 = io_op_bits_active_vint ? _GEN_956 : e_4_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1589 = io_op_bits_active_vint ? _GEN_957 : e_5_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1590 = io_op_bits_active_vint ? _GEN_958 : e_6_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1591 = io_op_bits_active_vint ? _GEN_959 : e_7_raw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1592 = io_op_bits_active_vint ? _GEN_1176 : e_0_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1593 = io_op_bits_active_vint ? _GEN_1177 : e_1_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1594 = io_op_bits_active_vint ? _GEN_1178 : e_2_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1595 = io_op_bits_active_vint ? _GEN_1179 : e_3_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1596 = io_op_bits_active_vint ? _GEN_1180 : e_4_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1597 = io_op_bits_active_vint ? _GEN_1181 : e_5_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1598 = io_op_bits_active_vint ? _GEN_1182 : e_6_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1599 = io_op_bits_active_vint ? _GEN_1183 : e_7_war_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1600 = io_op_bits_active_vint ? _GEN_1304 : e_0_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1601 = io_op_bits_active_vint ? _GEN_1305 : e_1_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1602 = io_op_bits_active_vint ? _GEN_1306 : e_2_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1603 = io_op_bits_active_vint ? _GEN_1307 : e_3_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1604 = io_op_bits_active_vint ? _GEN_1308 : e_4_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1605 = io_op_bits_active_vint ? _GEN_1309 : e_5_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1606 = io_op_bits_active_vint ? _GEN_1310 : e_6_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1607 = io_op_bits_active_vint ? _GEN_1311 : e_7_waw_5; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1608 = io_op_bits_active_vint ? _GEN_968 : e_0_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1609 = io_op_bits_active_vint ? _GEN_969 : e_1_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1610 = io_op_bits_active_vint ? _GEN_970 : e_2_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1611 = io_op_bits_active_vint ? _GEN_971 : e_3_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1612 = io_op_bits_active_vint ? _GEN_972 : e_4_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1613 = io_op_bits_active_vint ? _GEN_973 : e_5_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1614 = io_op_bits_active_vint ? _GEN_974 : e_6_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1615 = io_op_bits_active_vint ? _GEN_975 : e_7_raw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1616 = io_op_bits_active_vint ? _GEN_1192 : e_0_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1617 = io_op_bits_active_vint ? _GEN_1193 : e_1_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1618 = io_op_bits_active_vint ? _GEN_1194 : e_2_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1619 = io_op_bits_active_vint ? _GEN_1195 : e_3_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1620 = io_op_bits_active_vint ? _GEN_1196 : e_4_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1621 = io_op_bits_active_vint ? _GEN_1197 : e_5_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1622 = io_op_bits_active_vint ? _GEN_1198 : e_6_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1623 = io_op_bits_active_vint ? _GEN_1199 : e_7_war_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1624 = io_op_bits_active_vint ? _GEN_1320 : e_0_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1625 = io_op_bits_active_vint ? _GEN_1321 : e_1_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1626 = io_op_bits_active_vint ? _GEN_1322 : e_2_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1627 = io_op_bits_active_vint ? _GEN_1323 : e_3_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1628 = io_op_bits_active_vint ? _GEN_1324 : e_4_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1629 = io_op_bits_active_vint ? _GEN_1325 : e_5_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1630 = io_op_bits_active_vint ? _GEN_1326 : e_6_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1631 = io_op_bits_active_vint ? _GEN_1327 : e_7_waw_6; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1632 = io_op_bits_active_vint ? _GEN_984 : e_0_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1633 = io_op_bits_active_vint ? _GEN_985 : e_1_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1634 = io_op_bits_active_vint ? _GEN_986 : e_2_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1635 = io_op_bits_active_vint ? _GEN_987 : e_3_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1636 = io_op_bits_active_vint ? _GEN_988 : e_4_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1637 = io_op_bits_active_vint ? _GEN_989 : e_5_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1638 = io_op_bits_active_vint ? _GEN_990 : e_6_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1639 = io_op_bits_active_vint ? _GEN_991 : e_7_raw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 194:26]
  wire  _GEN_1640 = io_op_bits_active_vint ? _GEN_1208 : e_0_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1641 = io_op_bits_active_vint ? _GEN_1209 : e_1_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1642 = io_op_bits_active_vint ? _GEN_1210 : e_2_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1643 = io_op_bits_active_vint ? _GEN_1211 : e_3_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1644 = io_op_bits_active_vint ? _GEN_1212 : e_4_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1645 = io_op_bits_active_vint ? _GEN_1213 : e_5_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1646 = io_op_bits_active_vint ? _GEN_1214 : e_6_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1647 = io_op_bits_active_vint ? _GEN_1215 : e_7_war_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 195:26]
  wire  _GEN_1648 = io_op_bits_active_vint ? _GEN_1336 : e_0_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1649 = io_op_bits_active_vint ? _GEN_1337 : e_1_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1650 = io_op_bits_active_vint ? _GEN_1338 : e_2_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1651 = io_op_bits_active_vint ? _GEN_1339 : e_3_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1652 = io_op_bits_active_vint ? _GEN_1340 : e_4_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1653 = io_op_bits_active_vint ? _GEN_1341 : e_5_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1654 = io_op_bits_active_vint ? _GEN_1342 : e_6_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1655 = io_op_bits_active_vint ? _GEN_1343 : e_7_waw_7; // @[sequencer-master.scala 640:39 sequencer-master.scala 196:26]
  wire  _GEN_1656 = io_op_bits_active_vint ? _GEN_256 : e_0_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1657 = io_op_bits_active_vint ? _GEN_257 : e_1_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1658 = io_op_bits_active_vint ? _GEN_258 : e_2_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1659 = io_op_bits_active_vint ? _GEN_259 : e_3_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1660 = io_op_bits_active_vint ? _GEN_260 : e_4_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1661 = io_op_bits_active_vint ? _GEN_261 : e_5_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1662 = io_op_bits_active_vint ? _GEN_262 : e_6_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1663 = io_op_bits_active_vint ? _GEN_263 : e_7_last; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1672 = io_op_bits_active_vint ? _GEN_272 : e_0_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1673 = io_op_bits_active_vint ? _GEN_273 : e_1_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1674 = io_op_bits_active_vint ? _GEN_274 : e_2_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1675 = io_op_bits_active_vint ? _GEN_275 : e_3_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1676 = io_op_bits_active_vint ? _GEN_276 : e_4_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1677 = io_op_bits_active_vint ? _GEN_277 : e_5_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1678 = io_op_bits_active_vint ? _GEN_278 : e_6_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1679 = io_op_bits_active_vint ? _GEN_279 : e_7_active_viu; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1680 = io_op_bits_active_vint ? _GEN_280 : e_0_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1681 = io_op_bits_active_vint ? _GEN_281 : e_1_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1682 = io_op_bits_active_vint ? _GEN_282 : e_2_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1683 = io_op_bits_active_vint ? _GEN_283 : e_3_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1684 = io_op_bits_active_vint ? _GEN_284 : e_4_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1685 = io_op_bits_active_vint ? _GEN_285 : e_5_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1686 = io_op_bits_active_vint ? _GEN_286 : e_6_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_1687 = io_op_bits_active_vint ? _GEN_287 : e_7_fn_union; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1688 = io_op_bits_active_vint ? _GEN_328 : e_0_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1689 = io_op_bits_active_vint ? _GEN_329 : e_1_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1690 = io_op_bits_active_vint ? _GEN_330 : e_2_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1691 = io_op_bits_active_vint ? _GEN_331 : e_3_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1692 = io_op_bits_active_vint ? _GEN_332 : e_4_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1693 = io_op_bits_active_vint ? _GEN_333 : e_5_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1694 = io_op_bits_active_vint ? _GEN_334 : e_6_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1695 = io_op_bits_active_vint ? _GEN_335 : e_7_base_vp_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1696 = io_op_bits_active_vint ? _GEN_344 : e_0_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1697 = io_op_bits_active_vint ? _GEN_345 : e_1_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1698 = io_op_bits_active_vint ? _GEN_346 : e_2_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1699 = io_op_bits_active_vint ? _GEN_347 : e_3_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1700 = io_op_bits_active_vint ? _GEN_348 : e_4_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1701 = io_op_bits_active_vint ? _GEN_349 : e_5_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1702 = io_op_bits_active_vint ? _GEN_350 : e_6_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1703 = io_op_bits_active_vint ? _GEN_351 : e_7_base_vp_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1704 = io_op_bits_active_vint ? _GEN_352 : e_0_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1705 = io_op_bits_active_vint ? _GEN_353 : e_1_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1706 = io_op_bits_active_vint ? _GEN_354 : e_2_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1707 = io_op_bits_active_vint ? _GEN_355 : e_3_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1708 = io_op_bits_active_vint ? _GEN_356 : e_4_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1709 = io_op_bits_active_vint ? _GEN_357 : e_5_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1710 = io_op_bits_active_vint ? _GEN_358 : e_6_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1711 = io_op_bits_active_vint ? _GEN_359 : e_7_base_vp_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1712 = io_op_bits_active_vint ? _GEN_360 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1713 = io_op_bits_active_vint ? _GEN_361 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1714 = io_op_bits_active_vint ? _GEN_362 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1715 = io_op_bits_active_vint ? _GEN_363 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1716 = io_op_bits_active_vint ? _GEN_364 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1717 = io_op_bits_active_vint ? _GEN_365 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1718 = io_op_bits_active_vint ? _GEN_366 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1719 = io_op_bits_active_vint ? _GEN_367 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1720 = io_op_bits_active_vint ? _GEN_560 : e_0_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1721 = io_op_bits_active_vint ? _GEN_561 : e_1_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1722 = io_op_bits_active_vint ? _GEN_562 : e_2_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1723 = io_op_bits_active_vint ? _GEN_563 : e_3_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1724 = io_op_bits_active_vint ? _GEN_564 : e_4_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1725 = io_op_bits_active_vint ? _GEN_565 : e_5_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1726 = io_op_bits_active_vint ? _GEN_566 : e_6_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1727 = io_op_bits_active_vint ? _GEN_567 : e_7_base_vs1_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1728 = io_op_bits_active_vint ? _GEN_576 : e_0_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1729 = io_op_bits_active_vint ? _GEN_577 : e_1_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1730 = io_op_bits_active_vint ? _GEN_578 : e_2_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1731 = io_op_bits_active_vint ? _GEN_579 : e_3_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1732 = io_op_bits_active_vint ? _GEN_580 : e_4_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1733 = io_op_bits_active_vint ? _GEN_581 : e_5_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1734 = io_op_bits_active_vint ? _GEN_582 : e_6_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1735 = io_op_bits_active_vint ? _GEN_583 : e_7_base_vs1_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1736 = io_op_bits_active_vint ? _GEN_584 : e_0_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1737 = io_op_bits_active_vint ? _GEN_585 : e_1_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1738 = io_op_bits_active_vint ? _GEN_586 : e_2_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1739 = io_op_bits_active_vint ? _GEN_587 : e_3_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1740 = io_op_bits_active_vint ? _GEN_588 : e_4_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1741 = io_op_bits_active_vint ? _GEN_589 : e_5_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1742 = io_op_bits_active_vint ? _GEN_590 : e_6_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1743 = io_op_bits_active_vint ? _GEN_591 : e_7_base_vs1_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1744 = io_op_bits_active_vint ? _GEN_592 : e_0_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1745 = io_op_bits_active_vint ? _GEN_593 : e_1_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1746 = io_op_bits_active_vint ? _GEN_594 : e_2_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1747 = io_op_bits_active_vint ? _GEN_595 : e_3_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1748 = io_op_bits_active_vint ? _GEN_596 : e_4_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1749 = io_op_bits_active_vint ? _GEN_597 : e_5_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1750 = io_op_bits_active_vint ? _GEN_598 : e_6_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1751 = io_op_bits_active_vint ? _GEN_599 : e_7_base_vs1_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1752 = io_op_bits_active_vint ? _GEN_600 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1753 = io_op_bits_active_vint ? _GEN_601 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1754 = io_op_bits_active_vint ? _GEN_602 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1755 = io_op_bits_active_vint ? _GEN_603 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1756 = io_op_bits_active_vint ? _GEN_604 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1757 = io_op_bits_active_vint ? _GEN_605 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1758 = io_op_bits_active_vint ? _GEN_606 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1759 = io_op_bits_active_vint ? _GEN_607 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [63:0] _GEN_1760 = io_op_bits_active_vint ? _GEN_608 : e_0_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1761 = io_op_bits_active_vint ? _GEN_609 : e_1_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1762 = io_op_bits_active_vint ? _GEN_610 : e_2_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1763 = io_op_bits_active_vint ? _GEN_611 : e_3_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1764 = io_op_bits_active_vint ? _GEN_612 : e_4_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1765 = io_op_bits_active_vint ? _GEN_613 : e_5_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1766 = io_op_bits_active_vint ? _GEN_614 : e_6_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1767 = io_op_bits_active_vint ? _GEN_615 : e_7_sreg_ss1; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1768 = io_op_bits_active_vint ? _GEN_808 : e_0_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1769 = io_op_bits_active_vint ? _GEN_809 : e_1_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1770 = io_op_bits_active_vint ? _GEN_810 : e_2_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1771 = io_op_bits_active_vint ? _GEN_811 : e_3_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1772 = io_op_bits_active_vint ? _GEN_812 : e_4_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1773 = io_op_bits_active_vint ? _GEN_813 : e_5_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1774 = io_op_bits_active_vint ? _GEN_814 : e_6_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1775 = io_op_bits_active_vint ? _GEN_815 : e_7_base_vs2_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1776 = io_op_bits_active_vint ? _GEN_824 : e_0_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1777 = io_op_bits_active_vint ? _GEN_825 : e_1_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1778 = io_op_bits_active_vint ? _GEN_826 : e_2_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1779 = io_op_bits_active_vint ? _GEN_827 : e_3_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1780 = io_op_bits_active_vint ? _GEN_828 : e_4_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1781 = io_op_bits_active_vint ? _GEN_829 : e_5_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1782 = io_op_bits_active_vint ? _GEN_830 : e_6_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1783 = io_op_bits_active_vint ? _GEN_831 : e_7_base_vs2_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1784 = io_op_bits_active_vint ? _GEN_832 : e_0_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1785 = io_op_bits_active_vint ? _GEN_833 : e_1_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1786 = io_op_bits_active_vint ? _GEN_834 : e_2_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1787 = io_op_bits_active_vint ? _GEN_835 : e_3_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1788 = io_op_bits_active_vint ? _GEN_836 : e_4_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1789 = io_op_bits_active_vint ? _GEN_837 : e_5_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1790 = io_op_bits_active_vint ? _GEN_838 : e_6_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1791 = io_op_bits_active_vint ? _GEN_839 : e_7_base_vs2_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1792 = io_op_bits_active_vint ? _GEN_840 : e_0_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1793 = io_op_bits_active_vint ? _GEN_841 : e_1_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1794 = io_op_bits_active_vint ? _GEN_842 : e_2_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1795 = io_op_bits_active_vint ? _GEN_843 : e_3_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1796 = io_op_bits_active_vint ? _GEN_844 : e_4_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1797 = io_op_bits_active_vint ? _GEN_845 : e_5_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1798 = io_op_bits_active_vint ? _GEN_846 : e_6_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1799 = io_op_bits_active_vint ? _GEN_847 : e_7_base_vs2_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1800 = io_op_bits_active_vint ? _GEN_848 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1801 = io_op_bits_active_vint ? _GEN_849 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1802 = io_op_bits_active_vint ? _GEN_850 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1803 = io_op_bits_active_vint ? _GEN_851 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1804 = io_op_bits_active_vint ? _GEN_852 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1805 = io_op_bits_active_vint ? _GEN_853 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1806 = io_op_bits_active_vint ? _GEN_854 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1807 = io_op_bits_active_vint ? _GEN_855 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [63:0] _GEN_1808 = io_op_bits_active_vint ? _GEN_856 : e_0_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1809 = io_op_bits_active_vint ? _GEN_857 : e_1_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1810 = io_op_bits_active_vint ? _GEN_858 : e_2_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1811 = io_op_bits_active_vint ? _GEN_859 : e_3_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1812 = io_op_bits_active_vint ? _GEN_860 : e_4_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1813 = io_op_bits_active_vint ? _GEN_861 : e_5_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1814 = io_op_bits_active_vint ? _GEN_862 : e_6_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [63:0] _GEN_1815 = io_op_bits_active_vint ? _GEN_863 : e_7_sreg_ss2; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1816 = io_op_bits_active_vint ? _GEN_1040 : e_0_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1817 = io_op_bits_active_vint ? _GEN_1041 : e_1_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1818 = io_op_bits_active_vint ? _GEN_1042 : e_2_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1819 = io_op_bits_active_vint ? _GEN_1043 : e_3_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1820 = io_op_bits_active_vint ? _GEN_1044 : e_4_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1821 = io_op_bits_active_vint ? _GEN_1045 : e_5_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1822 = io_op_bits_active_vint ? _GEN_1046 : e_6_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1823 = io_op_bits_active_vint ? _GEN_1047 : e_7_base_vd_id; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1824 = io_op_bits_active_vint ? _GEN_1056 : e_0_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1825 = io_op_bits_active_vint ? _GEN_1057 : e_1_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1826 = io_op_bits_active_vint ? _GEN_1058 : e_2_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1827 = io_op_bits_active_vint ? _GEN_1059 : e_3_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1828 = io_op_bits_active_vint ? _GEN_1060 : e_4_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1829 = io_op_bits_active_vint ? _GEN_1061 : e_5_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1830 = io_op_bits_active_vint ? _GEN_1062 : e_6_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1831 = io_op_bits_active_vint ? _GEN_1063 : e_7_base_vd_scalar; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1832 = io_op_bits_active_vint ? _GEN_1064 : e_0_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1833 = io_op_bits_active_vint ? _GEN_1065 : e_1_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1834 = io_op_bits_active_vint ? _GEN_1066 : e_2_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1835 = io_op_bits_active_vint ? _GEN_1067 : e_3_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1836 = io_op_bits_active_vint ? _GEN_1068 : e_4_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1837 = io_op_bits_active_vint ? _GEN_1069 : e_5_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1838 = io_op_bits_active_vint ? _GEN_1070 : e_6_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire  _GEN_1839 = io_op_bits_active_vint ? _GEN_1071 : e_7_base_vd_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1840 = io_op_bits_active_vint ? _GEN_1072 : e_0_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1841 = io_op_bits_active_vint ? _GEN_1073 : e_1_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1842 = io_op_bits_active_vint ? _GEN_1074 : e_2_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1843 = io_op_bits_active_vint ? _GEN_1075 : e_3_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1844 = io_op_bits_active_vint ? _GEN_1076 : e_4_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1845 = io_op_bits_active_vint ? _GEN_1077 : e_5_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1846 = io_op_bits_active_vint ? _GEN_1078 : e_6_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1847 = io_op_bits_active_vint ? _GEN_1079 : e_7_base_vd_prec; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_1848 = io_op_bits_active_vint ? _GEN_1080 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1849 = io_op_bits_active_vint ? _GEN_1081 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1850 = io_op_bits_active_vint ? _GEN_1082 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1851 = io_op_bits_active_vint ? _GEN_1083 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1852 = io_op_bits_active_vint ? _GEN_1084 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1853 = io_op_bits_active_vint ? _GEN_1085 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1854 = io_op_bits_active_vint ? _GEN_1086 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [7:0] _GEN_1855 = io_op_bits_active_vint ? _GEN_1087 : 8'h0; // @[sequencer-master.scala 640:39 sequencer-master.scala 411:33]
  wire [1:0] _GEN_1856 = io_op_bits_active_vint ? _GEN_1344 : e_0_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1857 = io_op_bits_active_vint ? _GEN_1345 : e_1_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1858 = io_op_bits_active_vint ? _GEN_1346 : e_2_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1859 = io_op_bits_active_vint ? _GEN_1347 : e_3_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1860 = io_op_bits_active_vint ? _GEN_1348 : e_4_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1861 = io_op_bits_active_vint ? _GEN_1349 : e_5_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1862 = io_op_bits_active_vint ? _GEN_1350 : e_6_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [1:0] _GEN_1863 = io_op_bits_active_vint ? _GEN_1351 : e_7_rports; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1864 = io_op_bits_active_vint ? _GEN_1376 : e_0_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1865 = io_op_bits_active_vint ? _GEN_1377 : e_1_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1866 = io_op_bits_active_vint ? _GEN_1378 : e_2_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1867 = io_op_bits_active_vint ? _GEN_1379 : e_3_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1868 = io_op_bits_active_vint ? _GEN_1380 : e_4_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1869 = io_op_bits_active_vint ? _GEN_1381 : e_5_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1870 = io_op_bits_active_vint ? _GEN_1382 : e_6_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [3:0] _GEN_1871 = io_op_bits_active_vint ? _GEN_1383 : e_7_wport_sram; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1872 = io_op_bits_active_vint ? _GEN_1392 : e_0_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1873 = io_op_bits_active_vint ? _GEN_1393 : e_1_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1874 = io_op_bits_active_vint ? _GEN_1394 : e_2_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1875 = io_op_bits_active_vint ? _GEN_1395 : e_3_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1876 = io_op_bits_active_vint ? _GEN_1396 : e_4_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1877 = io_op_bits_active_vint ? _GEN_1397 : e_5_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1878 = io_op_bits_active_vint ? _GEN_1398 : e_6_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1879 = io_op_bits_active_vint ? _GEN_1399 : e_7_wport_pred; // @[sequencer-master.scala 640:39 sequencer-master.scala 109:14]
  wire [2:0] _GEN_1881 = io_op_bits_active_vint ? _T_1645 : tail; // @[sequencer-master.scala 640:39 sequencer-master.scala 265:66 sequencer-master.scala 407:17]
  wire  _GEN_1882 = _GEN_32729 | _GEN_1400; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1883 = _GEN_32730 | _GEN_1401; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1884 = _GEN_32731 | _GEN_1402; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1885 = _GEN_32732 | _GEN_1403; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1886 = _GEN_32733 | _GEN_1404; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1887 = _GEN_32734 | _GEN_1405; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1888 = _GEN_32735 | _GEN_1406; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1889 = _GEN_32736 | _GEN_1407; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_1898 = 3'h0 == tail ? 1'h0 : _GEN_1416; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1899 = 3'h1 == tail ? 1'h0 : _GEN_1417; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1900 = 3'h2 == tail ? 1'h0 : _GEN_1418; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1901 = 3'h3 == tail ? 1'h0 : _GEN_1419; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1902 = 3'h4 == tail ? 1'h0 : _GEN_1420; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1903 = 3'h5 == tail ? 1'h0 : _GEN_1421; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1904 = 3'h6 == tail ? 1'h0 : _GEN_1422; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1905 = 3'h7 == tail ? 1'h0 : _GEN_1423; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_1906 = 3'h0 == tail ? 1'h0 : _GEN_1424; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1907 = 3'h1 == tail ? 1'h0 : _GEN_1425; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1908 = 3'h2 == tail ? 1'h0 : _GEN_1426; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1909 = 3'h3 == tail ? 1'h0 : _GEN_1427; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1910 = 3'h4 == tail ? 1'h0 : _GEN_1428; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1911 = 3'h5 == tail ? 1'h0 : _GEN_1429; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1912 = 3'h6 == tail ? 1'h0 : _GEN_1430; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1913 = 3'h7 == tail ? 1'h0 : _GEN_1431; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_1914 = 3'h0 == tail ? 1'h0 : _GEN_1432; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1915 = 3'h1 == tail ? 1'h0 : _GEN_1433; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1916 = 3'h2 == tail ? 1'h0 : _GEN_1434; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1917 = 3'h3 == tail ? 1'h0 : _GEN_1435; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1918 = 3'h4 == tail ? 1'h0 : _GEN_1436; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1919 = 3'h5 == tail ? 1'h0 : _GEN_1437; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1920 = 3'h6 == tail ? 1'h0 : _GEN_1438; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1921 = 3'h7 == tail ? 1'h0 : _GEN_1439; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_1922 = 3'h0 == tail ? 1'h0 : _GEN_1440; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1923 = 3'h1 == tail ? 1'h0 : _GEN_1441; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1924 = 3'h2 == tail ? 1'h0 : _GEN_1442; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1925 = 3'h3 == tail ? 1'h0 : _GEN_1443; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1926 = 3'h4 == tail ? 1'h0 : _GEN_1444; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1927 = 3'h5 == tail ? 1'h0 : _GEN_1445; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1928 = 3'h6 == tail ? 1'h0 : _GEN_1446; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1929 = 3'h7 == tail ? 1'h0 : _GEN_1447; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_1930 = 3'h0 == tail ? 1'h0 : _GEN_1448; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1931 = 3'h1 == tail ? 1'h0 : _GEN_1449; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1932 = 3'h2 == tail ? 1'h0 : _GEN_1450; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1933 = 3'h3 == tail ? 1'h0 : _GEN_1451; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1934 = 3'h4 == tail ? 1'h0 : _GEN_1452; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1935 = 3'h5 == tail ? 1'h0 : _GEN_1453; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1936 = 3'h6 == tail ? 1'h0 : _GEN_1454; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1937 = 3'h7 == tail ? 1'h0 : _GEN_1455; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_1938 = _GEN_32729 | _GEN_1456; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1939 = _GEN_32730 | _GEN_1457; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1940 = _GEN_32731 | _GEN_1458; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1941 = _GEN_32732 | _GEN_1459; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1942 = _GEN_32733 | _GEN_1460; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1943 = _GEN_32734 | _GEN_1461; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1944 = _GEN_32735 | _GEN_1462; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1945 = _GEN_32736 | _GEN_1463; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_1946 = 3'h0 == tail ? 1'h0 : _GEN_1464; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1947 = 3'h1 == tail ? 1'h0 : _GEN_1465; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1948 = 3'h2 == tail ? 1'h0 : _GEN_1466; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1949 = 3'h3 == tail ? 1'h0 : _GEN_1467; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1950 = 3'h4 == tail ? 1'h0 : _GEN_1468; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1951 = 3'h5 == tail ? 1'h0 : _GEN_1469; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1952 = 3'h6 == tail ? 1'h0 : _GEN_1470; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1953 = 3'h7 == tail ? 1'h0 : _GEN_1471; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1954 = 3'h0 == tail ? 1'h0 : _GEN_1472; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1955 = 3'h1 == tail ? 1'h0 : _GEN_1473; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1956 = 3'h2 == tail ? 1'h0 : _GEN_1474; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1957 = 3'h3 == tail ? 1'h0 : _GEN_1475; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1958 = 3'h4 == tail ? 1'h0 : _GEN_1476; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1959 = 3'h5 == tail ? 1'h0 : _GEN_1477; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1960 = 3'h6 == tail ? 1'h0 : _GEN_1478; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1961 = 3'h7 == tail ? 1'h0 : _GEN_1479; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1962 = 3'h0 == tail ? 1'h0 : _GEN_1480; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1963 = 3'h1 == tail ? 1'h0 : _GEN_1481; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1964 = 3'h2 == tail ? 1'h0 : _GEN_1482; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1965 = 3'h3 == tail ? 1'h0 : _GEN_1483; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1966 = 3'h4 == tail ? 1'h0 : _GEN_1484; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1967 = 3'h5 == tail ? 1'h0 : _GEN_1485; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1968 = 3'h6 == tail ? 1'h0 : _GEN_1486; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1969 = 3'h7 == tail ? 1'h0 : _GEN_1487; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1970 = 3'h0 == tail ? 1'h0 : _GEN_1488; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1971 = 3'h1 == tail ? 1'h0 : _GEN_1489; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1972 = 3'h2 == tail ? 1'h0 : _GEN_1490; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1973 = 3'h3 == tail ? 1'h0 : _GEN_1491; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1974 = 3'h4 == tail ? 1'h0 : _GEN_1492; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1975 = 3'h5 == tail ? 1'h0 : _GEN_1493; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1976 = 3'h6 == tail ? 1'h0 : _GEN_1494; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1977 = 3'h7 == tail ? 1'h0 : _GEN_1495; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1978 = 3'h0 == tail ? 1'h0 : _GEN_1496; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1979 = 3'h1 == tail ? 1'h0 : _GEN_1497; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1980 = 3'h2 == tail ? 1'h0 : _GEN_1498; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1981 = 3'h3 == tail ? 1'h0 : _GEN_1499; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1982 = 3'h4 == tail ? 1'h0 : _GEN_1500; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1983 = 3'h5 == tail ? 1'h0 : _GEN_1501; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1984 = 3'h6 == tail ? 1'h0 : _GEN_1502; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1985 = 3'h7 == tail ? 1'h0 : _GEN_1503; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_1986 = 3'h0 == tail ? 1'h0 : _GEN_1504; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1987 = 3'h1 == tail ? 1'h0 : _GEN_1505; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1988 = 3'h2 == tail ? 1'h0 : _GEN_1506; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1989 = 3'h3 == tail ? 1'h0 : _GEN_1507; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1990 = 3'h4 == tail ? 1'h0 : _GEN_1508; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1991 = 3'h5 == tail ? 1'h0 : _GEN_1509; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1992 = 3'h6 == tail ? 1'h0 : _GEN_1510; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1993 = 3'h7 == tail ? 1'h0 : _GEN_1511; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_1994 = 3'h0 == tail ? 1'h0 : _GEN_1512; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1995 = 3'h1 == tail ? 1'h0 : _GEN_1513; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1996 = 3'h2 == tail ? 1'h0 : _GEN_1514; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1997 = 3'h3 == tail ? 1'h0 : _GEN_1515; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1998 = 3'h4 == tail ? 1'h0 : _GEN_1516; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_1999 = 3'h5 == tail ? 1'h0 : _GEN_1517; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2000 = 3'h6 == tail ? 1'h0 : _GEN_1518; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2001 = 3'h7 == tail ? 1'h0 : _GEN_1519; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2002 = 3'h0 == tail ? 1'h0 : _GEN_1520; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2003 = 3'h1 == tail ? 1'h0 : _GEN_1521; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2004 = 3'h2 == tail ? 1'h0 : _GEN_1522; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2005 = 3'h3 == tail ? 1'h0 : _GEN_1523; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2006 = 3'h4 == tail ? 1'h0 : _GEN_1524; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2007 = 3'h5 == tail ? 1'h0 : _GEN_1525; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2008 = 3'h6 == tail ? 1'h0 : _GEN_1526; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2009 = 3'h7 == tail ? 1'h0 : _GEN_1527; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2010 = 3'h0 == tail ? 1'h0 : _GEN_1528; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2011 = 3'h1 == tail ? 1'h0 : _GEN_1529; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2012 = 3'h2 == tail ? 1'h0 : _GEN_1530; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2013 = 3'h3 == tail ? 1'h0 : _GEN_1531; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2014 = 3'h4 == tail ? 1'h0 : _GEN_1532; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2015 = 3'h5 == tail ? 1'h0 : _GEN_1533; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2016 = 3'h6 == tail ? 1'h0 : _GEN_1534; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2017 = 3'h7 == tail ? 1'h0 : _GEN_1535; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2018 = 3'h0 == tail ? 1'h0 : _GEN_1536; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2019 = 3'h1 == tail ? 1'h0 : _GEN_1537; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2020 = 3'h2 == tail ? 1'h0 : _GEN_1538; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2021 = 3'h3 == tail ? 1'h0 : _GEN_1539; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2022 = 3'h4 == tail ? 1'h0 : _GEN_1540; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2023 = 3'h5 == tail ? 1'h0 : _GEN_1541; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2024 = 3'h6 == tail ? 1'h0 : _GEN_1542; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2025 = 3'h7 == tail ? 1'h0 : _GEN_1543; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2026 = 3'h0 == tail ? 1'h0 : _GEN_1544; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2027 = 3'h1 == tail ? 1'h0 : _GEN_1545; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2028 = 3'h2 == tail ? 1'h0 : _GEN_1546; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2029 = 3'h3 == tail ? 1'h0 : _GEN_1547; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2030 = 3'h4 == tail ? 1'h0 : _GEN_1548; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2031 = 3'h5 == tail ? 1'h0 : _GEN_1549; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2032 = 3'h6 == tail ? 1'h0 : _GEN_1550; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2033 = 3'h7 == tail ? 1'h0 : _GEN_1551; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2034 = 3'h0 == tail ? 1'h0 : _GEN_1552; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2035 = 3'h1 == tail ? 1'h0 : _GEN_1553; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2036 = 3'h2 == tail ? 1'h0 : _GEN_1554; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2037 = 3'h3 == tail ? 1'h0 : _GEN_1555; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2038 = 3'h4 == tail ? 1'h0 : _GEN_1556; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2039 = 3'h5 == tail ? 1'h0 : _GEN_1557; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2040 = 3'h6 == tail ? 1'h0 : _GEN_1558; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2041 = 3'h7 == tail ? 1'h0 : _GEN_1559; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2042 = 3'h0 == tail ? 1'h0 : _GEN_1560; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2043 = 3'h1 == tail ? 1'h0 : _GEN_1561; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2044 = 3'h2 == tail ? 1'h0 : _GEN_1562; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2045 = 3'h3 == tail ? 1'h0 : _GEN_1563; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2046 = 3'h4 == tail ? 1'h0 : _GEN_1564; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2047 = 3'h5 == tail ? 1'h0 : _GEN_1565; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2048 = 3'h6 == tail ? 1'h0 : _GEN_1566; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2049 = 3'h7 == tail ? 1'h0 : _GEN_1567; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2050 = 3'h0 == tail ? 1'h0 : _GEN_1568; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2051 = 3'h1 == tail ? 1'h0 : _GEN_1569; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2052 = 3'h2 == tail ? 1'h0 : _GEN_1570; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2053 = 3'h3 == tail ? 1'h0 : _GEN_1571; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2054 = 3'h4 == tail ? 1'h0 : _GEN_1572; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2055 = 3'h5 == tail ? 1'h0 : _GEN_1573; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2056 = 3'h6 == tail ? 1'h0 : _GEN_1574; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2057 = 3'h7 == tail ? 1'h0 : _GEN_1575; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2058 = 3'h0 == tail ? 1'h0 : _GEN_1576; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2059 = 3'h1 == tail ? 1'h0 : _GEN_1577; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2060 = 3'h2 == tail ? 1'h0 : _GEN_1578; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2061 = 3'h3 == tail ? 1'h0 : _GEN_1579; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2062 = 3'h4 == tail ? 1'h0 : _GEN_1580; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2063 = 3'h5 == tail ? 1'h0 : _GEN_1581; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2064 = 3'h6 == tail ? 1'h0 : _GEN_1582; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2065 = 3'h7 == tail ? 1'h0 : _GEN_1583; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2066 = 3'h0 == tail ? 1'h0 : _GEN_1584; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2067 = 3'h1 == tail ? 1'h0 : _GEN_1585; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2068 = 3'h2 == tail ? 1'h0 : _GEN_1586; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2069 = 3'h3 == tail ? 1'h0 : _GEN_1587; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2070 = 3'h4 == tail ? 1'h0 : _GEN_1588; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2071 = 3'h5 == tail ? 1'h0 : _GEN_1589; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2072 = 3'h6 == tail ? 1'h0 : _GEN_1590; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2073 = 3'h7 == tail ? 1'h0 : _GEN_1591; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2074 = 3'h0 == tail ? 1'h0 : _GEN_1592; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2075 = 3'h1 == tail ? 1'h0 : _GEN_1593; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2076 = 3'h2 == tail ? 1'h0 : _GEN_1594; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2077 = 3'h3 == tail ? 1'h0 : _GEN_1595; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2078 = 3'h4 == tail ? 1'h0 : _GEN_1596; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2079 = 3'h5 == tail ? 1'h0 : _GEN_1597; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2080 = 3'h6 == tail ? 1'h0 : _GEN_1598; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2081 = 3'h7 == tail ? 1'h0 : _GEN_1599; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2082 = 3'h0 == tail ? 1'h0 : _GEN_1600; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2083 = 3'h1 == tail ? 1'h0 : _GEN_1601; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2084 = 3'h2 == tail ? 1'h0 : _GEN_1602; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2085 = 3'h3 == tail ? 1'h0 : _GEN_1603; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2086 = 3'h4 == tail ? 1'h0 : _GEN_1604; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2087 = 3'h5 == tail ? 1'h0 : _GEN_1605; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2088 = 3'h6 == tail ? 1'h0 : _GEN_1606; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2089 = 3'h7 == tail ? 1'h0 : _GEN_1607; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2090 = 3'h0 == tail ? 1'h0 : _GEN_1608; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2091 = 3'h1 == tail ? 1'h0 : _GEN_1609; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2092 = 3'h2 == tail ? 1'h0 : _GEN_1610; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2093 = 3'h3 == tail ? 1'h0 : _GEN_1611; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2094 = 3'h4 == tail ? 1'h0 : _GEN_1612; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2095 = 3'h5 == tail ? 1'h0 : _GEN_1613; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2096 = 3'h6 == tail ? 1'h0 : _GEN_1614; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2097 = 3'h7 == tail ? 1'h0 : _GEN_1615; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2098 = 3'h0 == tail ? 1'h0 : _GEN_1616; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2099 = 3'h1 == tail ? 1'h0 : _GEN_1617; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2100 = 3'h2 == tail ? 1'h0 : _GEN_1618; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2101 = 3'h3 == tail ? 1'h0 : _GEN_1619; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2102 = 3'h4 == tail ? 1'h0 : _GEN_1620; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2103 = 3'h5 == tail ? 1'h0 : _GEN_1621; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2104 = 3'h6 == tail ? 1'h0 : _GEN_1622; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2105 = 3'h7 == tail ? 1'h0 : _GEN_1623; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2106 = 3'h0 == tail ? 1'h0 : _GEN_1624; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2107 = 3'h1 == tail ? 1'h0 : _GEN_1625; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2108 = 3'h2 == tail ? 1'h0 : _GEN_1626; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2109 = 3'h3 == tail ? 1'h0 : _GEN_1627; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2110 = 3'h4 == tail ? 1'h0 : _GEN_1628; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2111 = 3'h5 == tail ? 1'h0 : _GEN_1629; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2112 = 3'h6 == tail ? 1'h0 : _GEN_1630; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2113 = 3'h7 == tail ? 1'h0 : _GEN_1631; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2114 = 3'h0 == tail ? 1'h0 : _GEN_1632; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2115 = 3'h1 == tail ? 1'h0 : _GEN_1633; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2116 = 3'h2 == tail ? 1'h0 : _GEN_1634; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2117 = 3'h3 == tail ? 1'h0 : _GEN_1635; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2118 = 3'h4 == tail ? 1'h0 : _GEN_1636; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2119 = 3'h5 == tail ? 1'h0 : _GEN_1637; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2120 = 3'h6 == tail ? 1'h0 : _GEN_1638; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2121 = 3'h7 == tail ? 1'h0 : _GEN_1639; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_2122 = 3'h0 == tail ? 1'h0 : _GEN_1640; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2123 = 3'h1 == tail ? 1'h0 : _GEN_1641; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2124 = 3'h2 == tail ? 1'h0 : _GEN_1642; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2125 = 3'h3 == tail ? 1'h0 : _GEN_1643; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2126 = 3'h4 == tail ? 1'h0 : _GEN_1644; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2127 = 3'h5 == tail ? 1'h0 : _GEN_1645; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2128 = 3'h6 == tail ? 1'h0 : _GEN_1646; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2129 = 3'h7 == tail ? 1'h0 : _GEN_1647; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_2130 = 3'h0 == tail ? 1'h0 : _GEN_1648; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2131 = 3'h1 == tail ? 1'h0 : _GEN_1649; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2132 = 3'h2 == tail ? 1'h0 : _GEN_1650; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2133 = 3'h3 == tail ? 1'h0 : _GEN_1651; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2134 = 3'h4 == tail ? 1'h0 : _GEN_1652; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2135 = 3'h5 == tail ? 1'h0 : _GEN_1653; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2136 = 3'h6 == tail ? 1'h0 : _GEN_1654; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2137 = 3'h7 == tail ? 1'h0 : _GEN_1655; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_2138 = 3'h0 == tail ? 1'h0 : _GEN_1656; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2139 = 3'h1 == tail ? 1'h0 : _GEN_1657; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2140 = 3'h2 == tail ? 1'h0 : _GEN_1658; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2141 = 3'h3 == tail ? 1'h0 : _GEN_1659; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2142 = 3'h4 == tail ? 1'h0 : _GEN_1660; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2143 = 3'h5 == tail ? 1'h0 : _GEN_1661; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2144 = 3'h6 == tail ? 1'h0 : _GEN_1662; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2145 = 3'h7 == tail ? 1'h0 : _GEN_1663; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_2154 = _GEN_32729 | e_0_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2155 = _GEN_32730 | e_1_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2156 = _GEN_32731 | e_2_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2157 = _GEN_32732 | e_3_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2158 = _GEN_32733 | e_4_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2159 = _GEN_32734 | e_5_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2160 = _GEN_32735 | e_6_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_2161 = _GEN_32736 | e_7_active_vipu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_2162 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_1680; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2163 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_1681; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2164 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_1682; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2165 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_1683; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2166 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_1684; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2167 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_1685; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2168 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_1686; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_2169 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_1687; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [7:0] _GEN_2170 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_1720; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2171 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_1721; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2172 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_1722; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2173 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_1723; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2174 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_1724; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2175 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_1725; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2176 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_1726; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2177 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_1727; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2178 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_1906; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2179 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_1907; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2180 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_1908; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2181 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_1909; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2182 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_1910; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2183 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_1911; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2184 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_1912; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2185 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_1913; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2186 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_1728; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2187 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_1729; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2188 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_1730; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2189 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_1731; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2190 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_1732; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2191 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_1733; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2192 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_1734; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2193 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_1735; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2194 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_1736; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2195 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_1737; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2196 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_1738; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2197 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_1739; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2198 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_1740; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2199 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_1741; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2200 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_1742; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2201 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_1743; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2202 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_1744; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2203 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_1745; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2204 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_1746; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2205 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_1747; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2206 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_1748; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2207 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_1749; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2208 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_1750; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2209 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_1751; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2210 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_1752; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2211 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_1753; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2212 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_1754; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2213 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_1755; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2214 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_1756; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2215 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_1757; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2216 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_1758; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2217 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_1759; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_2218 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_1760; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2219 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_1761; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2220 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_1762; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2221 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_1763; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2222 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_1764; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2223 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_1765; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2224 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_1766; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2225 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_1767; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2226 = _T_189 ? _GEN_2218 : _GEN_1760; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2227 = _T_189 ? _GEN_2219 : _GEN_1761; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2228 = _T_189 ? _GEN_2220 : _GEN_1762; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2229 = _T_189 ? _GEN_2221 : _GEN_1763; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2230 = _T_189 ? _GEN_2222 : _GEN_1764; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2231 = _T_189 ? _GEN_2223 : _GEN_1765; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2232 = _T_189 ? _GEN_2224 : _GEN_1766; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2233 = _T_189 ? _GEN_2225 : _GEN_1767; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_2234 = io_op_bits_base_vs1_valid ? _GEN_2170 : _GEN_1720; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2235 = io_op_bits_base_vs1_valid ? _GEN_2171 : _GEN_1721; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2236 = io_op_bits_base_vs1_valid ? _GEN_2172 : _GEN_1722; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2237 = io_op_bits_base_vs1_valid ? _GEN_2173 : _GEN_1723; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2238 = io_op_bits_base_vs1_valid ? _GEN_2174 : _GEN_1724; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2239 = io_op_bits_base_vs1_valid ? _GEN_2175 : _GEN_1725; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2240 = io_op_bits_base_vs1_valid ? _GEN_2176 : _GEN_1726; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2241 = io_op_bits_base_vs1_valid ? _GEN_2177 : _GEN_1727; // @[sequencer-master.scala 328:47]
  wire  _GEN_2242 = io_op_bits_base_vs1_valid ? _GEN_2178 : _GEN_1906; // @[sequencer-master.scala 328:47]
  wire  _GEN_2243 = io_op_bits_base_vs1_valid ? _GEN_2179 : _GEN_1907; // @[sequencer-master.scala 328:47]
  wire  _GEN_2244 = io_op_bits_base_vs1_valid ? _GEN_2180 : _GEN_1908; // @[sequencer-master.scala 328:47]
  wire  _GEN_2245 = io_op_bits_base_vs1_valid ? _GEN_2181 : _GEN_1909; // @[sequencer-master.scala 328:47]
  wire  _GEN_2246 = io_op_bits_base_vs1_valid ? _GEN_2182 : _GEN_1910; // @[sequencer-master.scala 328:47]
  wire  _GEN_2247 = io_op_bits_base_vs1_valid ? _GEN_2183 : _GEN_1911; // @[sequencer-master.scala 328:47]
  wire  _GEN_2248 = io_op_bits_base_vs1_valid ? _GEN_2184 : _GEN_1912; // @[sequencer-master.scala 328:47]
  wire  _GEN_2249 = io_op_bits_base_vs1_valid ? _GEN_2185 : _GEN_1913; // @[sequencer-master.scala 328:47]
  wire  _GEN_2250 = io_op_bits_base_vs1_valid ? _GEN_2186 : _GEN_1728; // @[sequencer-master.scala 328:47]
  wire  _GEN_2251 = io_op_bits_base_vs1_valid ? _GEN_2187 : _GEN_1729; // @[sequencer-master.scala 328:47]
  wire  _GEN_2252 = io_op_bits_base_vs1_valid ? _GEN_2188 : _GEN_1730; // @[sequencer-master.scala 328:47]
  wire  _GEN_2253 = io_op_bits_base_vs1_valid ? _GEN_2189 : _GEN_1731; // @[sequencer-master.scala 328:47]
  wire  _GEN_2254 = io_op_bits_base_vs1_valid ? _GEN_2190 : _GEN_1732; // @[sequencer-master.scala 328:47]
  wire  _GEN_2255 = io_op_bits_base_vs1_valid ? _GEN_2191 : _GEN_1733; // @[sequencer-master.scala 328:47]
  wire  _GEN_2256 = io_op_bits_base_vs1_valid ? _GEN_2192 : _GEN_1734; // @[sequencer-master.scala 328:47]
  wire  _GEN_2257 = io_op_bits_base_vs1_valid ? _GEN_2193 : _GEN_1735; // @[sequencer-master.scala 328:47]
  wire  _GEN_2258 = io_op_bits_base_vs1_valid ? _GEN_2194 : _GEN_1736; // @[sequencer-master.scala 328:47]
  wire  _GEN_2259 = io_op_bits_base_vs1_valid ? _GEN_2195 : _GEN_1737; // @[sequencer-master.scala 328:47]
  wire  _GEN_2260 = io_op_bits_base_vs1_valid ? _GEN_2196 : _GEN_1738; // @[sequencer-master.scala 328:47]
  wire  _GEN_2261 = io_op_bits_base_vs1_valid ? _GEN_2197 : _GEN_1739; // @[sequencer-master.scala 328:47]
  wire  _GEN_2262 = io_op_bits_base_vs1_valid ? _GEN_2198 : _GEN_1740; // @[sequencer-master.scala 328:47]
  wire  _GEN_2263 = io_op_bits_base_vs1_valid ? _GEN_2199 : _GEN_1741; // @[sequencer-master.scala 328:47]
  wire  _GEN_2264 = io_op_bits_base_vs1_valid ? _GEN_2200 : _GEN_1742; // @[sequencer-master.scala 328:47]
  wire  _GEN_2265 = io_op_bits_base_vs1_valid ? _GEN_2201 : _GEN_1743; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2266 = io_op_bits_base_vs1_valid ? _GEN_2202 : _GEN_1744; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2267 = io_op_bits_base_vs1_valid ? _GEN_2203 : _GEN_1745; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2268 = io_op_bits_base_vs1_valid ? _GEN_2204 : _GEN_1746; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2269 = io_op_bits_base_vs1_valid ? _GEN_2205 : _GEN_1747; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2270 = io_op_bits_base_vs1_valid ? _GEN_2206 : _GEN_1748; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2271 = io_op_bits_base_vs1_valid ? _GEN_2207 : _GEN_1749; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2272 = io_op_bits_base_vs1_valid ? _GEN_2208 : _GEN_1750; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2273 = io_op_bits_base_vs1_valid ? _GEN_2209 : _GEN_1751; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2274 = io_op_bits_base_vs1_valid ? _GEN_2210 : _GEN_1752; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2275 = io_op_bits_base_vs1_valid ? _GEN_2211 : _GEN_1753; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2276 = io_op_bits_base_vs1_valid ? _GEN_2212 : _GEN_1754; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2277 = io_op_bits_base_vs1_valid ? _GEN_2213 : _GEN_1755; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2278 = io_op_bits_base_vs1_valid ? _GEN_2214 : _GEN_1756; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2279 = io_op_bits_base_vs1_valid ? _GEN_2215 : _GEN_1757; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2280 = io_op_bits_base_vs1_valid ? _GEN_2216 : _GEN_1758; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2281 = io_op_bits_base_vs1_valid ? _GEN_2217 : _GEN_1759; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2282 = io_op_bits_base_vs1_valid ? _GEN_2226 : _GEN_1760; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2283 = io_op_bits_base_vs1_valid ? _GEN_2227 : _GEN_1761; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2284 = io_op_bits_base_vs1_valid ? _GEN_2228 : _GEN_1762; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2285 = io_op_bits_base_vs1_valid ? _GEN_2229 : _GEN_1763; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2286 = io_op_bits_base_vs1_valid ? _GEN_2230 : _GEN_1764; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2287 = io_op_bits_base_vs1_valid ? _GEN_2231 : _GEN_1765; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2288 = io_op_bits_base_vs1_valid ? _GEN_2232 : _GEN_1766; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2289 = io_op_bits_base_vs1_valid ? _GEN_2233 : _GEN_1767; // @[sequencer-master.scala 328:47]
  wire  _GEN_2290 = _GEN_32729 | _GEN_1946; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2291 = _GEN_32730 | _GEN_1947; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2292 = _GEN_32731 | _GEN_1948; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2293 = _GEN_32732 | _GEN_1949; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2294 = _GEN_32733 | _GEN_1950; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2295 = _GEN_32734 | _GEN_1951; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2296 = _GEN_32735 | _GEN_1952; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2297 = _GEN_32736 | _GEN_1953; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2298 = _T_203 ? _GEN_2290 : _GEN_1946; // @[sequencer-master.scala 154:24]
  wire  _GEN_2299 = _T_203 ? _GEN_2291 : _GEN_1947; // @[sequencer-master.scala 154:24]
  wire  _GEN_2300 = _T_203 ? _GEN_2292 : _GEN_1948; // @[sequencer-master.scala 154:24]
  wire  _GEN_2301 = _T_203 ? _GEN_2293 : _GEN_1949; // @[sequencer-master.scala 154:24]
  wire  _GEN_2302 = _T_203 ? _GEN_2294 : _GEN_1950; // @[sequencer-master.scala 154:24]
  wire  _GEN_2303 = _T_203 ? _GEN_2295 : _GEN_1951; // @[sequencer-master.scala 154:24]
  wire  _GEN_2304 = _T_203 ? _GEN_2296 : _GEN_1952; // @[sequencer-master.scala 154:24]
  wire  _GEN_2305 = _T_203 ? _GEN_2297 : _GEN_1953; // @[sequencer-master.scala 154:24]
  wire  _GEN_2306 = _GEN_32729 | _GEN_1970; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2307 = _GEN_32730 | _GEN_1971; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2308 = _GEN_32731 | _GEN_1972; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2309 = _GEN_32732 | _GEN_1973; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2310 = _GEN_32733 | _GEN_1974; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2311 = _GEN_32734 | _GEN_1975; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2312 = _GEN_32735 | _GEN_1976; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2313 = _GEN_32736 | _GEN_1977; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2314 = _T_225 ? _GEN_2306 : _GEN_1970; // @[sequencer-master.scala 154:24]
  wire  _GEN_2315 = _T_225 ? _GEN_2307 : _GEN_1971; // @[sequencer-master.scala 154:24]
  wire  _GEN_2316 = _T_225 ? _GEN_2308 : _GEN_1972; // @[sequencer-master.scala 154:24]
  wire  _GEN_2317 = _T_225 ? _GEN_2309 : _GEN_1973; // @[sequencer-master.scala 154:24]
  wire  _GEN_2318 = _T_225 ? _GEN_2310 : _GEN_1974; // @[sequencer-master.scala 154:24]
  wire  _GEN_2319 = _T_225 ? _GEN_2311 : _GEN_1975; // @[sequencer-master.scala 154:24]
  wire  _GEN_2320 = _T_225 ? _GEN_2312 : _GEN_1976; // @[sequencer-master.scala 154:24]
  wire  _GEN_2321 = _T_225 ? _GEN_2313 : _GEN_1977; // @[sequencer-master.scala 154:24]
  wire  _GEN_2322 = _GEN_32729 | _GEN_1994; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2323 = _GEN_32730 | _GEN_1995; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2324 = _GEN_32731 | _GEN_1996; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2325 = _GEN_32732 | _GEN_1997; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2326 = _GEN_32733 | _GEN_1998; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2327 = _GEN_32734 | _GEN_1999; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2328 = _GEN_32735 | _GEN_2000; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2329 = _GEN_32736 | _GEN_2001; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2330 = _T_247 ? _GEN_2322 : _GEN_1994; // @[sequencer-master.scala 154:24]
  wire  _GEN_2331 = _T_247 ? _GEN_2323 : _GEN_1995; // @[sequencer-master.scala 154:24]
  wire  _GEN_2332 = _T_247 ? _GEN_2324 : _GEN_1996; // @[sequencer-master.scala 154:24]
  wire  _GEN_2333 = _T_247 ? _GEN_2325 : _GEN_1997; // @[sequencer-master.scala 154:24]
  wire  _GEN_2334 = _T_247 ? _GEN_2326 : _GEN_1998; // @[sequencer-master.scala 154:24]
  wire  _GEN_2335 = _T_247 ? _GEN_2327 : _GEN_1999; // @[sequencer-master.scala 154:24]
  wire  _GEN_2336 = _T_247 ? _GEN_2328 : _GEN_2000; // @[sequencer-master.scala 154:24]
  wire  _GEN_2337 = _T_247 ? _GEN_2329 : _GEN_2001; // @[sequencer-master.scala 154:24]
  wire  _GEN_2338 = _GEN_32729 | _GEN_2018; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2339 = _GEN_32730 | _GEN_2019; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2340 = _GEN_32731 | _GEN_2020; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2341 = _GEN_32732 | _GEN_2021; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2342 = _GEN_32733 | _GEN_2022; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2343 = _GEN_32734 | _GEN_2023; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2344 = _GEN_32735 | _GEN_2024; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2345 = _GEN_32736 | _GEN_2025; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2346 = _T_269 ? _GEN_2338 : _GEN_2018; // @[sequencer-master.scala 154:24]
  wire  _GEN_2347 = _T_269 ? _GEN_2339 : _GEN_2019; // @[sequencer-master.scala 154:24]
  wire  _GEN_2348 = _T_269 ? _GEN_2340 : _GEN_2020; // @[sequencer-master.scala 154:24]
  wire  _GEN_2349 = _T_269 ? _GEN_2341 : _GEN_2021; // @[sequencer-master.scala 154:24]
  wire  _GEN_2350 = _T_269 ? _GEN_2342 : _GEN_2022; // @[sequencer-master.scala 154:24]
  wire  _GEN_2351 = _T_269 ? _GEN_2343 : _GEN_2023; // @[sequencer-master.scala 154:24]
  wire  _GEN_2352 = _T_269 ? _GEN_2344 : _GEN_2024; // @[sequencer-master.scala 154:24]
  wire  _GEN_2353 = _T_269 ? _GEN_2345 : _GEN_2025; // @[sequencer-master.scala 154:24]
  wire  _GEN_2354 = _GEN_32729 | _GEN_2042; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2355 = _GEN_32730 | _GEN_2043; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2356 = _GEN_32731 | _GEN_2044; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2357 = _GEN_32732 | _GEN_2045; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2358 = _GEN_32733 | _GEN_2046; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2359 = _GEN_32734 | _GEN_2047; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2360 = _GEN_32735 | _GEN_2048; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2361 = _GEN_32736 | _GEN_2049; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2362 = _T_291 ? _GEN_2354 : _GEN_2042; // @[sequencer-master.scala 154:24]
  wire  _GEN_2363 = _T_291 ? _GEN_2355 : _GEN_2043; // @[sequencer-master.scala 154:24]
  wire  _GEN_2364 = _T_291 ? _GEN_2356 : _GEN_2044; // @[sequencer-master.scala 154:24]
  wire  _GEN_2365 = _T_291 ? _GEN_2357 : _GEN_2045; // @[sequencer-master.scala 154:24]
  wire  _GEN_2366 = _T_291 ? _GEN_2358 : _GEN_2046; // @[sequencer-master.scala 154:24]
  wire  _GEN_2367 = _T_291 ? _GEN_2359 : _GEN_2047; // @[sequencer-master.scala 154:24]
  wire  _GEN_2368 = _T_291 ? _GEN_2360 : _GEN_2048; // @[sequencer-master.scala 154:24]
  wire  _GEN_2369 = _T_291 ? _GEN_2361 : _GEN_2049; // @[sequencer-master.scala 154:24]
  wire  _GEN_2370 = _GEN_32729 | _GEN_2066; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2371 = _GEN_32730 | _GEN_2067; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2372 = _GEN_32731 | _GEN_2068; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2373 = _GEN_32732 | _GEN_2069; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2374 = _GEN_32733 | _GEN_2070; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2375 = _GEN_32734 | _GEN_2071; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2376 = _GEN_32735 | _GEN_2072; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2377 = _GEN_32736 | _GEN_2073; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2378 = _T_313 ? _GEN_2370 : _GEN_2066; // @[sequencer-master.scala 154:24]
  wire  _GEN_2379 = _T_313 ? _GEN_2371 : _GEN_2067; // @[sequencer-master.scala 154:24]
  wire  _GEN_2380 = _T_313 ? _GEN_2372 : _GEN_2068; // @[sequencer-master.scala 154:24]
  wire  _GEN_2381 = _T_313 ? _GEN_2373 : _GEN_2069; // @[sequencer-master.scala 154:24]
  wire  _GEN_2382 = _T_313 ? _GEN_2374 : _GEN_2070; // @[sequencer-master.scala 154:24]
  wire  _GEN_2383 = _T_313 ? _GEN_2375 : _GEN_2071; // @[sequencer-master.scala 154:24]
  wire  _GEN_2384 = _T_313 ? _GEN_2376 : _GEN_2072; // @[sequencer-master.scala 154:24]
  wire  _GEN_2385 = _T_313 ? _GEN_2377 : _GEN_2073; // @[sequencer-master.scala 154:24]
  wire  _GEN_2386 = _GEN_32729 | _GEN_2090; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2387 = _GEN_32730 | _GEN_2091; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2388 = _GEN_32731 | _GEN_2092; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2389 = _GEN_32732 | _GEN_2093; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2390 = _GEN_32733 | _GEN_2094; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2391 = _GEN_32734 | _GEN_2095; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2392 = _GEN_32735 | _GEN_2096; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2393 = _GEN_32736 | _GEN_2097; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2394 = _T_335 ? _GEN_2386 : _GEN_2090; // @[sequencer-master.scala 154:24]
  wire  _GEN_2395 = _T_335 ? _GEN_2387 : _GEN_2091; // @[sequencer-master.scala 154:24]
  wire  _GEN_2396 = _T_335 ? _GEN_2388 : _GEN_2092; // @[sequencer-master.scala 154:24]
  wire  _GEN_2397 = _T_335 ? _GEN_2389 : _GEN_2093; // @[sequencer-master.scala 154:24]
  wire  _GEN_2398 = _T_335 ? _GEN_2390 : _GEN_2094; // @[sequencer-master.scala 154:24]
  wire  _GEN_2399 = _T_335 ? _GEN_2391 : _GEN_2095; // @[sequencer-master.scala 154:24]
  wire  _GEN_2400 = _T_335 ? _GEN_2392 : _GEN_2096; // @[sequencer-master.scala 154:24]
  wire  _GEN_2401 = _T_335 ? _GEN_2393 : _GEN_2097; // @[sequencer-master.scala 154:24]
  wire  _GEN_2402 = _GEN_32729 | _GEN_2114; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2403 = _GEN_32730 | _GEN_2115; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2404 = _GEN_32731 | _GEN_2116; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2405 = _GEN_32732 | _GEN_2117; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2406 = _GEN_32733 | _GEN_2118; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2407 = _GEN_32734 | _GEN_2119; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2408 = _GEN_32735 | _GEN_2120; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2409 = _GEN_32736 | _GEN_2121; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2410 = _T_357 ? _GEN_2402 : _GEN_2114; // @[sequencer-master.scala 154:24]
  wire  _GEN_2411 = _T_357 ? _GEN_2403 : _GEN_2115; // @[sequencer-master.scala 154:24]
  wire  _GEN_2412 = _T_357 ? _GEN_2404 : _GEN_2116; // @[sequencer-master.scala 154:24]
  wire  _GEN_2413 = _T_357 ? _GEN_2405 : _GEN_2117; // @[sequencer-master.scala 154:24]
  wire  _GEN_2414 = _T_357 ? _GEN_2406 : _GEN_2118; // @[sequencer-master.scala 154:24]
  wire  _GEN_2415 = _T_357 ? _GEN_2407 : _GEN_2119; // @[sequencer-master.scala 154:24]
  wire  _GEN_2416 = _T_357 ? _GEN_2408 : _GEN_2120; // @[sequencer-master.scala 154:24]
  wire  _GEN_2417 = _T_357 ? _GEN_2409 : _GEN_2121; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_2418 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_1768; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2419 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_1769; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2420 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_1770; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2421 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_1771; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2422 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_1772; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2423 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_1773; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2424 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_1774; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2425 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_1775; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2426 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_1914; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2427 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_1915; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2428 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_1916; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2429 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_1917; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2430 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_1918; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2431 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_1919; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2432 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_1920; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2433 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_1921; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2434 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_1776; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2435 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_1777; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2436 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_1778; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2437 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_1779; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2438 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_1780; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2439 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_1781; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2440 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_1782; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2441 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_1783; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2442 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_1784; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2443 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_1785; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2444 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_1786; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2445 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_1787; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2446 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_1788; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2447 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_1789; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2448 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_1790; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2449 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_1791; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2450 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_1792; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2451 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_1793; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2452 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_1794; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2453 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_1795; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2454 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_1796; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2455 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_1797; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2456 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_1798; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_2457 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_1799; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_2458 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_1800; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2459 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_1801; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2460 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_1802; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2461 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_1803; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2462 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_1804; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2463 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_1805; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2464 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_1806; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_2465 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_1807; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_2466 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_1808; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2467 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_1809; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2468 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_1810; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2469 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_1811; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2470 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_1812; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2471 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_1813; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2472 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_1814; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2473 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_1815; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_2474 = _T_366 ? _GEN_2466 : _GEN_1808; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2475 = _T_366 ? _GEN_2467 : _GEN_1809; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2476 = _T_366 ? _GEN_2468 : _GEN_1810; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2477 = _T_366 ? _GEN_2469 : _GEN_1811; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2478 = _T_366 ? _GEN_2470 : _GEN_1812; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2479 = _T_366 ? _GEN_2471 : _GEN_1813; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2480 = _T_366 ? _GEN_2472 : _GEN_1814; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_2481 = _T_366 ? _GEN_2473 : _GEN_1815; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_2482 = io_op_bits_base_vs2_valid ? _GEN_2418 : _GEN_1768; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2483 = io_op_bits_base_vs2_valid ? _GEN_2419 : _GEN_1769; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2484 = io_op_bits_base_vs2_valid ? _GEN_2420 : _GEN_1770; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2485 = io_op_bits_base_vs2_valid ? _GEN_2421 : _GEN_1771; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2486 = io_op_bits_base_vs2_valid ? _GEN_2422 : _GEN_1772; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2487 = io_op_bits_base_vs2_valid ? _GEN_2423 : _GEN_1773; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2488 = io_op_bits_base_vs2_valid ? _GEN_2424 : _GEN_1774; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2489 = io_op_bits_base_vs2_valid ? _GEN_2425 : _GEN_1775; // @[sequencer-master.scala 328:47]
  wire  _GEN_2490 = io_op_bits_base_vs2_valid ? _GEN_2426 : _GEN_1914; // @[sequencer-master.scala 328:47]
  wire  _GEN_2491 = io_op_bits_base_vs2_valid ? _GEN_2427 : _GEN_1915; // @[sequencer-master.scala 328:47]
  wire  _GEN_2492 = io_op_bits_base_vs2_valid ? _GEN_2428 : _GEN_1916; // @[sequencer-master.scala 328:47]
  wire  _GEN_2493 = io_op_bits_base_vs2_valid ? _GEN_2429 : _GEN_1917; // @[sequencer-master.scala 328:47]
  wire  _GEN_2494 = io_op_bits_base_vs2_valid ? _GEN_2430 : _GEN_1918; // @[sequencer-master.scala 328:47]
  wire  _GEN_2495 = io_op_bits_base_vs2_valid ? _GEN_2431 : _GEN_1919; // @[sequencer-master.scala 328:47]
  wire  _GEN_2496 = io_op_bits_base_vs2_valid ? _GEN_2432 : _GEN_1920; // @[sequencer-master.scala 328:47]
  wire  _GEN_2497 = io_op_bits_base_vs2_valid ? _GEN_2433 : _GEN_1921; // @[sequencer-master.scala 328:47]
  wire  _GEN_2498 = io_op_bits_base_vs2_valid ? _GEN_2434 : _GEN_1776; // @[sequencer-master.scala 328:47]
  wire  _GEN_2499 = io_op_bits_base_vs2_valid ? _GEN_2435 : _GEN_1777; // @[sequencer-master.scala 328:47]
  wire  _GEN_2500 = io_op_bits_base_vs2_valid ? _GEN_2436 : _GEN_1778; // @[sequencer-master.scala 328:47]
  wire  _GEN_2501 = io_op_bits_base_vs2_valid ? _GEN_2437 : _GEN_1779; // @[sequencer-master.scala 328:47]
  wire  _GEN_2502 = io_op_bits_base_vs2_valid ? _GEN_2438 : _GEN_1780; // @[sequencer-master.scala 328:47]
  wire  _GEN_2503 = io_op_bits_base_vs2_valid ? _GEN_2439 : _GEN_1781; // @[sequencer-master.scala 328:47]
  wire  _GEN_2504 = io_op_bits_base_vs2_valid ? _GEN_2440 : _GEN_1782; // @[sequencer-master.scala 328:47]
  wire  _GEN_2505 = io_op_bits_base_vs2_valid ? _GEN_2441 : _GEN_1783; // @[sequencer-master.scala 328:47]
  wire  _GEN_2506 = io_op_bits_base_vs2_valid ? _GEN_2442 : _GEN_1784; // @[sequencer-master.scala 328:47]
  wire  _GEN_2507 = io_op_bits_base_vs2_valid ? _GEN_2443 : _GEN_1785; // @[sequencer-master.scala 328:47]
  wire  _GEN_2508 = io_op_bits_base_vs2_valid ? _GEN_2444 : _GEN_1786; // @[sequencer-master.scala 328:47]
  wire  _GEN_2509 = io_op_bits_base_vs2_valid ? _GEN_2445 : _GEN_1787; // @[sequencer-master.scala 328:47]
  wire  _GEN_2510 = io_op_bits_base_vs2_valid ? _GEN_2446 : _GEN_1788; // @[sequencer-master.scala 328:47]
  wire  _GEN_2511 = io_op_bits_base_vs2_valid ? _GEN_2447 : _GEN_1789; // @[sequencer-master.scala 328:47]
  wire  _GEN_2512 = io_op_bits_base_vs2_valid ? _GEN_2448 : _GEN_1790; // @[sequencer-master.scala 328:47]
  wire  _GEN_2513 = io_op_bits_base_vs2_valid ? _GEN_2449 : _GEN_1791; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2514 = io_op_bits_base_vs2_valid ? _GEN_2450 : _GEN_1792; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2515 = io_op_bits_base_vs2_valid ? _GEN_2451 : _GEN_1793; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2516 = io_op_bits_base_vs2_valid ? _GEN_2452 : _GEN_1794; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2517 = io_op_bits_base_vs2_valid ? _GEN_2453 : _GEN_1795; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2518 = io_op_bits_base_vs2_valid ? _GEN_2454 : _GEN_1796; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2519 = io_op_bits_base_vs2_valid ? _GEN_2455 : _GEN_1797; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2520 = io_op_bits_base_vs2_valid ? _GEN_2456 : _GEN_1798; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_2521 = io_op_bits_base_vs2_valid ? _GEN_2457 : _GEN_1799; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2522 = io_op_bits_base_vs2_valid ? _GEN_2458 : _GEN_1800; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2523 = io_op_bits_base_vs2_valid ? _GEN_2459 : _GEN_1801; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2524 = io_op_bits_base_vs2_valid ? _GEN_2460 : _GEN_1802; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2525 = io_op_bits_base_vs2_valid ? _GEN_2461 : _GEN_1803; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2526 = io_op_bits_base_vs2_valid ? _GEN_2462 : _GEN_1804; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2527 = io_op_bits_base_vs2_valid ? _GEN_2463 : _GEN_1805; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2528 = io_op_bits_base_vs2_valid ? _GEN_2464 : _GEN_1806; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_2529 = io_op_bits_base_vs2_valid ? _GEN_2465 : _GEN_1807; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2530 = io_op_bits_base_vs2_valid ? _GEN_2474 : _GEN_1808; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2531 = io_op_bits_base_vs2_valid ? _GEN_2475 : _GEN_1809; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2532 = io_op_bits_base_vs2_valid ? _GEN_2476 : _GEN_1810; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2533 = io_op_bits_base_vs2_valid ? _GEN_2477 : _GEN_1811; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2534 = io_op_bits_base_vs2_valid ? _GEN_2478 : _GEN_1812; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2535 = io_op_bits_base_vs2_valid ? _GEN_2479 : _GEN_1813; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2536 = io_op_bits_base_vs2_valid ? _GEN_2480 : _GEN_1814; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_2537 = io_op_bits_base_vs2_valid ? _GEN_2481 : _GEN_1815; // @[sequencer-master.scala 328:47]
  wire  _GEN_2538 = _GEN_32729 | _GEN_2298; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2539 = _GEN_32730 | _GEN_2299; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2540 = _GEN_32731 | _GEN_2300; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2541 = _GEN_32732 | _GEN_2301; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2542 = _GEN_32733 | _GEN_2302; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2543 = _GEN_32734 | _GEN_2303; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2544 = _GEN_32735 | _GEN_2304; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2545 = _GEN_32736 | _GEN_2305; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2546 = _T_380 ? _GEN_2538 : _GEN_2298; // @[sequencer-master.scala 154:24]
  wire  _GEN_2547 = _T_380 ? _GEN_2539 : _GEN_2299; // @[sequencer-master.scala 154:24]
  wire  _GEN_2548 = _T_380 ? _GEN_2540 : _GEN_2300; // @[sequencer-master.scala 154:24]
  wire  _GEN_2549 = _T_380 ? _GEN_2541 : _GEN_2301; // @[sequencer-master.scala 154:24]
  wire  _GEN_2550 = _T_380 ? _GEN_2542 : _GEN_2302; // @[sequencer-master.scala 154:24]
  wire  _GEN_2551 = _T_380 ? _GEN_2543 : _GEN_2303; // @[sequencer-master.scala 154:24]
  wire  _GEN_2552 = _T_380 ? _GEN_2544 : _GEN_2304; // @[sequencer-master.scala 154:24]
  wire  _GEN_2553 = _T_380 ? _GEN_2545 : _GEN_2305; // @[sequencer-master.scala 154:24]
  wire  _GEN_2554 = _GEN_32729 | _GEN_2314; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2555 = _GEN_32730 | _GEN_2315; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2556 = _GEN_32731 | _GEN_2316; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2557 = _GEN_32732 | _GEN_2317; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2558 = _GEN_32733 | _GEN_2318; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2559 = _GEN_32734 | _GEN_2319; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2560 = _GEN_32735 | _GEN_2320; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2561 = _GEN_32736 | _GEN_2321; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2562 = _T_402 ? _GEN_2554 : _GEN_2314; // @[sequencer-master.scala 154:24]
  wire  _GEN_2563 = _T_402 ? _GEN_2555 : _GEN_2315; // @[sequencer-master.scala 154:24]
  wire  _GEN_2564 = _T_402 ? _GEN_2556 : _GEN_2316; // @[sequencer-master.scala 154:24]
  wire  _GEN_2565 = _T_402 ? _GEN_2557 : _GEN_2317; // @[sequencer-master.scala 154:24]
  wire  _GEN_2566 = _T_402 ? _GEN_2558 : _GEN_2318; // @[sequencer-master.scala 154:24]
  wire  _GEN_2567 = _T_402 ? _GEN_2559 : _GEN_2319; // @[sequencer-master.scala 154:24]
  wire  _GEN_2568 = _T_402 ? _GEN_2560 : _GEN_2320; // @[sequencer-master.scala 154:24]
  wire  _GEN_2569 = _T_402 ? _GEN_2561 : _GEN_2321; // @[sequencer-master.scala 154:24]
  wire  _GEN_2570 = _GEN_32729 | _GEN_2330; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2571 = _GEN_32730 | _GEN_2331; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2572 = _GEN_32731 | _GEN_2332; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2573 = _GEN_32732 | _GEN_2333; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2574 = _GEN_32733 | _GEN_2334; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2575 = _GEN_32734 | _GEN_2335; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2576 = _GEN_32735 | _GEN_2336; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2577 = _GEN_32736 | _GEN_2337; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2578 = _T_424 ? _GEN_2570 : _GEN_2330; // @[sequencer-master.scala 154:24]
  wire  _GEN_2579 = _T_424 ? _GEN_2571 : _GEN_2331; // @[sequencer-master.scala 154:24]
  wire  _GEN_2580 = _T_424 ? _GEN_2572 : _GEN_2332; // @[sequencer-master.scala 154:24]
  wire  _GEN_2581 = _T_424 ? _GEN_2573 : _GEN_2333; // @[sequencer-master.scala 154:24]
  wire  _GEN_2582 = _T_424 ? _GEN_2574 : _GEN_2334; // @[sequencer-master.scala 154:24]
  wire  _GEN_2583 = _T_424 ? _GEN_2575 : _GEN_2335; // @[sequencer-master.scala 154:24]
  wire  _GEN_2584 = _T_424 ? _GEN_2576 : _GEN_2336; // @[sequencer-master.scala 154:24]
  wire  _GEN_2585 = _T_424 ? _GEN_2577 : _GEN_2337; // @[sequencer-master.scala 154:24]
  wire  _GEN_2586 = _GEN_32729 | _GEN_2346; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2587 = _GEN_32730 | _GEN_2347; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2588 = _GEN_32731 | _GEN_2348; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2589 = _GEN_32732 | _GEN_2349; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2590 = _GEN_32733 | _GEN_2350; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2591 = _GEN_32734 | _GEN_2351; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2592 = _GEN_32735 | _GEN_2352; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2593 = _GEN_32736 | _GEN_2353; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2594 = _T_446 ? _GEN_2586 : _GEN_2346; // @[sequencer-master.scala 154:24]
  wire  _GEN_2595 = _T_446 ? _GEN_2587 : _GEN_2347; // @[sequencer-master.scala 154:24]
  wire  _GEN_2596 = _T_446 ? _GEN_2588 : _GEN_2348; // @[sequencer-master.scala 154:24]
  wire  _GEN_2597 = _T_446 ? _GEN_2589 : _GEN_2349; // @[sequencer-master.scala 154:24]
  wire  _GEN_2598 = _T_446 ? _GEN_2590 : _GEN_2350; // @[sequencer-master.scala 154:24]
  wire  _GEN_2599 = _T_446 ? _GEN_2591 : _GEN_2351; // @[sequencer-master.scala 154:24]
  wire  _GEN_2600 = _T_446 ? _GEN_2592 : _GEN_2352; // @[sequencer-master.scala 154:24]
  wire  _GEN_2601 = _T_446 ? _GEN_2593 : _GEN_2353; // @[sequencer-master.scala 154:24]
  wire  _GEN_2602 = _GEN_32729 | _GEN_2362; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2603 = _GEN_32730 | _GEN_2363; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2604 = _GEN_32731 | _GEN_2364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2605 = _GEN_32732 | _GEN_2365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2606 = _GEN_32733 | _GEN_2366; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2607 = _GEN_32734 | _GEN_2367; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2608 = _GEN_32735 | _GEN_2368; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2609 = _GEN_32736 | _GEN_2369; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2610 = _T_468 ? _GEN_2602 : _GEN_2362; // @[sequencer-master.scala 154:24]
  wire  _GEN_2611 = _T_468 ? _GEN_2603 : _GEN_2363; // @[sequencer-master.scala 154:24]
  wire  _GEN_2612 = _T_468 ? _GEN_2604 : _GEN_2364; // @[sequencer-master.scala 154:24]
  wire  _GEN_2613 = _T_468 ? _GEN_2605 : _GEN_2365; // @[sequencer-master.scala 154:24]
  wire  _GEN_2614 = _T_468 ? _GEN_2606 : _GEN_2366; // @[sequencer-master.scala 154:24]
  wire  _GEN_2615 = _T_468 ? _GEN_2607 : _GEN_2367; // @[sequencer-master.scala 154:24]
  wire  _GEN_2616 = _T_468 ? _GEN_2608 : _GEN_2368; // @[sequencer-master.scala 154:24]
  wire  _GEN_2617 = _T_468 ? _GEN_2609 : _GEN_2369; // @[sequencer-master.scala 154:24]
  wire  _GEN_2618 = _GEN_32729 | _GEN_2378; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2619 = _GEN_32730 | _GEN_2379; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2620 = _GEN_32731 | _GEN_2380; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2621 = _GEN_32732 | _GEN_2381; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2622 = _GEN_32733 | _GEN_2382; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2623 = _GEN_32734 | _GEN_2383; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2624 = _GEN_32735 | _GEN_2384; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2625 = _GEN_32736 | _GEN_2385; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2626 = _T_490 ? _GEN_2618 : _GEN_2378; // @[sequencer-master.scala 154:24]
  wire  _GEN_2627 = _T_490 ? _GEN_2619 : _GEN_2379; // @[sequencer-master.scala 154:24]
  wire  _GEN_2628 = _T_490 ? _GEN_2620 : _GEN_2380; // @[sequencer-master.scala 154:24]
  wire  _GEN_2629 = _T_490 ? _GEN_2621 : _GEN_2381; // @[sequencer-master.scala 154:24]
  wire  _GEN_2630 = _T_490 ? _GEN_2622 : _GEN_2382; // @[sequencer-master.scala 154:24]
  wire  _GEN_2631 = _T_490 ? _GEN_2623 : _GEN_2383; // @[sequencer-master.scala 154:24]
  wire  _GEN_2632 = _T_490 ? _GEN_2624 : _GEN_2384; // @[sequencer-master.scala 154:24]
  wire  _GEN_2633 = _T_490 ? _GEN_2625 : _GEN_2385; // @[sequencer-master.scala 154:24]
  wire  _GEN_2634 = _GEN_32729 | _GEN_2394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2635 = _GEN_32730 | _GEN_2395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2636 = _GEN_32731 | _GEN_2396; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2637 = _GEN_32732 | _GEN_2397; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2638 = _GEN_32733 | _GEN_2398; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2639 = _GEN_32734 | _GEN_2399; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2640 = _GEN_32735 | _GEN_2400; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2641 = _GEN_32736 | _GEN_2401; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2642 = _T_512 ? _GEN_2634 : _GEN_2394; // @[sequencer-master.scala 154:24]
  wire  _GEN_2643 = _T_512 ? _GEN_2635 : _GEN_2395; // @[sequencer-master.scala 154:24]
  wire  _GEN_2644 = _T_512 ? _GEN_2636 : _GEN_2396; // @[sequencer-master.scala 154:24]
  wire  _GEN_2645 = _T_512 ? _GEN_2637 : _GEN_2397; // @[sequencer-master.scala 154:24]
  wire  _GEN_2646 = _T_512 ? _GEN_2638 : _GEN_2398; // @[sequencer-master.scala 154:24]
  wire  _GEN_2647 = _T_512 ? _GEN_2639 : _GEN_2399; // @[sequencer-master.scala 154:24]
  wire  _GEN_2648 = _T_512 ? _GEN_2640 : _GEN_2400; // @[sequencer-master.scala 154:24]
  wire  _GEN_2649 = _T_512 ? _GEN_2641 : _GEN_2401; // @[sequencer-master.scala 154:24]
  wire  _GEN_2650 = _GEN_32729 | _GEN_2410; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2651 = _GEN_32730 | _GEN_2411; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2652 = _GEN_32731 | _GEN_2412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2653 = _GEN_32732 | _GEN_2413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2654 = _GEN_32733 | _GEN_2414; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2655 = _GEN_32734 | _GEN_2415; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2656 = _GEN_32735 | _GEN_2416; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2657 = _GEN_32736 | _GEN_2417; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2658 = _T_534 ? _GEN_2650 : _GEN_2410; // @[sequencer-master.scala 154:24]
  wire  _GEN_2659 = _T_534 ? _GEN_2651 : _GEN_2411; // @[sequencer-master.scala 154:24]
  wire  _GEN_2660 = _T_534 ? _GEN_2652 : _GEN_2412; // @[sequencer-master.scala 154:24]
  wire  _GEN_2661 = _T_534 ? _GEN_2653 : _GEN_2413; // @[sequencer-master.scala 154:24]
  wire  _GEN_2662 = _T_534 ? _GEN_2654 : _GEN_2414; // @[sequencer-master.scala 154:24]
  wire  _GEN_2663 = _T_534 ? _GEN_2655 : _GEN_2415; // @[sequencer-master.scala 154:24]
  wire  _GEN_2664 = _T_534 ? _GEN_2656 : _GEN_2416; // @[sequencer-master.scala 154:24]
  wire  _GEN_2665 = _T_534 ? _GEN_2657 : _GEN_2417; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_2666 = 3'h0 == tail ? io_op_bits_base_vs3_id : e_0_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2667 = 3'h1 == tail ? io_op_bits_base_vs3_id : e_1_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2668 = 3'h2 == tail ? io_op_bits_base_vs3_id : e_2_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2669 = 3'h3 == tail ? io_op_bits_base_vs3_id : e_3_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2670 = 3'h4 == tail ? io_op_bits_base_vs3_id : e_4_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2671 = 3'h5 == tail ? io_op_bits_base_vs3_id : e_5_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2672 = 3'h6 == tail ? io_op_bits_base_vs3_id : e_6_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2673 = 3'h7 == tail ? io_op_bits_base_vs3_id : e_7_base_vs3_id; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2674 = 3'h0 == tail ? io_op_bits_base_vs3_valid : _GEN_1922; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2675 = 3'h1 == tail ? io_op_bits_base_vs3_valid : _GEN_1923; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2676 = 3'h2 == tail ? io_op_bits_base_vs3_valid : _GEN_1924; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2677 = 3'h3 == tail ? io_op_bits_base_vs3_valid : _GEN_1925; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2678 = 3'h4 == tail ? io_op_bits_base_vs3_valid : _GEN_1926; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2679 = 3'h5 == tail ? io_op_bits_base_vs3_valid : _GEN_1927; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2680 = 3'h6 == tail ? io_op_bits_base_vs3_valid : _GEN_1928; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2681 = 3'h7 == tail ? io_op_bits_base_vs3_valid : _GEN_1929; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_2682 = 3'h0 == tail ? io_op_bits_base_vs3_scalar : e_0_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2683 = 3'h1 == tail ? io_op_bits_base_vs3_scalar : e_1_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2684 = 3'h2 == tail ? io_op_bits_base_vs3_scalar : e_2_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2685 = 3'h3 == tail ? io_op_bits_base_vs3_scalar : e_3_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2686 = 3'h4 == tail ? io_op_bits_base_vs3_scalar : e_4_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2687 = 3'h5 == tail ? io_op_bits_base_vs3_scalar : e_5_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2688 = 3'h6 == tail ? io_op_bits_base_vs3_scalar : e_6_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2689 = 3'h7 == tail ? io_op_bits_base_vs3_scalar : e_7_base_vs3_scalar; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2690 = 3'h0 == tail ? io_op_bits_base_vs3_pred : e_0_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2691 = 3'h1 == tail ? io_op_bits_base_vs3_pred : e_1_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2692 = 3'h2 == tail ? io_op_bits_base_vs3_pred : e_2_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2693 = 3'h3 == tail ? io_op_bits_base_vs3_pred : e_3_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2694 = 3'h4 == tail ? io_op_bits_base_vs3_pred : e_4_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2695 = 3'h5 == tail ? io_op_bits_base_vs3_pred : e_5_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2696 = 3'h6 == tail ? io_op_bits_base_vs3_pred : e_6_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire  _GEN_2697 = 3'h7 == tail ? io_op_bits_base_vs3_pred : e_7_base_vs3_pred; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2698 = 3'h0 == tail ? io_op_bits_base_vs3_prec : e_0_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2699 = 3'h1 == tail ? io_op_bits_base_vs3_prec : e_1_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2700 = 3'h2 == tail ? io_op_bits_base_vs3_prec : e_2_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2701 = 3'h3 == tail ? io_op_bits_base_vs3_prec : e_3_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2702 = 3'h4 == tail ? io_op_bits_base_vs3_prec : e_4_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2703 = 3'h5 == tail ? io_op_bits_base_vs3_prec : e_5_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2704 = 3'h6 == tail ? io_op_bits_base_vs3_prec : e_6_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2705 = 3'h7 == tail ? io_op_bits_base_vs3_prec : e_7_base_vs3_prec; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2706 = 3'h0 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2707 = 3'h1 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2708 = 3'h2 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2709 = 3'h3 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2710 = 3'h4 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2711 = 3'h5 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2712 = 3'h6 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2713 = 3'h7 == tail ? io_op_bits_reg_vs3_id : 8'h0; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47 sequencer-master.scala 411:33]
  wire [63:0] _GEN_2714 = 3'h0 == tail ? io_op_bits_sreg_ss3 : e_0_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2715 = 3'h1 == tail ? io_op_bits_sreg_ss3 : e_1_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2716 = 3'h2 == tail ? io_op_bits_sreg_ss3 : e_2_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2717 = 3'h3 == tail ? io_op_bits_sreg_ss3 : e_3_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2718 = 3'h4 == tail ? io_op_bits_sreg_ss3 : e_4_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2719 = 3'h5 == tail ? io_op_bits_sreg_ss3 : e_5_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2720 = 3'h6 == tail ? io_op_bits_sreg_ss3 : e_6_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2721 = 3'h7 == tail ? io_op_bits_sreg_ss3 : e_7_sreg_ss3; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2722 = _T_543 ? _GEN_2714 : e_0_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2723 = _T_543 ? _GEN_2715 : e_1_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2724 = _T_543 ? _GEN_2716 : e_2_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2725 = _T_543 ? _GEN_2717 : e_3_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2726 = _T_543 ? _GEN_2718 : e_4_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2727 = _T_543 ? _GEN_2719 : e_5_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2728 = _T_543 ? _GEN_2720 : e_6_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2729 = _T_543 ? _GEN_2721 : e_7_sreg_ss3; // @[sequencer-master.scala 331:55 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2730 = io_op_bits_base_vs3_valid ? _GEN_2666 : e_0_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2731 = io_op_bits_base_vs3_valid ? _GEN_2667 : e_1_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2732 = io_op_bits_base_vs3_valid ? _GEN_2668 : e_2_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2733 = io_op_bits_base_vs3_valid ? _GEN_2669 : e_3_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2734 = io_op_bits_base_vs3_valid ? _GEN_2670 : e_4_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2735 = io_op_bits_base_vs3_valid ? _GEN_2671 : e_5_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2736 = io_op_bits_base_vs3_valid ? _GEN_2672 : e_6_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2737 = io_op_bits_base_vs3_valid ? _GEN_2673 : e_7_base_vs3_id; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2738 = io_op_bits_base_vs3_valid ? _GEN_2674 : _GEN_1922; // @[sequencer-master.scala 328:47]
  wire  _GEN_2739 = io_op_bits_base_vs3_valid ? _GEN_2675 : _GEN_1923; // @[sequencer-master.scala 328:47]
  wire  _GEN_2740 = io_op_bits_base_vs3_valid ? _GEN_2676 : _GEN_1924; // @[sequencer-master.scala 328:47]
  wire  _GEN_2741 = io_op_bits_base_vs3_valid ? _GEN_2677 : _GEN_1925; // @[sequencer-master.scala 328:47]
  wire  _GEN_2742 = io_op_bits_base_vs3_valid ? _GEN_2678 : _GEN_1926; // @[sequencer-master.scala 328:47]
  wire  _GEN_2743 = io_op_bits_base_vs3_valid ? _GEN_2679 : _GEN_1927; // @[sequencer-master.scala 328:47]
  wire  _GEN_2744 = io_op_bits_base_vs3_valid ? _GEN_2680 : _GEN_1928; // @[sequencer-master.scala 328:47]
  wire  _GEN_2745 = io_op_bits_base_vs3_valid ? _GEN_2681 : _GEN_1929; // @[sequencer-master.scala 328:47]
  wire  _GEN_2746 = io_op_bits_base_vs3_valid ? _GEN_2682 : e_0_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2747 = io_op_bits_base_vs3_valid ? _GEN_2683 : e_1_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2748 = io_op_bits_base_vs3_valid ? _GEN_2684 : e_2_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2749 = io_op_bits_base_vs3_valid ? _GEN_2685 : e_3_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2750 = io_op_bits_base_vs3_valid ? _GEN_2686 : e_4_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2751 = io_op_bits_base_vs3_valid ? _GEN_2687 : e_5_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2752 = io_op_bits_base_vs3_valid ? _GEN_2688 : e_6_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2753 = io_op_bits_base_vs3_valid ? _GEN_2689 : e_7_base_vs3_scalar; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2754 = io_op_bits_base_vs3_valid ? _GEN_2690 : e_0_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2755 = io_op_bits_base_vs3_valid ? _GEN_2691 : e_1_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2756 = io_op_bits_base_vs3_valid ? _GEN_2692 : e_2_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2757 = io_op_bits_base_vs3_valid ? _GEN_2693 : e_3_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2758 = io_op_bits_base_vs3_valid ? _GEN_2694 : e_4_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2759 = io_op_bits_base_vs3_valid ? _GEN_2695 : e_5_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2760 = io_op_bits_base_vs3_valid ? _GEN_2696 : e_6_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2761 = io_op_bits_base_vs3_valid ? _GEN_2697 : e_7_base_vs3_pred; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2762 = io_op_bits_base_vs3_valid ? _GEN_2698 : e_0_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2763 = io_op_bits_base_vs3_valid ? _GEN_2699 : e_1_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2764 = io_op_bits_base_vs3_valid ? _GEN_2700 : e_2_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2765 = io_op_bits_base_vs3_valid ? _GEN_2701 : e_3_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2766 = io_op_bits_base_vs3_valid ? _GEN_2702 : e_4_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2767 = io_op_bits_base_vs3_valid ? _GEN_2703 : e_5_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2768 = io_op_bits_base_vs3_valid ? _GEN_2704 : e_6_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [1:0] _GEN_2769 = io_op_bits_base_vs3_valid ? _GEN_2705 : e_7_base_vs3_prec; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [7:0] _GEN_2770 = io_op_bits_base_vs3_valid ? _GEN_2706 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2771 = io_op_bits_base_vs3_valid ? _GEN_2707 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2772 = io_op_bits_base_vs3_valid ? _GEN_2708 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2773 = io_op_bits_base_vs3_valid ? _GEN_2709 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2774 = io_op_bits_base_vs3_valid ? _GEN_2710 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2775 = io_op_bits_base_vs3_valid ? _GEN_2711 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2776 = io_op_bits_base_vs3_valid ? _GEN_2712 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [7:0] _GEN_2777 = io_op_bits_base_vs3_valid ? _GEN_2713 : 8'h0; // @[sequencer-master.scala 328:47 sequencer-master.scala 411:33]
  wire [63:0] _GEN_2778 = io_op_bits_base_vs3_valid ? _GEN_2722 : e_0_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2779 = io_op_bits_base_vs3_valid ? _GEN_2723 : e_1_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2780 = io_op_bits_base_vs3_valid ? _GEN_2724 : e_2_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2781 = io_op_bits_base_vs3_valid ? _GEN_2725 : e_3_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2782 = io_op_bits_base_vs3_valid ? _GEN_2726 : e_4_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2783 = io_op_bits_base_vs3_valid ? _GEN_2727 : e_5_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2784 = io_op_bits_base_vs3_valid ? _GEN_2728 : e_6_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire [63:0] _GEN_2785 = io_op_bits_base_vs3_valid ? _GEN_2729 : e_7_sreg_ss3; // @[sequencer-master.scala 328:47 sequencer-master.scala 109:14]
  wire  _GEN_2786 = _GEN_32729 | _GEN_2546; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2787 = _GEN_32730 | _GEN_2547; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2788 = _GEN_32731 | _GEN_2548; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2789 = _GEN_32732 | _GEN_2549; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2790 = _GEN_32733 | _GEN_2550; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2791 = _GEN_32734 | _GEN_2551; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2792 = _GEN_32735 | _GEN_2552; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2793 = _GEN_32736 | _GEN_2553; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2794 = _T_557 ? _GEN_2786 : _GEN_2546; // @[sequencer-master.scala 154:24]
  wire  _GEN_2795 = _T_557 ? _GEN_2787 : _GEN_2547; // @[sequencer-master.scala 154:24]
  wire  _GEN_2796 = _T_557 ? _GEN_2788 : _GEN_2548; // @[sequencer-master.scala 154:24]
  wire  _GEN_2797 = _T_557 ? _GEN_2789 : _GEN_2549; // @[sequencer-master.scala 154:24]
  wire  _GEN_2798 = _T_557 ? _GEN_2790 : _GEN_2550; // @[sequencer-master.scala 154:24]
  wire  _GEN_2799 = _T_557 ? _GEN_2791 : _GEN_2551; // @[sequencer-master.scala 154:24]
  wire  _GEN_2800 = _T_557 ? _GEN_2792 : _GEN_2552; // @[sequencer-master.scala 154:24]
  wire  _GEN_2801 = _T_557 ? _GEN_2793 : _GEN_2553; // @[sequencer-master.scala 154:24]
  wire  _GEN_2802 = _GEN_32729 | _GEN_2562; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2803 = _GEN_32730 | _GEN_2563; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2804 = _GEN_32731 | _GEN_2564; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2805 = _GEN_32732 | _GEN_2565; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2806 = _GEN_32733 | _GEN_2566; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2807 = _GEN_32734 | _GEN_2567; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2808 = _GEN_32735 | _GEN_2568; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2809 = _GEN_32736 | _GEN_2569; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2810 = _T_579 ? _GEN_2802 : _GEN_2562; // @[sequencer-master.scala 154:24]
  wire  _GEN_2811 = _T_579 ? _GEN_2803 : _GEN_2563; // @[sequencer-master.scala 154:24]
  wire  _GEN_2812 = _T_579 ? _GEN_2804 : _GEN_2564; // @[sequencer-master.scala 154:24]
  wire  _GEN_2813 = _T_579 ? _GEN_2805 : _GEN_2565; // @[sequencer-master.scala 154:24]
  wire  _GEN_2814 = _T_579 ? _GEN_2806 : _GEN_2566; // @[sequencer-master.scala 154:24]
  wire  _GEN_2815 = _T_579 ? _GEN_2807 : _GEN_2567; // @[sequencer-master.scala 154:24]
  wire  _GEN_2816 = _T_579 ? _GEN_2808 : _GEN_2568; // @[sequencer-master.scala 154:24]
  wire  _GEN_2817 = _T_579 ? _GEN_2809 : _GEN_2569; // @[sequencer-master.scala 154:24]
  wire  _GEN_2818 = _GEN_32729 | _GEN_2578; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2819 = _GEN_32730 | _GEN_2579; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2820 = _GEN_32731 | _GEN_2580; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2821 = _GEN_32732 | _GEN_2581; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2822 = _GEN_32733 | _GEN_2582; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2823 = _GEN_32734 | _GEN_2583; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2824 = _GEN_32735 | _GEN_2584; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2825 = _GEN_32736 | _GEN_2585; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2826 = _T_601 ? _GEN_2818 : _GEN_2578; // @[sequencer-master.scala 154:24]
  wire  _GEN_2827 = _T_601 ? _GEN_2819 : _GEN_2579; // @[sequencer-master.scala 154:24]
  wire  _GEN_2828 = _T_601 ? _GEN_2820 : _GEN_2580; // @[sequencer-master.scala 154:24]
  wire  _GEN_2829 = _T_601 ? _GEN_2821 : _GEN_2581; // @[sequencer-master.scala 154:24]
  wire  _GEN_2830 = _T_601 ? _GEN_2822 : _GEN_2582; // @[sequencer-master.scala 154:24]
  wire  _GEN_2831 = _T_601 ? _GEN_2823 : _GEN_2583; // @[sequencer-master.scala 154:24]
  wire  _GEN_2832 = _T_601 ? _GEN_2824 : _GEN_2584; // @[sequencer-master.scala 154:24]
  wire  _GEN_2833 = _T_601 ? _GEN_2825 : _GEN_2585; // @[sequencer-master.scala 154:24]
  wire  _GEN_2834 = _GEN_32729 | _GEN_2594; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2835 = _GEN_32730 | _GEN_2595; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2836 = _GEN_32731 | _GEN_2596; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2837 = _GEN_32732 | _GEN_2597; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2838 = _GEN_32733 | _GEN_2598; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2839 = _GEN_32734 | _GEN_2599; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2840 = _GEN_32735 | _GEN_2600; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2841 = _GEN_32736 | _GEN_2601; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2842 = _T_623 ? _GEN_2834 : _GEN_2594; // @[sequencer-master.scala 154:24]
  wire  _GEN_2843 = _T_623 ? _GEN_2835 : _GEN_2595; // @[sequencer-master.scala 154:24]
  wire  _GEN_2844 = _T_623 ? _GEN_2836 : _GEN_2596; // @[sequencer-master.scala 154:24]
  wire  _GEN_2845 = _T_623 ? _GEN_2837 : _GEN_2597; // @[sequencer-master.scala 154:24]
  wire  _GEN_2846 = _T_623 ? _GEN_2838 : _GEN_2598; // @[sequencer-master.scala 154:24]
  wire  _GEN_2847 = _T_623 ? _GEN_2839 : _GEN_2599; // @[sequencer-master.scala 154:24]
  wire  _GEN_2848 = _T_623 ? _GEN_2840 : _GEN_2600; // @[sequencer-master.scala 154:24]
  wire  _GEN_2849 = _T_623 ? _GEN_2841 : _GEN_2601; // @[sequencer-master.scala 154:24]
  wire  _GEN_2850 = _GEN_32729 | _GEN_2610; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2851 = _GEN_32730 | _GEN_2611; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2852 = _GEN_32731 | _GEN_2612; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2853 = _GEN_32732 | _GEN_2613; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2854 = _GEN_32733 | _GEN_2614; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2855 = _GEN_32734 | _GEN_2615; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2856 = _GEN_32735 | _GEN_2616; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2857 = _GEN_32736 | _GEN_2617; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2858 = _T_645 ? _GEN_2850 : _GEN_2610; // @[sequencer-master.scala 154:24]
  wire  _GEN_2859 = _T_645 ? _GEN_2851 : _GEN_2611; // @[sequencer-master.scala 154:24]
  wire  _GEN_2860 = _T_645 ? _GEN_2852 : _GEN_2612; // @[sequencer-master.scala 154:24]
  wire  _GEN_2861 = _T_645 ? _GEN_2853 : _GEN_2613; // @[sequencer-master.scala 154:24]
  wire  _GEN_2862 = _T_645 ? _GEN_2854 : _GEN_2614; // @[sequencer-master.scala 154:24]
  wire  _GEN_2863 = _T_645 ? _GEN_2855 : _GEN_2615; // @[sequencer-master.scala 154:24]
  wire  _GEN_2864 = _T_645 ? _GEN_2856 : _GEN_2616; // @[sequencer-master.scala 154:24]
  wire  _GEN_2865 = _T_645 ? _GEN_2857 : _GEN_2617; // @[sequencer-master.scala 154:24]
  wire  _GEN_2866 = _GEN_32729 | _GEN_2626; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2867 = _GEN_32730 | _GEN_2627; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2868 = _GEN_32731 | _GEN_2628; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2869 = _GEN_32732 | _GEN_2629; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2870 = _GEN_32733 | _GEN_2630; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2871 = _GEN_32734 | _GEN_2631; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2872 = _GEN_32735 | _GEN_2632; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2873 = _GEN_32736 | _GEN_2633; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2874 = _T_667 ? _GEN_2866 : _GEN_2626; // @[sequencer-master.scala 154:24]
  wire  _GEN_2875 = _T_667 ? _GEN_2867 : _GEN_2627; // @[sequencer-master.scala 154:24]
  wire  _GEN_2876 = _T_667 ? _GEN_2868 : _GEN_2628; // @[sequencer-master.scala 154:24]
  wire  _GEN_2877 = _T_667 ? _GEN_2869 : _GEN_2629; // @[sequencer-master.scala 154:24]
  wire  _GEN_2878 = _T_667 ? _GEN_2870 : _GEN_2630; // @[sequencer-master.scala 154:24]
  wire  _GEN_2879 = _T_667 ? _GEN_2871 : _GEN_2631; // @[sequencer-master.scala 154:24]
  wire  _GEN_2880 = _T_667 ? _GEN_2872 : _GEN_2632; // @[sequencer-master.scala 154:24]
  wire  _GEN_2881 = _T_667 ? _GEN_2873 : _GEN_2633; // @[sequencer-master.scala 154:24]
  wire  _GEN_2882 = _GEN_32729 | _GEN_2642; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2883 = _GEN_32730 | _GEN_2643; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2884 = _GEN_32731 | _GEN_2644; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2885 = _GEN_32732 | _GEN_2645; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2886 = _GEN_32733 | _GEN_2646; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2887 = _GEN_32734 | _GEN_2647; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2888 = _GEN_32735 | _GEN_2648; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2889 = _GEN_32736 | _GEN_2649; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2890 = _T_689 ? _GEN_2882 : _GEN_2642; // @[sequencer-master.scala 154:24]
  wire  _GEN_2891 = _T_689 ? _GEN_2883 : _GEN_2643; // @[sequencer-master.scala 154:24]
  wire  _GEN_2892 = _T_689 ? _GEN_2884 : _GEN_2644; // @[sequencer-master.scala 154:24]
  wire  _GEN_2893 = _T_689 ? _GEN_2885 : _GEN_2645; // @[sequencer-master.scala 154:24]
  wire  _GEN_2894 = _T_689 ? _GEN_2886 : _GEN_2646; // @[sequencer-master.scala 154:24]
  wire  _GEN_2895 = _T_689 ? _GEN_2887 : _GEN_2647; // @[sequencer-master.scala 154:24]
  wire  _GEN_2896 = _T_689 ? _GEN_2888 : _GEN_2648; // @[sequencer-master.scala 154:24]
  wire  _GEN_2897 = _T_689 ? _GEN_2889 : _GEN_2649; // @[sequencer-master.scala 154:24]
  wire  _GEN_2898 = _GEN_32729 | _GEN_2658; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2899 = _GEN_32730 | _GEN_2659; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2900 = _GEN_32731 | _GEN_2660; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2901 = _GEN_32732 | _GEN_2661; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2902 = _GEN_32733 | _GEN_2662; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2903 = _GEN_32734 | _GEN_2663; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2904 = _GEN_32735 | _GEN_2664; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2905 = _GEN_32736 | _GEN_2665; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_2906 = _T_711 ? _GEN_2898 : _GEN_2658; // @[sequencer-master.scala 154:24]
  wire  _GEN_2907 = _T_711 ? _GEN_2899 : _GEN_2659; // @[sequencer-master.scala 154:24]
  wire  _GEN_2908 = _T_711 ? _GEN_2900 : _GEN_2660; // @[sequencer-master.scala 154:24]
  wire  _GEN_2909 = _T_711 ? _GEN_2901 : _GEN_2661; // @[sequencer-master.scala 154:24]
  wire  _GEN_2910 = _T_711 ? _GEN_2902 : _GEN_2662; // @[sequencer-master.scala 154:24]
  wire  _GEN_2911 = _T_711 ? _GEN_2903 : _GEN_2663; // @[sequencer-master.scala 154:24]
  wire  _GEN_2912 = _T_711 ? _GEN_2904 : _GEN_2664; // @[sequencer-master.scala 154:24]
  wire  _GEN_2913 = _T_711 ? _GEN_2905 : _GEN_2665; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_2914 = 3'h0 == tail ? io_op_bits_base_vd_id : _GEN_1816; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2915 = 3'h1 == tail ? io_op_bits_base_vd_id : _GEN_1817; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2916 = 3'h2 == tail ? io_op_bits_base_vd_id : _GEN_1818; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2917 = 3'h3 == tail ? io_op_bits_base_vd_id : _GEN_1819; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2918 = 3'h4 == tail ? io_op_bits_base_vd_id : _GEN_1820; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2919 = 3'h5 == tail ? io_op_bits_base_vd_id : _GEN_1821; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2920 = 3'h6 == tail ? io_op_bits_base_vd_id : _GEN_1822; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2921 = 3'h7 == tail ? io_op_bits_base_vd_id : _GEN_1823; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2922 = 3'h0 == tail ? io_op_bits_base_vd_valid : _GEN_1930; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2923 = 3'h1 == tail ? io_op_bits_base_vd_valid : _GEN_1931; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2924 = 3'h2 == tail ? io_op_bits_base_vd_valid : _GEN_1932; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2925 = 3'h3 == tail ? io_op_bits_base_vd_valid : _GEN_1933; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2926 = 3'h4 == tail ? io_op_bits_base_vd_valid : _GEN_1934; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2927 = 3'h5 == tail ? io_op_bits_base_vd_valid : _GEN_1935; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2928 = 3'h6 == tail ? io_op_bits_base_vd_valid : _GEN_1936; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2929 = 3'h7 == tail ? io_op_bits_base_vd_valid : _GEN_1937; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2930 = 3'h0 == tail ? io_op_bits_base_vd_scalar : _GEN_1824; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2931 = 3'h1 == tail ? io_op_bits_base_vd_scalar : _GEN_1825; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2932 = 3'h2 == tail ? io_op_bits_base_vd_scalar : _GEN_1826; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2933 = 3'h3 == tail ? io_op_bits_base_vd_scalar : _GEN_1827; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2934 = 3'h4 == tail ? io_op_bits_base_vd_scalar : _GEN_1828; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2935 = 3'h5 == tail ? io_op_bits_base_vd_scalar : _GEN_1829; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2936 = 3'h6 == tail ? io_op_bits_base_vd_scalar : _GEN_1830; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2937 = 3'h7 == tail ? io_op_bits_base_vd_scalar : _GEN_1831; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2938 = 3'h0 == tail ? io_op_bits_base_vd_pred : _GEN_1832; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2939 = 3'h1 == tail ? io_op_bits_base_vd_pred : _GEN_1833; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2940 = 3'h2 == tail ? io_op_bits_base_vd_pred : _GEN_1834; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2941 = 3'h3 == tail ? io_op_bits_base_vd_pred : _GEN_1835; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2942 = 3'h4 == tail ? io_op_bits_base_vd_pred : _GEN_1836; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2943 = 3'h5 == tail ? io_op_bits_base_vd_pred : _GEN_1837; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2944 = 3'h6 == tail ? io_op_bits_base_vd_pred : _GEN_1838; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_2945 = 3'h7 == tail ? io_op_bits_base_vd_pred : _GEN_1839; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2946 = 3'h0 == tail ? io_op_bits_base_vd_prec : _GEN_1840; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2947 = 3'h1 == tail ? io_op_bits_base_vd_prec : _GEN_1841; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2948 = 3'h2 == tail ? io_op_bits_base_vd_prec : _GEN_1842; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2949 = 3'h3 == tail ? io_op_bits_base_vd_prec : _GEN_1843; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2950 = 3'h4 == tail ? io_op_bits_base_vd_prec : _GEN_1844; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2951 = 3'h5 == tail ? io_op_bits_base_vd_prec : _GEN_1845; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2952 = 3'h6 == tail ? io_op_bits_base_vd_prec : _GEN_1846; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_2953 = 3'h7 == tail ? io_op_bits_base_vd_prec : _GEN_1847; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_2954 = 3'h0 == tail ? io_op_bits_reg_vd_id : _GEN_1848; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2955 = 3'h1 == tail ? io_op_bits_reg_vd_id : _GEN_1849; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2956 = 3'h2 == tail ? io_op_bits_reg_vd_id : _GEN_1850; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2957 = 3'h3 == tail ? io_op_bits_reg_vd_id : _GEN_1851; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2958 = 3'h4 == tail ? io_op_bits_reg_vd_id : _GEN_1852; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2959 = 3'h5 == tail ? io_op_bits_reg_vd_id : _GEN_1853; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2960 = 3'h6 == tail ? io_op_bits_reg_vd_id : _GEN_1854; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2961 = 3'h7 == tail ? io_op_bits_reg_vd_id : _GEN_1855; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_2962 = io_op_bits_base_vd_valid ? _GEN_2914 : _GEN_1816; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2963 = io_op_bits_base_vd_valid ? _GEN_2915 : _GEN_1817; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2964 = io_op_bits_base_vd_valid ? _GEN_2916 : _GEN_1818; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2965 = io_op_bits_base_vd_valid ? _GEN_2917 : _GEN_1819; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2966 = io_op_bits_base_vd_valid ? _GEN_2918 : _GEN_1820; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2967 = io_op_bits_base_vd_valid ? _GEN_2919 : _GEN_1821; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2968 = io_op_bits_base_vd_valid ? _GEN_2920 : _GEN_1822; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_2969 = io_op_bits_base_vd_valid ? _GEN_2921 : _GEN_1823; // @[sequencer-master.scala 362:41]
  wire  _GEN_2970 = io_op_bits_base_vd_valid ? _GEN_2922 : _GEN_1930; // @[sequencer-master.scala 362:41]
  wire  _GEN_2971 = io_op_bits_base_vd_valid ? _GEN_2923 : _GEN_1931; // @[sequencer-master.scala 362:41]
  wire  _GEN_2972 = io_op_bits_base_vd_valid ? _GEN_2924 : _GEN_1932; // @[sequencer-master.scala 362:41]
  wire  _GEN_2973 = io_op_bits_base_vd_valid ? _GEN_2925 : _GEN_1933; // @[sequencer-master.scala 362:41]
  wire  _GEN_2974 = io_op_bits_base_vd_valid ? _GEN_2926 : _GEN_1934; // @[sequencer-master.scala 362:41]
  wire  _GEN_2975 = io_op_bits_base_vd_valid ? _GEN_2927 : _GEN_1935; // @[sequencer-master.scala 362:41]
  wire  _GEN_2976 = io_op_bits_base_vd_valid ? _GEN_2928 : _GEN_1936; // @[sequencer-master.scala 362:41]
  wire  _GEN_2977 = io_op_bits_base_vd_valid ? _GEN_2929 : _GEN_1937; // @[sequencer-master.scala 362:41]
  wire  _GEN_2978 = io_op_bits_base_vd_valid ? _GEN_2930 : _GEN_1824; // @[sequencer-master.scala 362:41]
  wire  _GEN_2979 = io_op_bits_base_vd_valid ? _GEN_2931 : _GEN_1825; // @[sequencer-master.scala 362:41]
  wire  _GEN_2980 = io_op_bits_base_vd_valid ? _GEN_2932 : _GEN_1826; // @[sequencer-master.scala 362:41]
  wire  _GEN_2981 = io_op_bits_base_vd_valid ? _GEN_2933 : _GEN_1827; // @[sequencer-master.scala 362:41]
  wire  _GEN_2982 = io_op_bits_base_vd_valid ? _GEN_2934 : _GEN_1828; // @[sequencer-master.scala 362:41]
  wire  _GEN_2983 = io_op_bits_base_vd_valid ? _GEN_2935 : _GEN_1829; // @[sequencer-master.scala 362:41]
  wire  _GEN_2984 = io_op_bits_base_vd_valid ? _GEN_2936 : _GEN_1830; // @[sequencer-master.scala 362:41]
  wire  _GEN_2985 = io_op_bits_base_vd_valid ? _GEN_2937 : _GEN_1831; // @[sequencer-master.scala 362:41]
  wire  _GEN_2986 = io_op_bits_base_vd_valid ? _GEN_2938 : _GEN_1832; // @[sequencer-master.scala 362:41]
  wire  _GEN_2987 = io_op_bits_base_vd_valid ? _GEN_2939 : _GEN_1833; // @[sequencer-master.scala 362:41]
  wire  _GEN_2988 = io_op_bits_base_vd_valid ? _GEN_2940 : _GEN_1834; // @[sequencer-master.scala 362:41]
  wire  _GEN_2989 = io_op_bits_base_vd_valid ? _GEN_2941 : _GEN_1835; // @[sequencer-master.scala 362:41]
  wire  _GEN_2990 = io_op_bits_base_vd_valid ? _GEN_2942 : _GEN_1836; // @[sequencer-master.scala 362:41]
  wire  _GEN_2991 = io_op_bits_base_vd_valid ? _GEN_2943 : _GEN_1837; // @[sequencer-master.scala 362:41]
  wire  _GEN_2992 = io_op_bits_base_vd_valid ? _GEN_2944 : _GEN_1838; // @[sequencer-master.scala 362:41]
  wire  _GEN_2993 = io_op_bits_base_vd_valid ? _GEN_2945 : _GEN_1839; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_2994 = io_op_bits_base_vd_valid ? _GEN_2946 : _GEN_1840; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_2995 = io_op_bits_base_vd_valid ? _GEN_2947 : _GEN_1841; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_2996 = io_op_bits_base_vd_valid ? _GEN_2948 : _GEN_1842; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_2997 = io_op_bits_base_vd_valid ? _GEN_2949 : _GEN_1843; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_2998 = io_op_bits_base_vd_valid ? _GEN_2950 : _GEN_1844; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_2999 = io_op_bits_base_vd_valid ? _GEN_2951 : _GEN_1845; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_3000 = io_op_bits_base_vd_valid ? _GEN_2952 : _GEN_1846; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_3001 = io_op_bits_base_vd_valid ? _GEN_2953 : _GEN_1847; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3002 = io_op_bits_base_vd_valid ? _GEN_2954 : _GEN_1848; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3003 = io_op_bits_base_vd_valid ? _GEN_2955 : _GEN_1849; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3004 = io_op_bits_base_vd_valid ? _GEN_2956 : _GEN_1850; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3005 = io_op_bits_base_vd_valid ? _GEN_2957 : _GEN_1851; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3006 = io_op_bits_base_vd_valid ? _GEN_2958 : _GEN_1852; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3007 = io_op_bits_base_vd_valid ? _GEN_2959 : _GEN_1853; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3008 = io_op_bits_base_vd_valid ? _GEN_2960 : _GEN_1854; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_3009 = io_op_bits_base_vd_valid ? _GEN_2961 : _GEN_1855; // @[sequencer-master.scala 362:41]
  wire  _GEN_3010 = _GEN_32729 | _GEN_1954; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3011 = _GEN_32730 | _GEN_1955; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3012 = _GEN_32731 | _GEN_1956; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3013 = _GEN_32732 | _GEN_1957; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3014 = _GEN_32733 | _GEN_1958; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3015 = _GEN_32734 | _GEN_1959; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3016 = _GEN_32735 | _GEN_1960; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3017 = _GEN_32736 | _GEN_1961; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3018 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3010 : _GEN_1954; // @[sequencer-master.scala 161:86]
  wire  _GEN_3019 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3011 : _GEN_1955; // @[sequencer-master.scala 161:86]
  wire  _GEN_3020 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3012 : _GEN_1956; // @[sequencer-master.scala 161:86]
  wire  _GEN_3021 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3013 : _GEN_1957; // @[sequencer-master.scala 161:86]
  wire  _GEN_3022 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3014 : _GEN_1958; // @[sequencer-master.scala 161:86]
  wire  _GEN_3023 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3015 : _GEN_1959; // @[sequencer-master.scala 161:86]
  wire  _GEN_3024 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3016 : _GEN_1960; // @[sequencer-master.scala 161:86]
  wire  _GEN_3025 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_3017 : _GEN_1961; // @[sequencer-master.scala 161:86]
  wire  _GEN_3026 = _GEN_32729 | _GEN_1978; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3027 = _GEN_32730 | _GEN_1979; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3028 = _GEN_32731 | _GEN_1980; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3029 = _GEN_32732 | _GEN_1981; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3030 = _GEN_32733 | _GEN_1982; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3031 = _GEN_32734 | _GEN_1983; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3032 = _GEN_32735 | _GEN_1984; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3033 = _GEN_32736 | _GEN_1985; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3034 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3026 : _GEN_1978; // @[sequencer-master.scala 161:86]
  wire  _GEN_3035 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3027 : _GEN_1979; // @[sequencer-master.scala 161:86]
  wire  _GEN_3036 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3028 : _GEN_1980; // @[sequencer-master.scala 161:86]
  wire  _GEN_3037 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3029 : _GEN_1981; // @[sequencer-master.scala 161:86]
  wire  _GEN_3038 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3030 : _GEN_1982; // @[sequencer-master.scala 161:86]
  wire  _GEN_3039 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3031 : _GEN_1983; // @[sequencer-master.scala 161:86]
  wire  _GEN_3040 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3032 : _GEN_1984; // @[sequencer-master.scala 161:86]
  wire  _GEN_3041 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_3033 : _GEN_1985; // @[sequencer-master.scala 161:86]
  wire  _GEN_3042 = _GEN_32729 | _GEN_2002; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3043 = _GEN_32730 | _GEN_2003; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3044 = _GEN_32731 | _GEN_2004; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3045 = _GEN_32732 | _GEN_2005; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3046 = _GEN_32733 | _GEN_2006; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3047 = _GEN_32734 | _GEN_2007; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3048 = _GEN_32735 | _GEN_2008; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3049 = _GEN_32736 | _GEN_2009; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3050 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3042 : _GEN_2002; // @[sequencer-master.scala 161:86]
  wire  _GEN_3051 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3043 : _GEN_2003; // @[sequencer-master.scala 161:86]
  wire  _GEN_3052 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3044 : _GEN_2004; // @[sequencer-master.scala 161:86]
  wire  _GEN_3053 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3045 : _GEN_2005; // @[sequencer-master.scala 161:86]
  wire  _GEN_3054 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3046 : _GEN_2006; // @[sequencer-master.scala 161:86]
  wire  _GEN_3055 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3047 : _GEN_2007; // @[sequencer-master.scala 161:86]
  wire  _GEN_3056 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3048 : _GEN_2008; // @[sequencer-master.scala 161:86]
  wire  _GEN_3057 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_3049 : _GEN_2009; // @[sequencer-master.scala 161:86]
  wire  _GEN_3058 = _GEN_32729 | _GEN_2026; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3059 = _GEN_32730 | _GEN_2027; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3060 = _GEN_32731 | _GEN_2028; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3061 = _GEN_32732 | _GEN_2029; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3062 = _GEN_32733 | _GEN_2030; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3063 = _GEN_32734 | _GEN_2031; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3064 = _GEN_32735 | _GEN_2032; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3065 = _GEN_32736 | _GEN_2033; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3066 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3058 : _GEN_2026; // @[sequencer-master.scala 161:86]
  wire  _GEN_3067 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3059 : _GEN_2027; // @[sequencer-master.scala 161:86]
  wire  _GEN_3068 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3060 : _GEN_2028; // @[sequencer-master.scala 161:86]
  wire  _GEN_3069 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3061 : _GEN_2029; // @[sequencer-master.scala 161:86]
  wire  _GEN_3070 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3062 : _GEN_2030; // @[sequencer-master.scala 161:86]
  wire  _GEN_3071 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3063 : _GEN_2031; // @[sequencer-master.scala 161:86]
  wire  _GEN_3072 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3064 : _GEN_2032; // @[sequencer-master.scala 161:86]
  wire  _GEN_3073 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_3065 : _GEN_2033; // @[sequencer-master.scala 161:86]
  wire  _GEN_3074 = _GEN_32729 | _GEN_2050; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3075 = _GEN_32730 | _GEN_2051; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3076 = _GEN_32731 | _GEN_2052; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3077 = _GEN_32732 | _GEN_2053; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3078 = _GEN_32733 | _GEN_2054; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3079 = _GEN_32734 | _GEN_2055; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3080 = _GEN_32735 | _GEN_2056; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3081 = _GEN_32736 | _GEN_2057; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3082 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3074 : _GEN_2050; // @[sequencer-master.scala 161:86]
  wire  _GEN_3083 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3075 : _GEN_2051; // @[sequencer-master.scala 161:86]
  wire  _GEN_3084 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3076 : _GEN_2052; // @[sequencer-master.scala 161:86]
  wire  _GEN_3085 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3077 : _GEN_2053; // @[sequencer-master.scala 161:86]
  wire  _GEN_3086 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3078 : _GEN_2054; // @[sequencer-master.scala 161:86]
  wire  _GEN_3087 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3079 : _GEN_2055; // @[sequencer-master.scala 161:86]
  wire  _GEN_3088 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3080 : _GEN_2056; // @[sequencer-master.scala 161:86]
  wire  _GEN_3089 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_3081 : _GEN_2057; // @[sequencer-master.scala 161:86]
  wire  _GEN_3090 = _GEN_32729 | _GEN_2074; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3091 = _GEN_32730 | _GEN_2075; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3092 = _GEN_32731 | _GEN_2076; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3093 = _GEN_32732 | _GEN_2077; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3094 = _GEN_32733 | _GEN_2078; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3095 = _GEN_32734 | _GEN_2079; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3096 = _GEN_32735 | _GEN_2080; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3097 = _GEN_32736 | _GEN_2081; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3098 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3090 : _GEN_2074; // @[sequencer-master.scala 161:86]
  wire  _GEN_3099 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3091 : _GEN_2075; // @[sequencer-master.scala 161:86]
  wire  _GEN_3100 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3092 : _GEN_2076; // @[sequencer-master.scala 161:86]
  wire  _GEN_3101 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3093 : _GEN_2077; // @[sequencer-master.scala 161:86]
  wire  _GEN_3102 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3094 : _GEN_2078; // @[sequencer-master.scala 161:86]
  wire  _GEN_3103 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3095 : _GEN_2079; // @[sequencer-master.scala 161:86]
  wire  _GEN_3104 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3096 : _GEN_2080; // @[sequencer-master.scala 161:86]
  wire  _GEN_3105 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_3097 : _GEN_2081; // @[sequencer-master.scala 161:86]
  wire  _GEN_3106 = _GEN_32729 | _GEN_2098; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3107 = _GEN_32730 | _GEN_2099; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3108 = _GEN_32731 | _GEN_2100; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3109 = _GEN_32732 | _GEN_2101; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3110 = _GEN_32733 | _GEN_2102; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3111 = _GEN_32734 | _GEN_2103; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3112 = _GEN_32735 | _GEN_2104; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3113 = _GEN_32736 | _GEN_2105; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3114 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3106 : _GEN_2098; // @[sequencer-master.scala 161:86]
  wire  _GEN_3115 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3107 : _GEN_2099; // @[sequencer-master.scala 161:86]
  wire  _GEN_3116 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3108 : _GEN_2100; // @[sequencer-master.scala 161:86]
  wire  _GEN_3117 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3109 : _GEN_2101; // @[sequencer-master.scala 161:86]
  wire  _GEN_3118 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3110 : _GEN_2102; // @[sequencer-master.scala 161:86]
  wire  _GEN_3119 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3111 : _GEN_2103; // @[sequencer-master.scala 161:86]
  wire  _GEN_3120 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3112 : _GEN_2104; // @[sequencer-master.scala 161:86]
  wire  _GEN_3121 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_3113 : _GEN_2105; // @[sequencer-master.scala 161:86]
  wire  _GEN_3122 = _GEN_32729 | _GEN_2122; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3123 = _GEN_32730 | _GEN_2123; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3124 = _GEN_32731 | _GEN_2124; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3125 = _GEN_32732 | _GEN_2125; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3126 = _GEN_32733 | _GEN_2126; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3127 = _GEN_32734 | _GEN_2127; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3128 = _GEN_32735 | _GEN_2128; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3129 = _GEN_32736 | _GEN_2129; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_3130 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3122 : _GEN_2122; // @[sequencer-master.scala 161:86]
  wire  _GEN_3131 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3123 : _GEN_2123; // @[sequencer-master.scala 161:86]
  wire  _GEN_3132 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3124 : _GEN_2124; // @[sequencer-master.scala 161:86]
  wire  _GEN_3133 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3125 : _GEN_2125; // @[sequencer-master.scala 161:86]
  wire  _GEN_3134 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3126 : _GEN_2126; // @[sequencer-master.scala 161:86]
  wire  _GEN_3135 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3127 : _GEN_2127; // @[sequencer-master.scala 161:86]
  wire  _GEN_3136 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3128 : _GEN_2128; // @[sequencer-master.scala 161:86]
  wire  _GEN_3137 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_3129 : _GEN_2129; // @[sequencer-master.scala 161:86]
  wire  _GEN_3138 = _GEN_32729 | _GEN_1962; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3139 = _GEN_32730 | _GEN_1963; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3140 = _GEN_32731 | _GEN_1964; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3141 = _GEN_32732 | _GEN_1965; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3142 = _GEN_32733 | _GEN_1966; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3143 = _GEN_32734 | _GEN_1967; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3144 = _GEN_32735 | _GEN_1968; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3145 = _GEN_32736 | _GEN_1969; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3146 = _T_1442 ? _GEN_3138 : _GEN_1962; // @[sequencer-master.scala 168:32]
  wire  _GEN_3147 = _T_1442 ? _GEN_3139 : _GEN_1963; // @[sequencer-master.scala 168:32]
  wire  _GEN_3148 = _T_1442 ? _GEN_3140 : _GEN_1964; // @[sequencer-master.scala 168:32]
  wire  _GEN_3149 = _T_1442 ? _GEN_3141 : _GEN_1965; // @[sequencer-master.scala 168:32]
  wire  _GEN_3150 = _T_1442 ? _GEN_3142 : _GEN_1966; // @[sequencer-master.scala 168:32]
  wire  _GEN_3151 = _T_1442 ? _GEN_3143 : _GEN_1967; // @[sequencer-master.scala 168:32]
  wire  _GEN_3152 = _T_1442 ? _GEN_3144 : _GEN_1968; // @[sequencer-master.scala 168:32]
  wire  _GEN_3153 = _T_1442 ? _GEN_3145 : _GEN_1969; // @[sequencer-master.scala 168:32]
  wire  _GEN_3154 = _GEN_32729 | _GEN_1986; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3155 = _GEN_32730 | _GEN_1987; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3156 = _GEN_32731 | _GEN_1988; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3157 = _GEN_32732 | _GEN_1989; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3158 = _GEN_32733 | _GEN_1990; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3159 = _GEN_32734 | _GEN_1991; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3160 = _GEN_32735 | _GEN_1992; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3161 = _GEN_32736 | _GEN_1993; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3162 = _T_1464 ? _GEN_3154 : _GEN_1986; // @[sequencer-master.scala 168:32]
  wire  _GEN_3163 = _T_1464 ? _GEN_3155 : _GEN_1987; // @[sequencer-master.scala 168:32]
  wire  _GEN_3164 = _T_1464 ? _GEN_3156 : _GEN_1988; // @[sequencer-master.scala 168:32]
  wire  _GEN_3165 = _T_1464 ? _GEN_3157 : _GEN_1989; // @[sequencer-master.scala 168:32]
  wire  _GEN_3166 = _T_1464 ? _GEN_3158 : _GEN_1990; // @[sequencer-master.scala 168:32]
  wire  _GEN_3167 = _T_1464 ? _GEN_3159 : _GEN_1991; // @[sequencer-master.scala 168:32]
  wire  _GEN_3168 = _T_1464 ? _GEN_3160 : _GEN_1992; // @[sequencer-master.scala 168:32]
  wire  _GEN_3169 = _T_1464 ? _GEN_3161 : _GEN_1993; // @[sequencer-master.scala 168:32]
  wire  _GEN_3170 = _GEN_32729 | _GEN_2010; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3171 = _GEN_32730 | _GEN_2011; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3172 = _GEN_32731 | _GEN_2012; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3173 = _GEN_32732 | _GEN_2013; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3174 = _GEN_32733 | _GEN_2014; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3175 = _GEN_32734 | _GEN_2015; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3176 = _GEN_32735 | _GEN_2016; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3177 = _GEN_32736 | _GEN_2017; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3178 = _T_1486 ? _GEN_3170 : _GEN_2010; // @[sequencer-master.scala 168:32]
  wire  _GEN_3179 = _T_1486 ? _GEN_3171 : _GEN_2011; // @[sequencer-master.scala 168:32]
  wire  _GEN_3180 = _T_1486 ? _GEN_3172 : _GEN_2012; // @[sequencer-master.scala 168:32]
  wire  _GEN_3181 = _T_1486 ? _GEN_3173 : _GEN_2013; // @[sequencer-master.scala 168:32]
  wire  _GEN_3182 = _T_1486 ? _GEN_3174 : _GEN_2014; // @[sequencer-master.scala 168:32]
  wire  _GEN_3183 = _T_1486 ? _GEN_3175 : _GEN_2015; // @[sequencer-master.scala 168:32]
  wire  _GEN_3184 = _T_1486 ? _GEN_3176 : _GEN_2016; // @[sequencer-master.scala 168:32]
  wire  _GEN_3185 = _T_1486 ? _GEN_3177 : _GEN_2017; // @[sequencer-master.scala 168:32]
  wire  _GEN_3186 = _GEN_32729 | _GEN_2034; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3187 = _GEN_32730 | _GEN_2035; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3188 = _GEN_32731 | _GEN_2036; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3189 = _GEN_32732 | _GEN_2037; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3190 = _GEN_32733 | _GEN_2038; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3191 = _GEN_32734 | _GEN_2039; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3192 = _GEN_32735 | _GEN_2040; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3193 = _GEN_32736 | _GEN_2041; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3194 = _T_1508 ? _GEN_3186 : _GEN_2034; // @[sequencer-master.scala 168:32]
  wire  _GEN_3195 = _T_1508 ? _GEN_3187 : _GEN_2035; // @[sequencer-master.scala 168:32]
  wire  _GEN_3196 = _T_1508 ? _GEN_3188 : _GEN_2036; // @[sequencer-master.scala 168:32]
  wire  _GEN_3197 = _T_1508 ? _GEN_3189 : _GEN_2037; // @[sequencer-master.scala 168:32]
  wire  _GEN_3198 = _T_1508 ? _GEN_3190 : _GEN_2038; // @[sequencer-master.scala 168:32]
  wire  _GEN_3199 = _T_1508 ? _GEN_3191 : _GEN_2039; // @[sequencer-master.scala 168:32]
  wire  _GEN_3200 = _T_1508 ? _GEN_3192 : _GEN_2040; // @[sequencer-master.scala 168:32]
  wire  _GEN_3201 = _T_1508 ? _GEN_3193 : _GEN_2041; // @[sequencer-master.scala 168:32]
  wire  _GEN_3202 = _GEN_32729 | _GEN_2058; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3203 = _GEN_32730 | _GEN_2059; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3204 = _GEN_32731 | _GEN_2060; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3205 = _GEN_32732 | _GEN_2061; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3206 = _GEN_32733 | _GEN_2062; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3207 = _GEN_32734 | _GEN_2063; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3208 = _GEN_32735 | _GEN_2064; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3209 = _GEN_32736 | _GEN_2065; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3210 = _T_1530 ? _GEN_3202 : _GEN_2058; // @[sequencer-master.scala 168:32]
  wire  _GEN_3211 = _T_1530 ? _GEN_3203 : _GEN_2059; // @[sequencer-master.scala 168:32]
  wire  _GEN_3212 = _T_1530 ? _GEN_3204 : _GEN_2060; // @[sequencer-master.scala 168:32]
  wire  _GEN_3213 = _T_1530 ? _GEN_3205 : _GEN_2061; // @[sequencer-master.scala 168:32]
  wire  _GEN_3214 = _T_1530 ? _GEN_3206 : _GEN_2062; // @[sequencer-master.scala 168:32]
  wire  _GEN_3215 = _T_1530 ? _GEN_3207 : _GEN_2063; // @[sequencer-master.scala 168:32]
  wire  _GEN_3216 = _T_1530 ? _GEN_3208 : _GEN_2064; // @[sequencer-master.scala 168:32]
  wire  _GEN_3217 = _T_1530 ? _GEN_3209 : _GEN_2065; // @[sequencer-master.scala 168:32]
  wire  _GEN_3218 = _GEN_32729 | _GEN_2082; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3219 = _GEN_32730 | _GEN_2083; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3220 = _GEN_32731 | _GEN_2084; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3221 = _GEN_32732 | _GEN_2085; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3222 = _GEN_32733 | _GEN_2086; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3223 = _GEN_32734 | _GEN_2087; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3224 = _GEN_32735 | _GEN_2088; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3225 = _GEN_32736 | _GEN_2089; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3226 = _T_1552 ? _GEN_3218 : _GEN_2082; // @[sequencer-master.scala 168:32]
  wire  _GEN_3227 = _T_1552 ? _GEN_3219 : _GEN_2083; // @[sequencer-master.scala 168:32]
  wire  _GEN_3228 = _T_1552 ? _GEN_3220 : _GEN_2084; // @[sequencer-master.scala 168:32]
  wire  _GEN_3229 = _T_1552 ? _GEN_3221 : _GEN_2085; // @[sequencer-master.scala 168:32]
  wire  _GEN_3230 = _T_1552 ? _GEN_3222 : _GEN_2086; // @[sequencer-master.scala 168:32]
  wire  _GEN_3231 = _T_1552 ? _GEN_3223 : _GEN_2087; // @[sequencer-master.scala 168:32]
  wire  _GEN_3232 = _T_1552 ? _GEN_3224 : _GEN_2088; // @[sequencer-master.scala 168:32]
  wire  _GEN_3233 = _T_1552 ? _GEN_3225 : _GEN_2089; // @[sequencer-master.scala 168:32]
  wire  _GEN_3234 = _GEN_32729 | _GEN_2106; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3235 = _GEN_32730 | _GEN_2107; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3236 = _GEN_32731 | _GEN_2108; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3237 = _GEN_32732 | _GEN_2109; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3238 = _GEN_32733 | _GEN_2110; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3239 = _GEN_32734 | _GEN_2111; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3240 = _GEN_32735 | _GEN_2112; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3241 = _GEN_32736 | _GEN_2113; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3242 = _T_1574 ? _GEN_3234 : _GEN_2106; // @[sequencer-master.scala 168:32]
  wire  _GEN_3243 = _T_1574 ? _GEN_3235 : _GEN_2107; // @[sequencer-master.scala 168:32]
  wire  _GEN_3244 = _T_1574 ? _GEN_3236 : _GEN_2108; // @[sequencer-master.scala 168:32]
  wire  _GEN_3245 = _T_1574 ? _GEN_3237 : _GEN_2109; // @[sequencer-master.scala 168:32]
  wire  _GEN_3246 = _T_1574 ? _GEN_3238 : _GEN_2110; // @[sequencer-master.scala 168:32]
  wire  _GEN_3247 = _T_1574 ? _GEN_3239 : _GEN_2111; // @[sequencer-master.scala 168:32]
  wire  _GEN_3248 = _T_1574 ? _GEN_3240 : _GEN_2112; // @[sequencer-master.scala 168:32]
  wire  _GEN_3249 = _T_1574 ? _GEN_3241 : _GEN_2113; // @[sequencer-master.scala 168:32]
  wire  _GEN_3250 = _GEN_32729 | _GEN_2130; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3251 = _GEN_32730 | _GEN_2131; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3252 = _GEN_32731 | _GEN_2132; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3253 = _GEN_32732 | _GEN_2133; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3254 = _GEN_32733 | _GEN_2134; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3255 = _GEN_32734 | _GEN_2135; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3256 = _GEN_32735 | _GEN_2136; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3257 = _GEN_32736 | _GEN_2137; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_3258 = _T_1596 ? _GEN_3250 : _GEN_2130; // @[sequencer-master.scala 168:32]
  wire  _GEN_3259 = _T_1596 ? _GEN_3251 : _GEN_2131; // @[sequencer-master.scala 168:32]
  wire  _GEN_3260 = _T_1596 ? _GEN_3252 : _GEN_2132; // @[sequencer-master.scala 168:32]
  wire  _GEN_3261 = _T_1596 ? _GEN_3253 : _GEN_2133; // @[sequencer-master.scala 168:32]
  wire  _GEN_3262 = _T_1596 ? _GEN_3254 : _GEN_2134; // @[sequencer-master.scala 168:32]
  wire  _GEN_3263 = _T_1596 ? _GEN_3255 : _GEN_2135; // @[sequencer-master.scala 168:32]
  wire  _GEN_3264 = _T_1596 ? _GEN_3256 : _GEN_2136; // @[sequencer-master.scala 168:32]
  wire  _GEN_3265 = _T_1596 ? _GEN_3257 : _GEN_2137; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_3266 = 3'h0 == tail ? _T_1615[1:0] : _GEN_1856; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3267 = 3'h1 == tail ? _T_1615[1:0] : _GEN_1857; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3268 = 3'h2 == tail ? _T_1615[1:0] : _GEN_1858; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3269 = 3'h3 == tail ? _T_1615[1:0] : _GEN_1859; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3270 = 3'h4 == tail ? _T_1615[1:0] : _GEN_1860; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3271 = 3'h5 == tail ? _T_1615[1:0] : _GEN_1861; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3272 = 3'h6 == tail ? _T_1615[1:0] : _GEN_1862; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_3273 = 3'h7 == tail ? _T_1615[1:0] : _GEN_1863; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_3274 = 3'h0 == tail ? 4'h0 : _GEN_1864; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3275 = 3'h1 == tail ? 4'h0 : _GEN_1865; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3276 = 3'h2 == tail ? 4'h0 : _GEN_1866; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3277 = 3'h3 == tail ? 4'h0 : _GEN_1867; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3278 = 3'h4 == tail ? 4'h0 : _GEN_1868; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3279 = 3'h5 == tail ? 4'h0 : _GEN_1869; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3280 = 3'h6 == tail ? 4'h0 : _GEN_1870; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_3281 = 3'h7 == tail ? 4'h0 : _GEN_1871; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_3282 = 3'h0 == tail ? 3'h0 : _GEN_1872; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3283 = 3'h1 == tail ? 3'h0 : _GEN_1873; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3284 = 3'h2 == tail ? 3'h0 : _GEN_1874; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3285 = 3'h3 == tail ? 3'h0 : _GEN_1875; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3286 = 3'h4 == tail ? 3'h0 : _GEN_1876; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3287 = 3'h5 == tail ? 3'h0 : _GEN_1877; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3288 = 3'h6 == tail ? 3'h0 : _GEN_1878; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_3289 = 3'h7 == tail ? 3'h0 : _GEN_1879; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [3:0] _T_1837 = _T_1789[3:0] + 4'h1; // @[sequencer-master.scala 247:56]
  wire [3:0] _GEN_3290 = 3'h0 == tail ? _T_1837 : _GEN_3274; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3291 = 3'h1 == tail ? _T_1837 : _GEN_3275; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3292 = 3'h2 == tail ? _T_1837 : _GEN_3276; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3293 = 3'h3 == tail ? _T_1837 : _GEN_3277; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3294 = 3'h4 == tail ? _T_1837 : _GEN_3278; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3295 = 3'h5 == tail ? _T_1837 : _GEN_3279; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3296 = 3'h6 == tail ? _T_1837 : _GEN_3280; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3297 = 3'h7 == tail ? _T_1837 : _GEN_3281; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_3298 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3290 : _GEN_3274; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3299 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3291 : _GEN_3275; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3300 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3292 : _GEN_3276; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3301 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3293 : _GEN_3277; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3302 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3294 : _GEN_3278; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3303 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3295 : _GEN_3279; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3304 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3296 : _GEN_3280; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_3305 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_3297 : _GEN_3281; // @[sequencer-master.scala 235:47]
  wire [2:0] _GEN_3306 = 3'h0 == tail ? _T_1837[2:0] : _GEN_3282; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3307 = 3'h1 == tail ? _T_1837[2:0] : _GEN_3283; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3308 = 3'h2 == tail ? _T_1837[2:0] : _GEN_3284; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3309 = 3'h3 == tail ? _T_1837[2:0] : _GEN_3285; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3310 = 3'h4 == tail ? _T_1837[2:0] : _GEN_3286; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3311 = 3'h5 == tail ? _T_1837[2:0] : _GEN_3287; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3312 = 3'h6 == tail ? _T_1837[2:0] : _GEN_3288; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3313 = 3'h7 == tail ? _T_1837[2:0] : _GEN_3289; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_3314 = io_op_bits_base_vd_pred ? _GEN_3306 : _GEN_3282; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3315 = io_op_bits_base_vd_pred ? _GEN_3307 : _GEN_3283; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3316 = io_op_bits_base_vd_pred ? _GEN_3308 : _GEN_3284; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3317 = io_op_bits_base_vd_pred ? _GEN_3309 : _GEN_3285; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3318 = io_op_bits_base_vd_pred ? _GEN_3310 : _GEN_3286; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3319 = io_op_bits_base_vd_pred ? _GEN_3311 : _GEN_3287; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3320 = io_op_bits_base_vd_pred ? _GEN_3312 : _GEN_3288; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_3321 = io_op_bits_base_vd_pred ? _GEN_3313 : _GEN_3289; // @[sequencer-master.scala 236:45]
  wire  _GEN_3322 = io_op_bits_active_vipred ? _GEN_1882 : _GEN_1400; // @[sequencer-master.scala 641:41]
  wire  _GEN_3323 = io_op_bits_active_vipred ? _GEN_1883 : _GEN_1401; // @[sequencer-master.scala 641:41]
  wire  _GEN_3324 = io_op_bits_active_vipred ? _GEN_1884 : _GEN_1402; // @[sequencer-master.scala 641:41]
  wire  _GEN_3325 = io_op_bits_active_vipred ? _GEN_1885 : _GEN_1403; // @[sequencer-master.scala 641:41]
  wire  _GEN_3326 = io_op_bits_active_vipred ? _GEN_1886 : _GEN_1404; // @[sequencer-master.scala 641:41]
  wire  _GEN_3327 = io_op_bits_active_vipred ? _GEN_1887 : _GEN_1405; // @[sequencer-master.scala 641:41]
  wire  _GEN_3328 = io_op_bits_active_vipred ? _GEN_1888 : _GEN_1406; // @[sequencer-master.scala 641:41]
  wire  _GEN_3329 = io_op_bits_active_vipred ? _GEN_1889 : _GEN_1407; // @[sequencer-master.scala 641:41]
  wire  _GEN_3338 = io_op_bits_active_vipred ? _GEN_1898 : _GEN_1416; // @[sequencer-master.scala 641:41]
  wire  _GEN_3339 = io_op_bits_active_vipred ? _GEN_1899 : _GEN_1417; // @[sequencer-master.scala 641:41]
  wire  _GEN_3340 = io_op_bits_active_vipred ? _GEN_1900 : _GEN_1418; // @[sequencer-master.scala 641:41]
  wire  _GEN_3341 = io_op_bits_active_vipred ? _GEN_1901 : _GEN_1419; // @[sequencer-master.scala 641:41]
  wire  _GEN_3342 = io_op_bits_active_vipred ? _GEN_1902 : _GEN_1420; // @[sequencer-master.scala 641:41]
  wire  _GEN_3343 = io_op_bits_active_vipred ? _GEN_1903 : _GEN_1421; // @[sequencer-master.scala 641:41]
  wire  _GEN_3344 = io_op_bits_active_vipred ? _GEN_1904 : _GEN_1422; // @[sequencer-master.scala 641:41]
  wire  _GEN_3345 = io_op_bits_active_vipred ? _GEN_1905 : _GEN_1423; // @[sequencer-master.scala 641:41]
  wire  _GEN_3346 = io_op_bits_active_vipred ? _GEN_2242 : _GEN_1424; // @[sequencer-master.scala 641:41]
  wire  _GEN_3347 = io_op_bits_active_vipred ? _GEN_2243 : _GEN_1425; // @[sequencer-master.scala 641:41]
  wire  _GEN_3348 = io_op_bits_active_vipred ? _GEN_2244 : _GEN_1426; // @[sequencer-master.scala 641:41]
  wire  _GEN_3349 = io_op_bits_active_vipred ? _GEN_2245 : _GEN_1427; // @[sequencer-master.scala 641:41]
  wire  _GEN_3350 = io_op_bits_active_vipred ? _GEN_2246 : _GEN_1428; // @[sequencer-master.scala 641:41]
  wire  _GEN_3351 = io_op_bits_active_vipred ? _GEN_2247 : _GEN_1429; // @[sequencer-master.scala 641:41]
  wire  _GEN_3352 = io_op_bits_active_vipred ? _GEN_2248 : _GEN_1430; // @[sequencer-master.scala 641:41]
  wire  _GEN_3353 = io_op_bits_active_vipred ? _GEN_2249 : _GEN_1431; // @[sequencer-master.scala 641:41]
  wire  _GEN_3354 = io_op_bits_active_vipred ? _GEN_2490 : _GEN_1432; // @[sequencer-master.scala 641:41]
  wire  _GEN_3355 = io_op_bits_active_vipred ? _GEN_2491 : _GEN_1433; // @[sequencer-master.scala 641:41]
  wire  _GEN_3356 = io_op_bits_active_vipred ? _GEN_2492 : _GEN_1434; // @[sequencer-master.scala 641:41]
  wire  _GEN_3357 = io_op_bits_active_vipred ? _GEN_2493 : _GEN_1435; // @[sequencer-master.scala 641:41]
  wire  _GEN_3358 = io_op_bits_active_vipred ? _GEN_2494 : _GEN_1436; // @[sequencer-master.scala 641:41]
  wire  _GEN_3359 = io_op_bits_active_vipred ? _GEN_2495 : _GEN_1437; // @[sequencer-master.scala 641:41]
  wire  _GEN_3360 = io_op_bits_active_vipred ? _GEN_2496 : _GEN_1438; // @[sequencer-master.scala 641:41]
  wire  _GEN_3361 = io_op_bits_active_vipred ? _GEN_2497 : _GEN_1439; // @[sequencer-master.scala 641:41]
  wire  _GEN_3362 = io_op_bits_active_vipred ? _GEN_2738 : _GEN_1440; // @[sequencer-master.scala 641:41]
  wire  _GEN_3363 = io_op_bits_active_vipred ? _GEN_2739 : _GEN_1441; // @[sequencer-master.scala 641:41]
  wire  _GEN_3364 = io_op_bits_active_vipred ? _GEN_2740 : _GEN_1442; // @[sequencer-master.scala 641:41]
  wire  _GEN_3365 = io_op_bits_active_vipred ? _GEN_2741 : _GEN_1443; // @[sequencer-master.scala 641:41]
  wire  _GEN_3366 = io_op_bits_active_vipred ? _GEN_2742 : _GEN_1444; // @[sequencer-master.scala 641:41]
  wire  _GEN_3367 = io_op_bits_active_vipred ? _GEN_2743 : _GEN_1445; // @[sequencer-master.scala 641:41]
  wire  _GEN_3368 = io_op_bits_active_vipred ? _GEN_2744 : _GEN_1446; // @[sequencer-master.scala 641:41]
  wire  _GEN_3369 = io_op_bits_active_vipred ? _GEN_2745 : _GEN_1447; // @[sequencer-master.scala 641:41]
  wire  _GEN_3370 = io_op_bits_active_vipred ? _GEN_2970 : _GEN_1448; // @[sequencer-master.scala 641:41]
  wire  _GEN_3371 = io_op_bits_active_vipred ? _GEN_2971 : _GEN_1449; // @[sequencer-master.scala 641:41]
  wire  _GEN_3372 = io_op_bits_active_vipred ? _GEN_2972 : _GEN_1450; // @[sequencer-master.scala 641:41]
  wire  _GEN_3373 = io_op_bits_active_vipred ? _GEN_2973 : _GEN_1451; // @[sequencer-master.scala 641:41]
  wire  _GEN_3374 = io_op_bits_active_vipred ? _GEN_2974 : _GEN_1452; // @[sequencer-master.scala 641:41]
  wire  _GEN_3375 = io_op_bits_active_vipred ? _GEN_2975 : _GEN_1453; // @[sequencer-master.scala 641:41]
  wire  _GEN_3376 = io_op_bits_active_vipred ? _GEN_2976 : _GEN_1454; // @[sequencer-master.scala 641:41]
  wire  _GEN_3377 = io_op_bits_active_vipred ? _GEN_2977 : _GEN_1455; // @[sequencer-master.scala 641:41]
  wire  _GEN_3378 = io_op_bits_active_vipred ? _GEN_1938 : _GEN_1456; // @[sequencer-master.scala 641:41]
  wire  _GEN_3379 = io_op_bits_active_vipred ? _GEN_1939 : _GEN_1457; // @[sequencer-master.scala 641:41]
  wire  _GEN_3380 = io_op_bits_active_vipred ? _GEN_1940 : _GEN_1458; // @[sequencer-master.scala 641:41]
  wire  _GEN_3381 = io_op_bits_active_vipred ? _GEN_1941 : _GEN_1459; // @[sequencer-master.scala 641:41]
  wire  _GEN_3382 = io_op_bits_active_vipred ? _GEN_1942 : _GEN_1460; // @[sequencer-master.scala 641:41]
  wire  _GEN_3383 = io_op_bits_active_vipred ? _GEN_1943 : _GEN_1461; // @[sequencer-master.scala 641:41]
  wire  _GEN_3384 = io_op_bits_active_vipred ? _GEN_1944 : _GEN_1462; // @[sequencer-master.scala 641:41]
  wire  _GEN_3385 = io_op_bits_active_vipred ? _GEN_1945 : _GEN_1463; // @[sequencer-master.scala 641:41]
  wire  _GEN_3386 = io_op_bits_active_vipred ? _GEN_2794 : _GEN_1464; // @[sequencer-master.scala 641:41]
  wire  _GEN_3387 = io_op_bits_active_vipred ? _GEN_2795 : _GEN_1465; // @[sequencer-master.scala 641:41]
  wire  _GEN_3388 = io_op_bits_active_vipred ? _GEN_2796 : _GEN_1466; // @[sequencer-master.scala 641:41]
  wire  _GEN_3389 = io_op_bits_active_vipred ? _GEN_2797 : _GEN_1467; // @[sequencer-master.scala 641:41]
  wire  _GEN_3390 = io_op_bits_active_vipred ? _GEN_2798 : _GEN_1468; // @[sequencer-master.scala 641:41]
  wire  _GEN_3391 = io_op_bits_active_vipred ? _GEN_2799 : _GEN_1469; // @[sequencer-master.scala 641:41]
  wire  _GEN_3392 = io_op_bits_active_vipred ? _GEN_2800 : _GEN_1470; // @[sequencer-master.scala 641:41]
  wire  _GEN_3393 = io_op_bits_active_vipred ? _GEN_2801 : _GEN_1471; // @[sequencer-master.scala 641:41]
  wire  _GEN_3394 = io_op_bits_active_vipred ? _GEN_3018 : _GEN_1472; // @[sequencer-master.scala 641:41]
  wire  _GEN_3395 = io_op_bits_active_vipred ? _GEN_3019 : _GEN_1473; // @[sequencer-master.scala 641:41]
  wire  _GEN_3396 = io_op_bits_active_vipred ? _GEN_3020 : _GEN_1474; // @[sequencer-master.scala 641:41]
  wire  _GEN_3397 = io_op_bits_active_vipred ? _GEN_3021 : _GEN_1475; // @[sequencer-master.scala 641:41]
  wire  _GEN_3398 = io_op_bits_active_vipred ? _GEN_3022 : _GEN_1476; // @[sequencer-master.scala 641:41]
  wire  _GEN_3399 = io_op_bits_active_vipred ? _GEN_3023 : _GEN_1477; // @[sequencer-master.scala 641:41]
  wire  _GEN_3400 = io_op_bits_active_vipred ? _GEN_3024 : _GEN_1478; // @[sequencer-master.scala 641:41]
  wire  _GEN_3401 = io_op_bits_active_vipred ? _GEN_3025 : _GEN_1479; // @[sequencer-master.scala 641:41]
  wire  _GEN_3402 = io_op_bits_active_vipred ? _GEN_3146 : _GEN_1480; // @[sequencer-master.scala 641:41]
  wire  _GEN_3403 = io_op_bits_active_vipred ? _GEN_3147 : _GEN_1481; // @[sequencer-master.scala 641:41]
  wire  _GEN_3404 = io_op_bits_active_vipred ? _GEN_3148 : _GEN_1482; // @[sequencer-master.scala 641:41]
  wire  _GEN_3405 = io_op_bits_active_vipred ? _GEN_3149 : _GEN_1483; // @[sequencer-master.scala 641:41]
  wire  _GEN_3406 = io_op_bits_active_vipred ? _GEN_3150 : _GEN_1484; // @[sequencer-master.scala 641:41]
  wire  _GEN_3407 = io_op_bits_active_vipred ? _GEN_3151 : _GEN_1485; // @[sequencer-master.scala 641:41]
  wire  _GEN_3408 = io_op_bits_active_vipred ? _GEN_3152 : _GEN_1486; // @[sequencer-master.scala 641:41]
  wire  _GEN_3409 = io_op_bits_active_vipred ? _GEN_3153 : _GEN_1487; // @[sequencer-master.scala 641:41]
  wire  _GEN_3410 = io_op_bits_active_vipred ? _GEN_2810 : _GEN_1488; // @[sequencer-master.scala 641:41]
  wire  _GEN_3411 = io_op_bits_active_vipred ? _GEN_2811 : _GEN_1489; // @[sequencer-master.scala 641:41]
  wire  _GEN_3412 = io_op_bits_active_vipred ? _GEN_2812 : _GEN_1490; // @[sequencer-master.scala 641:41]
  wire  _GEN_3413 = io_op_bits_active_vipred ? _GEN_2813 : _GEN_1491; // @[sequencer-master.scala 641:41]
  wire  _GEN_3414 = io_op_bits_active_vipred ? _GEN_2814 : _GEN_1492; // @[sequencer-master.scala 641:41]
  wire  _GEN_3415 = io_op_bits_active_vipred ? _GEN_2815 : _GEN_1493; // @[sequencer-master.scala 641:41]
  wire  _GEN_3416 = io_op_bits_active_vipred ? _GEN_2816 : _GEN_1494; // @[sequencer-master.scala 641:41]
  wire  _GEN_3417 = io_op_bits_active_vipred ? _GEN_2817 : _GEN_1495; // @[sequencer-master.scala 641:41]
  wire  _GEN_3418 = io_op_bits_active_vipred ? _GEN_3034 : _GEN_1496; // @[sequencer-master.scala 641:41]
  wire  _GEN_3419 = io_op_bits_active_vipred ? _GEN_3035 : _GEN_1497; // @[sequencer-master.scala 641:41]
  wire  _GEN_3420 = io_op_bits_active_vipred ? _GEN_3036 : _GEN_1498; // @[sequencer-master.scala 641:41]
  wire  _GEN_3421 = io_op_bits_active_vipred ? _GEN_3037 : _GEN_1499; // @[sequencer-master.scala 641:41]
  wire  _GEN_3422 = io_op_bits_active_vipred ? _GEN_3038 : _GEN_1500; // @[sequencer-master.scala 641:41]
  wire  _GEN_3423 = io_op_bits_active_vipred ? _GEN_3039 : _GEN_1501; // @[sequencer-master.scala 641:41]
  wire  _GEN_3424 = io_op_bits_active_vipred ? _GEN_3040 : _GEN_1502; // @[sequencer-master.scala 641:41]
  wire  _GEN_3425 = io_op_bits_active_vipred ? _GEN_3041 : _GEN_1503; // @[sequencer-master.scala 641:41]
  wire  _GEN_3426 = io_op_bits_active_vipred ? _GEN_3162 : _GEN_1504; // @[sequencer-master.scala 641:41]
  wire  _GEN_3427 = io_op_bits_active_vipred ? _GEN_3163 : _GEN_1505; // @[sequencer-master.scala 641:41]
  wire  _GEN_3428 = io_op_bits_active_vipred ? _GEN_3164 : _GEN_1506; // @[sequencer-master.scala 641:41]
  wire  _GEN_3429 = io_op_bits_active_vipred ? _GEN_3165 : _GEN_1507; // @[sequencer-master.scala 641:41]
  wire  _GEN_3430 = io_op_bits_active_vipred ? _GEN_3166 : _GEN_1508; // @[sequencer-master.scala 641:41]
  wire  _GEN_3431 = io_op_bits_active_vipred ? _GEN_3167 : _GEN_1509; // @[sequencer-master.scala 641:41]
  wire  _GEN_3432 = io_op_bits_active_vipred ? _GEN_3168 : _GEN_1510; // @[sequencer-master.scala 641:41]
  wire  _GEN_3433 = io_op_bits_active_vipred ? _GEN_3169 : _GEN_1511; // @[sequencer-master.scala 641:41]
  wire  _GEN_3434 = io_op_bits_active_vipred ? _GEN_2826 : _GEN_1512; // @[sequencer-master.scala 641:41]
  wire  _GEN_3435 = io_op_bits_active_vipred ? _GEN_2827 : _GEN_1513; // @[sequencer-master.scala 641:41]
  wire  _GEN_3436 = io_op_bits_active_vipred ? _GEN_2828 : _GEN_1514; // @[sequencer-master.scala 641:41]
  wire  _GEN_3437 = io_op_bits_active_vipred ? _GEN_2829 : _GEN_1515; // @[sequencer-master.scala 641:41]
  wire  _GEN_3438 = io_op_bits_active_vipred ? _GEN_2830 : _GEN_1516; // @[sequencer-master.scala 641:41]
  wire  _GEN_3439 = io_op_bits_active_vipred ? _GEN_2831 : _GEN_1517; // @[sequencer-master.scala 641:41]
  wire  _GEN_3440 = io_op_bits_active_vipred ? _GEN_2832 : _GEN_1518; // @[sequencer-master.scala 641:41]
  wire  _GEN_3441 = io_op_bits_active_vipred ? _GEN_2833 : _GEN_1519; // @[sequencer-master.scala 641:41]
  wire  _GEN_3442 = io_op_bits_active_vipred ? _GEN_3050 : _GEN_1520; // @[sequencer-master.scala 641:41]
  wire  _GEN_3443 = io_op_bits_active_vipred ? _GEN_3051 : _GEN_1521; // @[sequencer-master.scala 641:41]
  wire  _GEN_3444 = io_op_bits_active_vipred ? _GEN_3052 : _GEN_1522; // @[sequencer-master.scala 641:41]
  wire  _GEN_3445 = io_op_bits_active_vipred ? _GEN_3053 : _GEN_1523; // @[sequencer-master.scala 641:41]
  wire  _GEN_3446 = io_op_bits_active_vipred ? _GEN_3054 : _GEN_1524; // @[sequencer-master.scala 641:41]
  wire  _GEN_3447 = io_op_bits_active_vipred ? _GEN_3055 : _GEN_1525; // @[sequencer-master.scala 641:41]
  wire  _GEN_3448 = io_op_bits_active_vipred ? _GEN_3056 : _GEN_1526; // @[sequencer-master.scala 641:41]
  wire  _GEN_3449 = io_op_bits_active_vipred ? _GEN_3057 : _GEN_1527; // @[sequencer-master.scala 641:41]
  wire  _GEN_3450 = io_op_bits_active_vipred ? _GEN_3178 : _GEN_1528; // @[sequencer-master.scala 641:41]
  wire  _GEN_3451 = io_op_bits_active_vipred ? _GEN_3179 : _GEN_1529; // @[sequencer-master.scala 641:41]
  wire  _GEN_3452 = io_op_bits_active_vipred ? _GEN_3180 : _GEN_1530; // @[sequencer-master.scala 641:41]
  wire  _GEN_3453 = io_op_bits_active_vipred ? _GEN_3181 : _GEN_1531; // @[sequencer-master.scala 641:41]
  wire  _GEN_3454 = io_op_bits_active_vipred ? _GEN_3182 : _GEN_1532; // @[sequencer-master.scala 641:41]
  wire  _GEN_3455 = io_op_bits_active_vipred ? _GEN_3183 : _GEN_1533; // @[sequencer-master.scala 641:41]
  wire  _GEN_3456 = io_op_bits_active_vipred ? _GEN_3184 : _GEN_1534; // @[sequencer-master.scala 641:41]
  wire  _GEN_3457 = io_op_bits_active_vipred ? _GEN_3185 : _GEN_1535; // @[sequencer-master.scala 641:41]
  wire  _GEN_3458 = io_op_bits_active_vipred ? _GEN_2842 : _GEN_1536; // @[sequencer-master.scala 641:41]
  wire  _GEN_3459 = io_op_bits_active_vipred ? _GEN_2843 : _GEN_1537; // @[sequencer-master.scala 641:41]
  wire  _GEN_3460 = io_op_bits_active_vipred ? _GEN_2844 : _GEN_1538; // @[sequencer-master.scala 641:41]
  wire  _GEN_3461 = io_op_bits_active_vipred ? _GEN_2845 : _GEN_1539; // @[sequencer-master.scala 641:41]
  wire  _GEN_3462 = io_op_bits_active_vipred ? _GEN_2846 : _GEN_1540; // @[sequencer-master.scala 641:41]
  wire  _GEN_3463 = io_op_bits_active_vipred ? _GEN_2847 : _GEN_1541; // @[sequencer-master.scala 641:41]
  wire  _GEN_3464 = io_op_bits_active_vipred ? _GEN_2848 : _GEN_1542; // @[sequencer-master.scala 641:41]
  wire  _GEN_3465 = io_op_bits_active_vipred ? _GEN_2849 : _GEN_1543; // @[sequencer-master.scala 641:41]
  wire  _GEN_3466 = io_op_bits_active_vipred ? _GEN_3066 : _GEN_1544; // @[sequencer-master.scala 641:41]
  wire  _GEN_3467 = io_op_bits_active_vipred ? _GEN_3067 : _GEN_1545; // @[sequencer-master.scala 641:41]
  wire  _GEN_3468 = io_op_bits_active_vipred ? _GEN_3068 : _GEN_1546; // @[sequencer-master.scala 641:41]
  wire  _GEN_3469 = io_op_bits_active_vipred ? _GEN_3069 : _GEN_1547; // @[sequencer-master.scala 641:41]
  wire  _GEN_3470 = io_op_bits_active_vipred ? _GEN_3070 : _GEN_1548; // @[sequencer-master.scala 641:41]
  wire  _GEN_3471 = io_op_bits_active_vipred ? _GEN_3071 : _GEN_1549; // @[sequencer-master.scala 641:41]
  wire  _GEN_3472 = io_op_bits_active_vipred ? _GEN_3072 : _GEN_1550; // @[sequencer-master.scala 641:41]
  wire  _GEN_3473 = io_op_bits_active_vipred ? _GEN_3073 : _GEN_1551; // @[sequencer-master.scala 641:41]
  wire  _GEN_3474 = io_op_bits_active_vipred ? _GEN_3194 : _GEN_1552; // @[sequencer-master.scala 641:41]
  wire  _GEN_3475 = io_op_bits_active_vipred ? _GEN_3195 : _GEN_1553; // @[sequencer-master.scala 641:41]
  wire  _GEN_3476 = io_op_bits_active_vipred ? _GEN_3196 : _GEN_1554; // @[sequencer-master.scala 641:41]
  wire  _GEN_3477 = io_op_bits_active_vipred ? _GEN_3197 : _GEN_1555; // @[sequencer-master.scala 641:41]
  wire  _GEN_3478 = io_op_bits_active_vipred ? _GEN_3198 : _GEN_1556; // @[sequencer-master.scala 641:41]
  wire  _GEN_3479 = io_op_bits_active_vipred ? _GEN_3199 : _GEN_1557; // @[sequencer-master.scala 641:41]
  wire  _GEN_3480 = io_op_bits_active_vipred ? _GEN_3200 : _GEN_1558; // @[sequencer-master.scala 641:41]
  wire  _GEN_3481 = io_op_bits_active_vipred ? _GEN_3201 : _GEN_1559; // @[sequencer-master.scala 641:41]
  wire  _GEN_3482 = io_op_bits_active_vipred ? _GEN_2858 : _GEN_1560; // @[sequencer-master.scala 641:41]
  wire  _GEN_3483 = io_op_bits_active_vipred ? _GEN_2859 : _GEN_1561; // @[sequencer-master.scala 641:41]
  wire  _GEN_3484 = io_op_bits_active_vipred ? _GEN_2860 : _GEN_1562; // @[sequencer-master.scala 641:41]
  wire  _GEN_3485 = io_op_bits_active_vipred ? _GEN_2861 : _GEN_1563; // @[sequencer-master.scala 641:41]
  wire  _GEN_3486 = io_op_bits_active_vipred ? _GEN_2862 : _GEN_1564; // @[sequencer-master.scala 641:41]
  wire  _GEN_3487 = io_op_bits_active_vipred ? _GEN_2863 : _GEN_1565; // @[sequencer-master.scala 641:41]
  wire  _GEN_3488 = io_op_bits_active_vipred ? _GEN_2864 : _GEN_1566; // @[sequencer-master.scala 641:41]
  wire  _GEN_3489 = io_op_bits_active_vipred ? _GEN_2865 : _GEN_1567; // @[sequencer-master.scala 641:41]
  wire  _GEN_3490 = io_op_bits_active_vipred ? _GEN_3082 : _GEN_1568; // @[sequencer-master.scala 641:41]
  wire  _GEN_3491 = io_op_bits_active_vipred ? _GEN_3083 : _GEN_1569; // @[sequencer-master.scala 641:41]
  wire  _GEN_3492 = io_op_bits_active_vipred ? _GEN_3084 : _GEN_1570; // @[sequencer-master.scala 641:41]
  wire  _GEN_3493 = io_op_bits_active_vipred ? _GEN_3085 : _GEN_1571; // @[sequencer-master.scala 641:41]
  wire  _GEN_3494 = io_op_bits_active_vipred ? _GEN_3086 : _GEN_1572; // @[sequencer-master.scala 641:41]
  wire  _GEN_3495 = io_op_bits_active_vipred ? _GEN_3087 : _GEN_1573; // @[sequencer-master.scala 641:41]
  wire  _GEN_3496 = io_op_bits_active_vipred ? _GEN_3088 : _GEN_1574; // @[sequencer-master.scala 641:41]
  wire  _GEN_3497 = io_op_bits_active_vipred ? _GEN_3089 : _GEN_1575; // @[sequencer-master.scala 641:41]
  wire  _GEN_3498 = io_op_bits_active_vipred ? _GEN_3210 : _GEN_1576; // @[sequencer-master.scala 641:41]
  wire  _GEN_3499 = io_op_bits_active_vipred ? _GEN_3211 : _GEN_1577; // @[sequencer-master.scala 641:41]
  wire  _GEN_3500 = io_op_bits_active_vipred ? _GEN_3212 : _GEN_1578; // @[sequencer-master.scala 641:41]
  wire  _GEN_3501 = io_op_bits_active_vipred ? _GEN_3213 : _GEN_1579; // @[sequencer-master.scala 641:41]
  wire  _GEN_3502 = io_op_bits_active_vipred ? _GEN_3214 : _GEN_1580; // @[sequencer-master.scala 641:41]
  wire  _GEN_3503 = io_op_bits_active_vipred ? _GEN_3215 : _GEN_1581; // @[sequencer-master.scala 641:41]
  wire  _GEN_3504 = io_op_bits_active_vipred ? _GEN_3216 : _GEN_1582; // @[sequencer-master.scala 641:41]
  wire  _GEN_3505 = io_op_bits_active_vipred ? _GEN_3217 : _GEN_1583; // @[sequencer-master.scala 641:41]
  wire  _GEN_3506 = io_op_bits_active_vipred ? _GEN_2874 : _GEN_1584; // @[sequencer-master.scala 641:41]
  wire  _GEN_3507 = io_op_bits_active_vipred ? _GEN_2875 : _GEN_1585; // @[sequencer-master.scala 641:41]
  wire  _GEN_3508 = io_op_bits_active_vipred ? _GEN_2876 : _GEN_1586; // @[sequencer-master.scala 641:41]
  wire  _GEN_3509 = io_op_bits_active_vipred ? _GEN_2877 : _GEN_1587; // @[sequencer-master.scala 641:41]
  wire  _GEN_3510 = io_op_bits_active_vipred ? _GEN_2878 : _GEN_1588; // @[sequencer-master.scala 641:41]
  wire  _GEN_3511 = io_op_bits_active_vipred ? _GEN_2879 : _GEN_1589; // @[sequencer-master.scala 641:41]
  wire  _GEN_3512 = io_op_bits_active_vipred ? _GEN_2880 : _GEN_1590; // @[sequencer-master.scala 641:41]
  wire  _GEN_3513 = io_op_bits_active_vipred ? _GEN_2881 : _GEN_1591; // @[sequencer-master.scala 641:41]
  wire  _GEN_3514 = io_op_bits_active_vipred ? _GEN_3098 : _GEN_1592; // @[sequencer-master.scala 641:41]
  wire  _GEN_3515 = io_op_bits_active_vipred ? _GEN_3099 : _GEN_1593; // @[sequencer-master.scala 641:41]
  wire  _GEN_3516 = io_op_bits_active_vipred ? _GEN_3100 : _GEN_1594; // @[sequencer-master.scala 641:41]
  wire  _GEN_3517 = io_op_bits_active_vipred ? _GEN_3101 : _GEN_1595; // @[sequencer-master.scala 641:41]
  wire  _GEN_3518 = io_op_bits_active_vipred ? _GEN_3102 : _GEN_1596; // @[sequencer-master.scala 641:41]
  wire  _GEN_3519 = io_op_bits_active_vipred ? _GEN_3103 : _GEN_1597; // @[sequencer-master.scala 641:41]
  wire  _GEN_3520 = io_op_bits_active_vipred ? _GEN_3104 : _GEN_1598; // @[sequencer-master.scala 641:41]
  wire  _GEN_3521 = io_op_bits_active_vipred ? _GEN_3105 : _GEN_1599; // @[sequencer-master.scala 641:41]
  wire  _GEN_3522 = io_op_bits_active_vipred ? _GEN_3226 : _GEN_1600; // @[sequencer-master.scala 641:41]
  wire  _GEN_3523 = io_op_bits_active_vipred ? _GEN_3227 : _GEN_1601; // @[sequencer-master.scala 641:41]
  wire  _GEN_3524 = io_op_bits_active_vipred ? _GEN_3228 : _GEN_1602; // @[sequencer-master.scala 641:41]
  wire  _GEN_3525 = io_op_bits_active_vipred ? _GEN_3229 : _GEN_1603; // @[sequencer-master.scala 641:41]
  wire  _GEN_3526 = io_op_bits_active_vipred ? _GEN_3230 : _GEN_1604; // @[sequencer-master.scala 641:41]
  wire  _GEN_3527 = io_op_bits_active_vipred ? _GEN_3231 : _GEN_1605; // @[sequencer-master.scala 641:41]
  wire  _GEN_3528 = io_op_bits_active_vipred ? _GEN_3232 : _GEN_1606; // @[sequencer-master.scala 641:41]
  wire  _GEN_3529 = io_op_bits_active_vipred ? _GEN_3233 : _GEN_1607; // @[sequencer-master.scala 641:41]
  wire  _GEN_3530 = io_op_bits_active_vipred ? _GEN_2890 : _GEN_1608; // @[sequencer-master.scala 641:41]
  wire  _GEN_3531 = io_op_bits_active_vipred ? _GEN_2891 : _GEN_1609; // @[sequencer-master.scala 641:41]
  wire  _GEN_3532 = io_op_bits_active_vipred ? _GEN_2892 : _GEN_1610; // @[sequencer-master.scala 641:41]
  wire  _GEN_3533 = io_op_bits_active_vipred ? _GEN_2893 : _GEN_1611; // @[sequencer-master.scala 641:41]
  wire  _GEN_3534 = io_op_bits_active_vipred ? _GEN_2894 : _GEN_1612; // @[sequencer-master.scala 641:41]
  wire  _GEN_3535 = io_op_bits_active_vipred ? _GEN_2895 : _GEN_1613; // @[sequencer-master.scala 641:41]
  wire  _GEN_3536 = io_op_bits_active_vipred ? _GEN_2896 : _GEN_1614; // @[sequencer-master.scala 641:41]
  wire  _GEN_3537 = io_op_bits_active_vipred ? _GEN_2897 : _GEN_1615; // @[sequencer-master.scala 641:41]
  wire  _GEN_3538 = io_op_bits_active_vipred ? _GEN_3114 : _GEN_1616; // @[sequencer-master.scala 641:41]
  wire  _GEN_3539 = io_op_bits_active_vipred ? _GEN_3115 : _GEN_1617; // @[sequencer-master.scala 641:41]
  wire  _GEN_3540 = io_op_bits_active_vipred ? _GEN_3116 : _GEN_1618; // @[sequencer-master.scala 641:41]
  wire  _GEN_3541 = io_op_bits_active_vipred ? _GEN_3117 : _GEN_1619; // @[sequencer-master.scala 641:41]
  wire  _GEN_3542 = io_op_bits_active_vipred ? _GEN_3118 : _GEN_1620; // @[sequencer-master.scala 641:41]
  wire  _GEN_3543 = io_op_bits_active_vipred ? _GEN_3119 : _GEN_1621; // @[sequencer-master.scala 641:41]
  wire  _GEN_3544 = io_op_bits_active_vipred ? _GEN_3120 : _GEN_1622; // @[sequencer-master.scala 641:41]
  wire  _GEN_3545 = io_op_bits_active_vipred ? _GEN_3121 : _GEN_1623; // @[sequencer-master.scala 641:41]
  wire  _GEN_3546 = io_op_bits_active_vipred ? _GEN_3242 : _GEN_1624; // @[sequencer-master.scala 641:41]
  wire  _GEN_3547 = io_op_bits_active_vipred ? _GEN_3243 : _GEN_1625; // @[sequencer-master.scala 641:41]
  wire  _GEN_3548 = io_op_bits_active_vipred ? _GEN_3244 : _GEN_1626; // @[sequencer-master.scala 641:41]
  wire  _GEN_3549 = io_op_bits_active_vipred ? _GEN_3245 : _GEN_1627; // @[sequencer-master.scala 641:41]
  wire  _GEN_3550 = io_op_bits_active_vipred ? _GEN_3246 : _GEN_1628; // @[sequencer-master.scala 641:41]
  wire  _GEN_3551 = io_op_bits_active_vipred ? _GEN_3247 : _GEN_1629; // @[sequencer-master.scala 641:41]
  wire  _GEN_3552 = io_op_bits_active_vipred ? _GEN_3248 : _GEN_1630; // @[sequencer-master.scala 641:41]
  wire  _GEN_3553 = io_op_bits_active_vipred ? _GEN_3249 : _GEN_1631; // @[sequencer-master.scala 641:41]
  wire  _GEN_3554 = io_op_bits_active_vipred ? _GEN_2906 : _GEN_1632; // @[sequencer-master.scala 641:41]
  wire  _GEN_3555 = io_op_bits_active_vipred ? _GEN_2907 : _GEN_1633; // @[sequencer-master.scala 641:41]
  wire  _GEN_3556 = io_op_bits_active_vipred ? _GEN_2908 : _GEN_1634; // @[sequencer-master.scala 641:41]
  wire  _GEN_3557 = io_op_bits_active_vipred ? _GEN_2909 : _GEN_1635; // @[sequencer-master.scala 641:41]
  wire  _GEN_3558 = io_op_bits_active_vipred ? _GEN_2910 : _GEN_1636; // @[sequencer-master.scala 641:41]
  wire  _GEN_3559 = io_op_bits_active_vipred ? _GEN_2911 : _GEN_1637; // @[sequencer-master.scala 641:41]
  wire  _GEN_3560 = io_op_bits_active_vipred ? _GEN_2912 : _GEN_1638; // @[sequencer-master.scala 641:41]
  wire  _GEN_3561 = io_op_bits_active_vipred ? _GEN_2913 : _GEN_1639; // @[sequencer-master.scala 641:41]
  wire  _GEN_3562 = io_op_bits_active_vipred ? _GEN_3130 : _GEN_1640; // @[sequencer-master.scala 641:41]
  wire  _GEN_3563 = io_op_bits_active_vipred ? _GEN_3131 : _GEN_1641; // @[sequencer-master.scala 641:41]
  wire  _GEN_3564 = io_op_bits_active_vipred ? _GEN_3132 : _GEN_1642; // @[sequencer-master.scala 641:41]
  wire  _GEN_3565 = io_op_bits_active_vipred ? _GEN_3133 : _GEN_1643; // @[sequencer-master.scala 641:41]
  wire  _GEN_3566 = io_op_bits_active_vipred ? _GEN_3134 : _GEN_1644; // @[sequencer-master.scala 641:41]
  wire  _GEN_3567 = io_op_bits_active_vipred ? _GEN_3135 : _GEN_1645; // @[sequencer-master.scala 641:41]
  wire  _GEN_3568 = io_op_bits_active_vipred ? _GEN_3136 : _GEN_1646; // @[sequencer-master.scala 641:41]
  wire  _GEN_3569 = io_op_bits_active_vipred ? _GEN_3137 : _GEN_1647; // @[sequencer-master.scala 641:41]
  wire  _GEN_3570 = io_op_bits_active_vipred ? _GEN_3258 : _GEN_1648; // @[sequencer-master.scala 641:41]
  wire  _GEN_3571 = io_op_bits_active_vipred ? _GEN_3259 : _GEN_1649; // @[sequencer-master.scala 641:41]
  wire  _GEN_3572 = io_op_bits_active_vipred ? _GEN_3260 : _GEN_1650; // @[sequencer-master.scala 641:41]
  wire  _GEN_3573 = io_op_bits_active_vipred ? _GEN_3261 : _GEN_1651; // @[sequencer-master.scala 641:41]
  wire  _GEN_3574 = io_op_bits_active_vipred ? _GEN_3262 : _GEN_1652; // @[sequencer-master.scala 641:41]
  wire  _GEN_3575 = io_op_bits_active_vipred ? _GEN_3263 : _GEN_1653; // @[sequencer-master.scala 641:41]
  wire  _GEN_3576 = io_op_bits_active_vipred ? _GEN_3264 : _GEN_1654; // @[sequencer-master.scala 641:41]
  wire  _GEN_3577 = io_op_bits_active_vipred ? _GEN_3265 : _GEN_1655; // @[sequencer-master.scala 641:41]
  wire  _GEN_3578 = io_op_bits_active_vipred ? _GEN_2138 : _GEN_1656; // @[sequencer-master.scala 641:41]
  wire  _GEN_3579 = io_op_bits_active_vipred ? _GEN_2139 : _GEN_1657; // @[sequencer-master.scala 641:41]
  wire  _GEN_3580 = io_op_bits_active_vipred ? _GEN_2140 : _GEN_1658; // @[sequencer-master.scala 641:41]
  wire  _GEN_3581 = io_op_bits_active_vipred ? _GEN_2141 : _GEN_1659; // @[sequencer-master.scala 641:41]
  wire  _GEN_3582 = io_op_bits_active_vipred ? _GEN_2142 : _GEN_1660; // @[sequencer-master.scala 641:41]
  wire  _GEN_3583 = io_op_bits_active_vipred ? _GEN_2143 : _GEN_1661; // @[sequencer-master.scala 641:41]
  wire  _GEN_3584 = io_op_bits_active_vipred ? _GEN_2144 : _GEN_1662; // @[sequencer-master.scala 641:41]
  wire  _GEN_3585 = io_op_bits_active_vipred ? _GEN_2145 : _GEN_1663; // @[sequencer-master.scala 641:41]
  wire  _GEN_3594 = io_op_bits_active_vipred ? _GEN_2154 : e_0_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3595 = io_op_bits_active_vipred ? _GEN_2155 : e_1_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3596 = io_op_bits_active_vipred ? _GEN_2156 : e_2_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3597 = io_op_bits_active_vipred ? _GEN_2157 : e_3_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3598 = io_op_bits_active_vipred ? _GEN_2158 : e_4_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3599 = io_op_bits_active_vipred ? _GEN_2159 : e_5_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3600 = io_op_bits_active_vipred ? _GEN_2160 : e_6_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3601 = io_op_bits_active_vipred ? _GEN_2161 : e_7_active_vipu; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [9:0] _GEN_3602 = io_op_bits_active_vipred ? _GEN_2162 : _GEN_1680; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3603 = io_op_bits_active_vipred ? _GEN_2163 : _GEN_1681; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3604 = io_op_bits_active_vipred ? _GEN_2164 : _GEN_1682; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3605 = io_op_bits_active_vipred ? _GEN_2165 : _GEN_1683; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3606 = io_op_bits_active_vipred ? _GEN_2166 : _GEN_1684; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3607 = io_op_bits_active_vipred ? _GEN_2167 : _GEN_1685; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3608 = io_op_bits_active_vipred ? _GEN_2168 : _GEN_1686; // @[sequencer-master.scala 641:41]
  wire [9:0] _GEN_3609 = io_op_bits_active_vipred ? _GEN_2169 : _GEN_1687; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3610 = io_op_bits_active_vipred ? _GEN_2234 : _GEN_1720; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3611 = io_op_bits_active_vipred ? _GEN_2235 : _GEN_1721; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3612 = io_op_bits_active_vipred ? _GEN_2236 : _GEN_1722; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3613 = io_op_bits_active_vipred ? _GEN_2237 : _GEN_1723; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3614 = io_op_bits_active_vipred ? _GEN_2238 : _GEN_1724; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3615 = io_op_bits_active_vipred ? _GEN_2239 : _GEN_1725; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3616 = io_op_bits_active_vipred ? _GEN_2240 : _GEN_1726; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3617 = io_op_bits_active_vipred ? _GEN_2241 : _GEN_1727; // @[sequencer-master.scala 641:41]
  wire  _GEN_3618 = io_op_bits_active_vipred ? _GEN_2250 : _GEN_1728; // @[sequencer-master.scala 641:41]
  wire  _GEN_3619 = io_op_bits_active_vipred ? _GEN_2251 : _GEN_1729; // @[sequencer-master.scala 641:41]
  wire  _GEN_3620 = io_op_bits_active_vipred ? _GEN_2252 : _GEN_1730; // @[sequencer-master.scala 641:41]
  wire  _GEN_3621 = io_op_bits_active_vipred ? _GEN_2253 : _GEN_1731; // @[sequencer-master.scala 641:41]
  wire  _GEN_3622 = io_op_bits_active_vipred ? _GEN_2254 : _GEN_1732; // @[sequencer-master.scala 641:41]
  wire  _GEN_3623 = io_op_bits_active_vipred ? _GEN_2255 : _GEN_1733; // @[sequencer-master.scala 641:41]
  wire  _GEN_3624 = io_op_bits_active_vipred ? _GEN_2256 : _GEN_1734; // @[sequencer-master.scala 641:41]
  wire  _GEN_3625 = io_op_bits_active_vipred ? _GEN_2257 : _GEN_1735; // @[sequencer-master.scala 641:41]
  wire  _GEN_3626 = io_op_bits_active_vipred ? _GEN_2258 : _GEN_1736; // @[sequencer-master.scala 641:41]
  wire  _GEN_3627 = io_op_bits_active_vipred ? _GEN_2259 : _GEN_1737; // @[sequencer-master.scala 641:41]
  wire  _GEN_3628 = io_op_bits_active_vipred ? _GEN_2260 : _GEN_1738; // @[sequencer-master.scala 641:41]
  wire  _GEN_3629 = io_op_bits_active_vipred ? _GEN_2261 : _GEN_1739; // @[sequencer-master.scala 641:41]
  wire  _GEN_3630 = io_op_bits_active_vipred ? _GEN_2262 : _GEN_1740; // @[sequencer-master.scala 641:41]
  wire  _GEN_3631 = io_op_bits_active_vipred ? _GEN_2263 : _GEN_1741; // @[sequencer-master.scala 641:41]
  wire  _GEN_3632 = io_op_bits_active_vipred ? _GEN_2264 : _GEN_1742; // @[sequencer-master.scala 641:41]
  wire  _GEN_3633 = io_op_bits_active_vipred ? _GEN_2265 : _GEN_1743; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3634 = io_op_bits_active_vipred ? _GEN_2266 : _GEN_1744; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3635 = io_op_bits_active_vipred ? _GEN_2267 : _GEN_1745; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3636 = io_op_bits_active_vipred ? _GEN_2268 : _GEN_1746; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3637 = io_op_bits_active_vipred ? _GEN_2269 : _GEN_1747; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3638 = io_op_bits_active_vipred ? _GEN_2270 : _GEN_1748; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3639 = io_op_bits_active_vipred ? _GEN_2271 : _GEN_1749; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3640 = io_op_bits_active_vipred ? _GEN_2272 : _GEN_1750; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3641 = io_op_bits_active_vipred ? _GEN_2273 : _GEN_1751; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3642 = io_op_bits_active_vipred ? _GEN_2274 : _GEN_1752; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3643 = io_op_bits_active_vipred ? _GEN_2275 : _GEN_1753; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3644 = io_op_bits_active_vipred ? _GEN_2276 : _GEN_1754; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3645 = io_op_bits_active_vipred ? _GEN_2277 : _GEN_1755; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3646 = io_op_bits_active_vipred ? _GEN_2278 : _GEN_1756; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3647 = io_op_bits_active_vipred ? _GEN_2279 : _GEN_1757; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3648 = io_op_bits_active_vipred ? _GEN_2280 : _GEN_1758; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3649 = io_op_bits_active_vipred ? _GEN_2281 : _GEN_1759; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3650 = io_op_bits_active_vipred ? _GEN_2282 : _GEN_1760; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3651 = io_op_bits_active_vipred ? _GEN_2283 : _GEN_1761; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3652 = io_op_bits_active_vipred ? _GEN_2284 : _GEN_1762; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3653 = io_op_bits_active_vipred ? _GEN_2285 : _GEN_1763; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3654 = io_op_bits_active_vipred ? _GEN_2286 : _GEN_1764; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3655 = io_op_bits_active_vipred ? _GEN_2287 : _GEN_1765; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3656 = io_op_bits_active_vipred ? _GEN_2288 : _GEN_1766; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3657 = io_op_bits_active_vipred ? _GEN_2289 : _GEN_1767; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3658 = io_op_bits_active_vipred ? _GEN_2482 : _GEN_1768; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3659 = io_op_bits_active_vipred ? _GEN_2483 : _GEN_1769; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3660 = io_op_bits_active_vipred ? _GEN_2484 : _GEN_1770; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3661 = io_op_bits_active_vipred ? _GEN_2485 : _GEN_1771; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3662 = io_op_bits_active_vipred ? _GEN_2486 : _GEN_1772; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3663 = io_op_bits_active_vipred ? _GEN_2487 : _GEN_1773; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3664 = io_op_bits_active_vipred ? _GEN_2488 : _GEN_1774; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3665 = io_op_bits_active_vipred ? _GEN_2489 : _GEN_1775; // @[sequencer-master.scala 641:41]
  wire  _GEN_3666 = io_op_bits_active_vipred ? _GEN_2498 : _GEN_1776; // @[sequencer-master.scala 641:41]
  wire  _GEN_3667 = io_op_bits_active_vipred ? _GEN_2499 : _GEN_1777; // @[sequencer-master.scala 641:41]
  wire  _GEN_3668 = io_op_bits_active_vipred ? _GEN_2500 : _GEN_1778; // @[sequencer-master.scala 641:41]
  wire  _GEN_3669 = io_op_bits_active_vipred ? _GEN_2501 : _GEN_1779; // @[sequencer-master.scala 641:41]
  wire  _GEN_3670 = io_op_bits_active_vipred ? _GEN_2502 : _GEN_1780; // @[sequencer-master.scala 641:41]
  wire  _GEN_3671 = io_op_bits_active_vipred ? _GEN_2503 : _GEN_1781; // @[sequencer-master.scala 641:41]
  wire  _GEN_3672 = io_op_bits_active_vipred ? _GEN_2504 : _GEN_1782; // @[sequencer-master.scala 641:41]
  wire  _GEN_3673 = io_op_bits_active_vipred ? _GEN_2505 : _GEN_1783; // @[sequencer-master.scala 641:41]
  wire  _GEN_3674 = io_op_bits_active_vipred ? _GEN_2506 : _GEN_1784; // @[sequencer-master.scala 641:41]
  wire  _GEN_3675 = io_op_bits_active_vipred ? _GEN_2507 : _GEN_1785; // @[sequencer-master.scala 641:41]
  wire  _GEN_3676 = io_op_bits_active_vipred ? _GEN_2508 : _GEN_1786; // @[sequencer-master.scala 641:41]
  wire  _GEN_3677 = io_op_bits_active_vipred ? _GEN_2509 : _GEN_1787; // @[sequencer-master.scala 641:41]
  wire  _GEN_3678 = io_op_bits_active_vipred ? _GEN_2510 : _GEN_1788; // @[sequencer-master.scala 641:41]
  wire  _GEN_3679 = io_op_bits_active_vipred ? _GEN_2511 : _GEN_1789; // @[sequencer-master.scala 641:41]
  wire  _GEN_3680 = io_op_bits_active_vipred ? _GEN_2512 : _GEN_1790; // @[sequencer-master.scala 641:41]
  wire  _GEN_3681 = io_op_bits_active_vipred ? _GEN_2513 : _GEN_1791; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3682 = io_op_bits_active_vipred ? _GEN_2514 : _GEN_1792; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3683 = io_op_bits_active_vipred ? _GEN_2515 : _GEN_1793; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3684 = io_op_bits_active_vipred ? _GEN_2516 : _GEN_1794; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3685 = io_op_bits_active_vipred ? _GEN_2517 : _GEN_1795; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3686 = io_op_bits_active_vipred ? _GEN_2518 : _GEN_1796; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3687 = io_op_bits_active_vipred ? _GEN_2519 : _GEN_1797; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3688 = io_op_bits_active_vipred ? _GEN_2520 : _GEN_1798; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3689 = io_op_bits_active_vipred ? _GEN_2521 : _GEN_1799; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3690 = io_op_bits_active_vipred ? _GEN_2522 : _GEN_1800; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3691 = io_op_bits_active_vipred ? _GEN_2523 : _GEN_1801; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3692 = io_op_bits_active_vipred ? _GEN_2524 : _GEN_1802; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3693 = io_op_bits_active_vipred ? _GEN_2525 : _GEN_1803; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3694 = io_op_bits_active_vipred ? _GEN_2526 : _GEN_1804; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3695 = io_op_bits_active_vipred ? _GEN_2527 : _GEN_1805; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3696 = io_op_bits_active_vipred ? _GEN_2528 : _GEN_1806; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3697 = io_op_bits_active_vipred ? _GEN_2529 : _GEN_1807; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3698 = io_op_bits_active_vipred ? _GEN_2530 : _GEN_1808; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3699 = io_op_bits_active_vipred ? _GEN_2531 : _GEN_1809; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3700 = io_op_bits_active_vipred ? _GEN_2532 : _GEN_1810; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3701 = io_op_bits_active_vipred ? _GEN_2533 : _GEN_1811; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3702 = io_op_bits_active_vipred ? _GEN_2534 : _GEN_1812; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3703 = io_op_bits_active_vipred ? _GEN_2535 : _GEN_1813; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3704 = io_op_bits_active_vipred ? _GEN_2536 : _GEN_1814; // @[sequencer-master.scala 641:41]
  wire [63:0] _GEN_3705 = io_op_bits_active_vipred ? _GEN_2537 : _GEN_1815; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3706 = io_op_bits_active_vipred ? _GEN_2730 : e_0_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3707 = io_op_bits_active_vipred ? _GEN_2731 : e_1_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3708 = io_op_bits_active_vipred ? _GEN_2732 : e_2_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3709 = io_op_bits_active_vipred ? _GEN_2733 : e_3_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3710 = io_op_bits_active_vipred ? _GEN_2734 : e_4_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3711 = io_op_bits_active_vipred ? _GEN_2735 : e_5_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3712 = io_op_bits_active_vipred ? _GEN_2736 : e_6_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3713 = io_op_bits_active_vipred ? _GEN_2737 : e_7_base_vs3_id; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3714 = io_op_bits_active_vipred ? _GEN_2746 : e_0_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3715 = io_op_bits_active_vipred ? _GEN_2747 : e_1_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3716 = io_op_bits_active_vipred ? _GEN_2748 : e_2_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3717 = io_op_bits_active_vipred ? _GEN_2749 : e_3_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3718 = io_op_bits_active_vipred ? _GEN_2750 : e_4_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3719 = io_op_bits_active_vipred ? _GEN_2751 : e_5_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3720 = io_op_bits_active_vipred ? _GEN_2752 : e_6_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3721 = io_op_bits_active_vipred ? _GEN_2753 : e_7_base_vs3_scalar; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3722 = io_op_bits_active_vipred ? _GEN_2754 : e_0_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3723 = io_op_bits_active_vipred ? _GEN_2755 : e_1_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3724 = io_op_bits_active_vipred ? _GEN_2756 : e_2_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3725 = io_op_bits_active_vipred ? _GEN_2757 : e_3_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3726 = io_op_bits_active_vipred ? _GEN_2758 : e_4_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3727 = io_op_bits_active_vipred ? _GEN_2759 : e_5_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3728 = io_op_bits_active_vipred ? _GEN_2760 : e_6_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire  _GEN_3729 = io_op_bits_active_vipred ? _GEN_2761 : e_7_base_vs3_pred; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3730 = io_op_bits_active_vipred ? _GEN_2762 : e_0_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3731 = io_op_bits_active_vipred ? _GEN_2763 : e_1_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3732 = io_op_bits_active_vipred ? _GEN_2764 : e_2_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3733 = io_op_bits_active_vipred ? _GEN_2765 : e_3_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3734 = io_op_bits_active_vipred ? _GEN_2766 : e_4_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3735 = io_op_bits_active_vipred ? _GEN_2767 : e_5_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3736 = io_op_bits_active_vipred ? _GEN_2768 : e_6_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [1:0] _GEN_3737 = io_op_bits_active_vipred ? _GEN_2769 : e_7_base_vs3_prec; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3738 = io_op_bits_active_vipred ? _GEN_2770 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3739 = io_op_bits_active_vipred ? _GEN_2771 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3740 = io_op_bits_active_vipred ? _GEN_2772 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3741 = io_op_bits_active_vipred ? _GEN_2773 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3742 = io_op_bits_active_vipred ? _GEN_2774 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3743 = io_op_bits_active_vipred ? _GEN_2775 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3744 = io_op_bits_active_vipred ? _GEN_2776 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [7:0] _GEN_3745 = io_op_bits_active_vipred ? _GEN_2777 : 8'h0; // @[sequencer-master.scala 641:41 sequencer-master.scala 411:33]
  wire [63:0] _GEN_3746 = io_op_bits_active_vipred ? _GEN_2778 : e_0_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3747 = io_op_bits_active_vipred ? _GEN_2779 : e_1_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3748 = io_op_bits_active_vipred ? _GEN_2780 : e_2_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3749 = io_op_bits_active_vipred ? _GEN_2781 : e_3_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3750 = io_op_bits_active_vipred ? _GEN_2782 : e_4_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3751 = io_op_bits_active_vipred ? _GEN_2783 : e_5_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3752 = io_op_bits_active_vipred ? _GEN_2784 : e_6_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [63:0] _GEN_3753 = io_op_bits_active_vipred ? _GEN_2785 : e_7_sreg_ss3; // @[sequencer-master.scala 641:41 sequencer-master.scala 109:14]
  wire [7:0] _GEN_3754 = io_op_bits_active_vipred ? _GEN_2962 : _GEN_1816; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3755 = io_op_bits_active_vipred ? _GEN_2963 : _GEN_1817; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3756 = io_op_bits_active_vipred ? _GEN_2964 : _GEN_1818; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3757 = io_op_bits_active_vipred ? _GEN_2965 : _GEN_1819; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3758 = io_op_bits_active_vipred ? _GEN_2966 : _GEN_1820; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3759 = io_op_bits_active_vipred ? _GEN_2967 : _GEN_1821; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3760 = io_op_bits_active_vipred ? _GEN_2968 : _GEN_1822; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3761 = io_op_bits_active_vipred ? _GEN_2969 : _GEN_1823; // @[sequencer-master.scala 641:41]
  wire  _GEN_3762 = io_op_bits_active_vipred ? _GEN_2978 : _GEN_1824; // @[sequencer-master.scala 641:41]
  wire  _GEN_3763 = io_op_bits_active_vipred ? _GEN_2979 : _GEN_1825; // @[sequencer-master.scala 641:41]
  wire  _GEN_3764 = io_op_bits_active_vipred ? _GEN_2980 : _GEN_1826; // @[sequencer-master.scala 641:41]
  wire  _GEN_3765 = io_op_bits_active_vipred ? _GEN_2981 : _GEN_1827; // @[sequencer-master.scala 641:41]
  wire  _GEN_3766 = io_op_bits_active_vipred ? _GEN_2982 : _GEN_1828; // @[sequencer-master.scala 641:41]
  wire  _GEN_3767 = io_op_bits_active_vipred ? _GEN_2983 : _GEN_1829; // @[sequencer-master.scala 641:41]
  wire  _GEN_3768 = io_op_bits_active_vipred ? _GEN_2984 : _GEN_1830; // @[sequencer-master.scala 641:41]
  wire  _GEN_3769 = io_op_bits_active_vipred ? _GEN_2985 : _GEN_1831; // @[sequencer-master.scala 641:41]
  wire  _GEN_3770 = io_op_bits_active_vipred ? _GEN_2986 : _GEN_1832; // @[sequencer-master.scala 641:41]
  wire  _GEN_3771 = io_op_bits_active_vipred ? _GEN_2987 : _GEN_1833; // @[sequencer-master.scala 641:41]
  wire  _GEN_3772 = io_op_bits_active_vipred ? _GEN_2988 : _GEN_1834; // @[sequencer-master.scala 641:41]
  wire  _GEN_3773 = io_op_bits_active_vipred ? _GEN_2989 : _GEN_1835; // @[sequencer-master.scala 641:41]
  wire  _GEN_3774 = io_op_bits_active_vipred ? _GEN_2990 : _GEN_1836; // @[sequencer-master.scala 641:41]
  wire  _GEN_3775 = io_op_bits_active_vipred ? _GEN_2991 : _GEN_1837; // @[sequencer-master.scala 641:41]
  wire  _GEN_3776 = io_op_bits_active_vipred ? _GEN_2992 : _GEN_1838; // @[sequencer-master.scala 641:41]
  wire  _GEN_3777 = io_op_bits_active_vipred ? _GEN_2993 : _GEN_1839; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3778 = io_op_bits_active_vipred ? _GEN_2994 : _GEN_1840; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3779 = io_op_bits_active_vipred ? _GEN_2995 : _GEN_1841; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3780 = io_op_bits_active_vipred ? _GEN_2996 : _GEN_1842; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3781 = io_op_bits_active_vipred ? _GEN_2997 : _GEN_1843; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3782 = io_op_bits_active_vipred ? _GEN_2998 : _GEN_1844; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3783 = io_op_bits_active_vipred ? _GEN_2999 : _GEN_1845; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3784 = io_op_bits_active_vipred ? _GEN_3000 : _GEN_1846; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3785 = io_op_bits_active_vipred ? _GEN_3001 : _GEN_1847; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3786 = io_op_bits_active_vipred ? _GEN_3002 : _GEN_1848; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3787 = io_op_bits_active_vipred ? _GEN_3003 : _GEN_1849; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3788 = io_op_bits_active_vipred ? _GEN_3004 : _GEN_1850; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3789 = io_op_bits_active_vipred ? _GEN_3005 : _GEN_1851; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3790 = io_op_bits_active_vipred ? _GEN_3006 : _GEN_1852; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3791 = io_op_bits_active_vipred ? _GEN_3007 : _GEN_1853; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3792 = io_op_bits_active_vipred ? _GEN_3008 : _GEN_1854; // @[sequencer-master.scala 641:41]
  wire [7:0] _GEN_3793 = io_op_bits_active_vipred ? _GEN_3009 : _GEN_1855; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3794 = io_op_bits_active_vipred ? _GEN_3266 : _GEN_1856; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3795 = io_op_bits_active_vipred ? _GEN_3267 : _GEN_1857; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3796 = io_op_bits_active_vipred ? _GEN_3268 : _GEN_1858; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3797 = io_op_bits_active_vipred ? _GEN_3269 : _GEN_1859; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3798 = io_op_bits_active_vipred ? _GEN_3270 : _GEN_1860; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3799 = io_op_bits_active_vipred ? _GEN_3271 : _GEN_1861; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3800 = io_op_bits_active_vipred ? _GEN_3272 : _GEN_1862; // @[sequencer-master.scala 641:41]
  wire [1:0] _GEN_3801 = io_op_bits_active_vipred ? _GEN_3273 : _GEN_1863; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3802 = io_op_bits_active_vipred ? _GEN_3298 : _GEN_1864; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3803 = io_op_bits_active_vipred ? _GEN_3299 : _GEN_1865; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3804 = io_op_bits_active_vipred ? _GEN_3300 : _GEN_1866; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3805 = io_op_bits_active_vipred ? _GEN_3301 : _GEN_1867; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3806 = io_op_bits_active_vipred ? _GEN_3302 : _GEN_1868; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3807 = io_op_bits_active_vipred ? _GEN_3303 : _GEN_1869; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3808 = io_op_bits_active_vipred ? _GEN_3304 : _GEN_1870; // @[sequencer-master.scala 641:41]
  wire [3:0] _GEN_3809 = io_op_bits_active_vipred ? _GEN_3305 : _GEN_1871; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3810 = io_op_bits_active_vipred ? _GEN_3314 : _GEN_1872; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3811 = io_op_bits_active_vipred ? _GEN_3315 : _GEN_1873; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3812 = io_op_bits_active_vipred ? _GEN_3316 : _GEN_1874; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3813 = io_op_bits_active_vipred ? _GEN_3317 : _GEN_1875; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3814 = io_op_bits_active_vipred ? _GEN_3318 : _GEN_1876; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3815 = io_op_bits_active_vipred ? _GEN_3319 : _GEN_1877; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3816 = io_op_bits_active_vipred ? _GEN_3320 : _GEN_1878; // @[sequencer-master.scala 641:41]
  wire [2:0] _GEN_3817 = io_op_bits_active_vipred ? _GEN_3321 : _GEN_1879; // @[sequencer-master.scala 641:41]
  wire  _GEN_3818 = io_op_bits_active_vipred | io_op_bits_active_vint; // @[sequencer-master.scala 641:41 sequencer-master.scala 265:41]
  wire [2:0] _GEN_3819 = io_op_bits_active_vipred ? _T_1645 : _GEN_1881; // @[sequencer-master.scala 641:41 sequencer-master.scala 265:66]
  wire  _GEN_3820 = _GEN_32729 | _GEN_3322; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3821 = _GEN_32730 | _GEN_3323; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3822 = _GEN_32731 | _GEN_3324; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3823 = _GEN_32732 | _GEN_3325; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3824 = _GEN_32733 | _GEN_3326; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3825 = _GEN_32734 | _GEN_3327; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3826 = _GEN_32735 | _GEN_3328; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3827 = _GEN_32736 | _GEN_3329; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_3836 = 3'h0 == tail ? 1'h0 : _GEN_3338; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3837 = 3'h1 == tail ? 1'h0 : _GEN_3339; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3838 = 3'h2 == tail ? 1'h0 : _GEN_3340; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3839 = 3'h3 == tail ? 1'h0 : _GEN_3341; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3840 = 3'h4 == tail ? 1'h0 : _GEN_3342; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3841 = 3'h5 == tail ? 1'h0 : _GEN_3343; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3842 = 3'h6 == tail ? 1'h0 : _GEN_3344; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3843 = 3'h7 == tail ? 1'h0 : _GEN_3345; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_3844 = 3'h0 == tail ? 1'h0 : _GEN_3346; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3845 = 3'h1 == tail ? 1'h0 : _GEN_3347; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3846 = 3'h2 == tail ? 1'h0 : _GEN_3348; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3847 = 3'h3 == tail ? 1'h0 : _GEN_3349; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3848 = 3'h4 == tail ? 1'h0 : _GEN_3350; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3849 = 3'h5 == tail ? 1'h0 : _GEN_3351; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3850 = 3'h6 == tail ? 1'h0 : _GEN_3352; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3851 = 3'h7 == tail ? 1'h0 : _GEN_3353; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_3852 = 3'h0 == tail ? 1'h0 : _GEN_3354; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3853 = 3'h1 == tail ? 1'h0 : _GEN_3355; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3854 = 3'h2 == tail ? 1'h0 : _GEN_3356; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3855 = 3'h3 == tail ? 1'h0 : _GEN_3357; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3856 = 3'h4 == tail ? 1'h0 : _GEN_3358; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3857 = 3'h5 == tail ? 1'h0 : _GEN_3359; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3858 = 3'h6 == tail ? 1'h0 : _GEN_3360; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3859 = 3'h7 == tail ? 1'h0 : _GEN_3361; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_3860 = 3'h0 == tail ? 1'h0 : _GEN_3362; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3861 = 3'h1 == tail ? 1'h0 : _GEN_3363; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3862 = 3'h2 == tail ? 1'h0 : _GEN_3364; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3863 = 3'h3 == tail ? 1'h0 : _GEN_3365; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3864 = 3'h4 == tail ? 1'h0 : _GEN_3366; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3865 = 3'h5 == tail ? 1'h0 : _GEN_3367; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3866 = 3'h6 == tail ? 1'h0 : _GEN_3368; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3867 = 3'h7 == tail ? 1'h0 : _GEN_3369; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_3868 = 3'h0 == tail ? 1'h0 : _GEN_3370; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3869 = 3'h1 == tail ? 1'h0 : _GEN_3371; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3870 = 3'h2 == tail ? 1'h0 : _GEN_3372; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3871 = 3'h3 == tail ? 1'h0 : _GEN_3373; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3872 = 3'h4 == tail ? 1'h0 : _GEN_3374; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3873 = 3'h5 == tail ? 1'h0 : _GEN_3375; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3874 = 3'h6 == tail ? 1'h0 : _GEN_3376; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3875 = 3'h7 == tail ? 1'h0 : _GEN_3377; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_3876 = _GEN_32729 | _GEN_3378; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3877 = _GEN_32730 | _GEN_3379; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3878 = _GEN_32731 | _GEN_3380; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3879 = _GEN_32732 | _GEN_3381; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3880 = _GEN_32733 | _GEN_3382; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3881 = _GEN_32734 | _GEN_3383; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3882 = _GEN_32735 | _GEN_3384; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3883 = _GEN_32736 | _GEN_3385; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_3884 = 3'h0 == tail ? 1'h0 : _GEN_3386; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3885 = 3'h1 == tail ? 1'h0 : _GEN_3387; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3886 = 3'h2 == tail ? 1'h0 : _GEN_3388; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3887 = 3'h3 == tail ? 1'h0 : _GEN_3389; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3888 = 3'h4 == tail ? 1'h0 : _GEN_3390; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3889 = 3'h5 == tail ? 1'h0 : _GEN_3391; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3890 = 3'h6 == tail ? 1'h0 : _GEN_3392; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3891 = 3'h7 == tail ? 1'h0 : _GEN_3393; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3892 = 3'h0 == tail ? 1'h0 : _GEN_3394; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3893 = 3'h1 == tail ? 1'h0 : _GEN_3395; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3894 = 3'h2 == tail ? 1'h0 : _GEN_3396; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3895 = 3'h3 == tail ? 1'h0 : _GEN_3397; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3896 = 3'h4 == tail ? 1'h0 : _GEN_3398; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3897 = 3'h5 == tail ? 1'h0 : _GEN_3399; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3898 = 3'h6 == tail ? 1'h0 : _GEN_3400; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3899 = 3'h7 == tail ? 1'h0 : _GEN_3401; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3900 = 3'h0 == tail ? 1'h0 : _GEN_3402; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3901 = 3'h1 == tail ? 1'h0 : _GEN_3403; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3902 = 3'h2 == tail ? 1'h0 : _GEN_3404; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3903 = 3'h3 == tail ? 1'h0 : _GEN_3405; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3904 = 3'h4 == tail ? 1'h0 : _GEN_3406; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3905 = 3'h5 == tail ? 1'h0 : _GEN_3407; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3906 = 3'h6 == tail ? 1'h0 : _GEN_3408; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3907 = 3'h7 == tail ? 1'h0 : _GEN_3409; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3908 = 3'h0 == tail ? 1'h0 : _GEN_3410; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3909 = 3'h1 == tail ? 1'h0 : _GEN_3411; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3910 = 3'h2 == tail ? 1'h0 : _GEN_3412; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3911 = 3'h3 == tail ? 1'h0 : _GEN_3413; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3912 = 3'h4 == tail ? 1'h0 : _GEN_3414; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3913 = 3'h5 == tail ? 1'h0 : _GEN_3415; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3914 = 3'h6 == tail ? 1'h0 : _GEN_3416; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3915 = 3'h7 == tail ? 1'h0 : _GEN_3417; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3916 = 3'h0 == tail ? 1'h0 : _GEN_3418; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3917 = 3'h1 == tail ? 1'h0 : _GEN_3419; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3918 = 3'h2 == tail ? 1'h0 : _GEN_3420; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3919 = 3'h3 == tail ? 1'h0 : _GEN_3421; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3920 = 3'h4 == tail ? 1'h0 : _GEN_3422; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3921 = 3'h5 == tail ? 1'h0 : _GEN_3423; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3922 = 3'h6 == tail ? 1'h0 : _GEN_3424; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3923 = 3'h7 == tail ? 1'h0 : _GEN_3425; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3924 = 3'h0 == tail ? 1'h0 : _GEN_3426; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3925 = 3'h1 == tail ? 1'h0 : _GEN_3427; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3926 = 3'h2 == tail ? 1'h0 : _GEN_3428; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3927 = 3'h3 == tail ? 1'h0 : _GEN_3429; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3928 = 3'h4 == tail ? 1'h0 : _GEN_3430; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3929 = 3'h5 == tail ? 1'h0 : _GEN_3431; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3930 = 3'h6 == tail ? 1'h0 : _GEN_3432; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3931 = 3'h7 == tail ? 1'h0 : _GEN_3433; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3932 = 3'h0 == tail ? 1'h0 : _GEN_3434; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3933 = 3'h1 == tail ? 1'h0 : _GEN_3435; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3934 = 3'h2 == tail ? 1'h0 : _GEN_3436; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3935 = 3'h3 == tail ? 1'h0 : _GEN_3437; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3936 = 3'h4 == tail ? 1'h0 : _GEN_3438; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3937 = 3'h5 == tail ? 1'h0 : _GEN_3439; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3938 = 3'h6 == tail ? 1'h0 : _GEN_3440; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3939 = 3'h7 == tail ? 1'h0 : _GEN_3441; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3940 = 3'h0 == tail ? 1'h0 : _GEN_3442; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3941 = 3'h1 == tail ? 1'h0 : _GEN_3443; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3942 = 3'h2 == tail ? 1'h0 : _GEN_3444; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3943 = 3'h3 == tail ? 1'h0 : _GEN_3445; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3944 = 3'h4 == tail ? 1'h0 : _GEN_3446; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3945 = 3'h5 == tail ? 1'h0 : _GEN_3447; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3946 = 3'h6 == tail ? 1'h0 : _GEN_3448; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3947 = 3'h7 == tail ? 1'h0 : _GEN_3449; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3948 = 3'h0 == tail ? 1'h0 : _GEN_3450; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3949 = 3'h1 == tail ? 1'h0 : _GEN_3451; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3950 = 3'h2 == tail ? 1'h0 : _GEN_3452; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3951 = 3'h3 == tail ? 1'h0 : _GEN_3453; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3952 = 3'h4 == tail ? 1'h0 : _GEN_3454; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3953 = 3'h5 == tail ? 1'h0 : _GEN_3455; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3954 = 3'h6 == tail ? 1'h0 : _GEN_3456; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3955 = 3'h7 == tail ? 1'h0 : _GEN_3457; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3956 = 3'h0 == tail ? 1'h0 : _GEN_3458; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3957 = 3'h1 == tail ? 1'h0 : _GEN_3459; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3958 = 3'h2 == tail ? 1'h0 : _GEN_3460; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3959 = 3'h3 == tail ? 1'h0 : _GEN_3461; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3960 = 3'h4 == tail ? 1'h0 : _GEN_3462; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3961 = 3'h5 == tail ? 1'h0 : _GEN_3463; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3962 = 3'h6 == tail ? 1'h0 : _GEN_3464; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3963 = 3'h7 == tail ? 1'h0 : _GEN_3465; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3964 = 3'h0 == tail ? 1'h0 : _GEN_3466; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3965 = 3'h1 == tail ? 1'h0 : _GEN_3467; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3966 = 3'h2 == tail ? 1'h0 : _GEN_3468; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3967 = 3'h3 == tail ? 1'h0 : _GEN_3469; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3968 = 3'h4 == tail ? 1'h0 : _GEN_3470; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3969 = 3'h5 == tail ? 1'h0 : _GEN_3471; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3970 = 3'h6 == tail ? 1'h0 : _GEN_3472; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3971 = 3'h7 == tail ? 1'h0 : _GEN_3473; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3972 = 3'h0 == tail ? 1'h0 : _GEN_3474; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3973 = 3'h1 == tail ? 1'h0 : _GEN_3475; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3974 = 3'h2 == tail ? 1'h0 : _GEN_3476; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3975 = 3'h3 == tail ? 1'h0 : _GEN_3477; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3976 = 3'h4 == tail ? 1'h0 : _GEN_3478; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3977 = 3'h5 == tail ? 1'h0 : _GEN_3479; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3978 = 3'h6 == tail ? 1'h0 : _GEN_3480; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3979 = 3'h7 == tail ? 1'h0 : _GEN_3481; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3980 = 3'h0 == tail ? 1'h0 : _GEN_3482; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3981 = 3'h1 == tail ? 1'h0 : _GEN_3483; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3982 = 3'h2 == tail ? 1'h0 : _GEN_3484; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3983 = 3'h3 == tail ? 1'h0 : _GEN_3485; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3984 = 3'h4 == tail ? 1'h0 : _GEN_3486; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3985 = 3'h5 == tail ? 1'h0 : _GEN_3487; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3986 = 3'h6 == tail ? 1'h0 : _GEN_3488; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3987 = 3'h7 == tail ? 1'h0 : _GEN_3489; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_3988 = 3'h0 == tail ? 1'h0 : _GEN_3490; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3989 = 3'h1 == tail ? 1'h0 : _GEN_3491; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3990 = 3'h2 == tail ? 1'h0 : _GEN_3492; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3991 = 3'h3 == tail ? 1'h0 : _GEN_3493; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3992 = 3'h4 == tail ? 1'h0 : _GEN_3494; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3993 = 3'h5 == tail ? 1'h0 : _GEN_3495; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3994 = 3'h6 == tail ? 1'h0 : _GEN_3496; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3995 = 3'h7 == tail ? 1'h0 : _GEN_3497; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_3996 = 3'h0 == tail ? 1'h0 : _GEN_3498; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3997 = 3'h1 == tail ? 1'h0 : _GEN_3499; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3998 = 3'h2 == tail ? 1'h0 : _GEN_3500; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_3999 = 3'h3 == tail ? 1'h0 : _GEN_3501; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4000 = 3'h4 == tail ? 1'h0 : _GEN_3502; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4001 = 3'h5 == tail ? 1'h0 : _GEN_3503; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4002 = 3'h6 == tail ? 1'h0 : _GEN_3504; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4003 = 3'h7 == tail ? 1'h0 : _GEN_3505; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4004 = 3'h0 == tail ? 1'h0 : _GEN_3506; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4005 = 3'h1 == tail ? 1'h0 : _GEN_3507; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4006 = 3'h2 == tail ? 1'h0 : _GEN_3508; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4007 = 3'h3 == tail ? 1'h0 : _GEN_3509; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4008 = 3'h4 == tail ? 1'h0 : _GEN_3510; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4009 = 3'h5 == tail ? 1'h0 : _GEN_3511; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4010 = 3'h6 == tail ? 1'h0 : _GEN_3512; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4011 = 3'h7 == tail ? 1'h0 : _GEN_3513; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4012 = 3'h0 == tail ? 1'h0 : _GEN_3514; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4013 = 3'h1 == tail ? 1'h0 : _GEN_3515; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4014 = 3'h2 == tail ? 1'h0 : _GEN_3516; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4015 = 3'h3 == tail ? 1'h0 : _GEN_3517; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4016 = 3'h4 == tail ? 1'h0 : _GEN_3518; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4017 = 3'h5 == tail ? 1'h0 : _GEN_3519; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4018 = 3'h6 == tail ? 1'h0 : _GEN_3520; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4019 = 3'h7 == tail ? 1'h0 : _GEN_3521; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4020 = 3'h0 == tail ? 1'h0 : _GEN_3522; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4021 = 3'h1 == tail ? 1'h0 : _GEN_3523; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4022 = 3'h2 == tail ? 1'h0 : _GEN_3524; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4023 = 3'h3 == tail ? 1'h0 : _GEN_3525; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4024 = 3'h4 == tail ? 1'h0 : _GEN_3526; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4025 = 3'h5 == tail ? 1'h0 : _GEN_3527; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4026 = 3'h6 == tail ? 1'h0 : _GEN_3528; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4027 = 3'h7 == tail ? 1'h0 : _GEN_3529; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4028 = 3'h0 == tail ? 1'h0 : _GEN_3530; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4029 = 3'h1 == tail ? 1'h0 : _GEN_3531; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4030 = 3'h2 == tail ? 1'h0 : _GEN_3532; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4031 = 3'h3 == tail ? 1'h0 : _GEN_3533; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4032 = 3'h4 == tail ? 1'h0 : _GEN_3534; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4033 = 3'h5 == tail ? 1'h0 : _GEN_3535; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4034 = 3'h6 == tail ? 1'h0 : _GEN_3536; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4035 = 3'h7 == tail ? 1'h0 : _GEN_3537; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4036 = 3'h0 == tail ? 1'h0 : _GEN_3538; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4037 = 3'h1 == tail ? 1'h0 : _GEN_3539; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4038 = 3'h2 == tail ? 1'h0 : _GEN_3540; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4039 = 3'h3 == tail ? 1'h0 : _GEN_3541; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4040 = 3'h4 == tail ? 1'h0 : _GEN_3542; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4041 = 3'h5 == tail ? 1'h0 : _GEN_3543; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4042 = 3'h6 == tail ? 1'h0 : _GEN_3544; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4043 = 3'h7 == tail ? 1'h0 : _GEN_3545; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4044 = 3'h0 == tail ? 1'h0 : _GEN_3546; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4045 = 3'h1 == tail ? 1'h0 : _GEN_3547; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4046 = 3'h2 == tail ? 1'h0 : _GEN_3548; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4047 = 3'h3 == tail ? 1'h0 : _GEN_3549; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4048 = 3'h4 == tail ? 1'h0 : _GEN_3550; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4049 = 3'h5 == tail ? 1'h0 : _GEN_3551; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4050 = 3'h6 == tail ? 1'h0 : _GEN_3552; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4051 = 3'h7 == tail ? 1'h0 : _GEN_3553; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4052 = 3'h0 == tail ? 1'h0 : _GEN_3554; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4053 = 3'h1 == tail ? 1'h0 : _GEN_3555; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4054 = 3'h2 == tail ? 1'h0 : _GEN_3556; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4055 = 3'h3 == tail ? 1'h0 : _GEN_3557; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4056 = 3'h4 == tail ? 1'h0 : _GEN_3558; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4057 = 3'h5 == tail ? 1'h0 : _GEN_3559; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4058 = 3'h6 == tail ? 1'h0 : _GEN_3560; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4059 = 3'h7 == tail ? 1'h0 : _GEN_3561; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_4060 = 3'h0 == tail ? 1'h0 : _GEN_3562; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4061 = 3'h1 == tail ? 1'h0 : _GEN_3563; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4062 = 3'h2 == tail ? 1'h0 : _GEN_3564; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4063 = 3'h3 == tail ? 1'h0 : _GEN_3565; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4064 = 3'h4 == tail ? 1'h0 : _GEN_3566; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4065 = 3'h5 == tail ? 1'h0 : _GEN_3567; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4066 = 3'h6 == tail ? 1'h0 : _GEN_3568; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4067 = 3'h7 == tail ? 1'h0 : _GEN_3569; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_4068 = 3'h0 == tail ? 1'h0 : _GEN_3570; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4069 = 3'h1 == tail ? 1'h0 : _GEN_3571; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4070 = 3'h2 == tail ? 1'h0 : _GEN_3572; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4071 = 3'h3 == tail ? 1'h0 : _GEN_3573; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4072 = 3'h4 == tail ? 1'h0 : _GEN_3574; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4073 = 3'h5 == tail ? 1'h0 : _GEN_3575; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4074 = 3'h6 == tail ? 1'h0 : _GEN_3576; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4075 = 3'h7 == tail ? 1'h0 : _GEN_3577; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_4076 = 3'h0 == tail ? 1'h0 : _GEN_3578; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4077 = 3'h1 == tail ? 1'h0 : _GEN_3579; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4078 = 3'h2 == tail ? 1'h0 : _GEN_3580; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4079 = 3'h3 == tail ? 1'h0 : _GEN_3581; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4080 = 3'h4 == tail ? 1'h0 : _GEN_3582; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4081 = 3'h5 == tail ? 1'h0 : _GEN_3583; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4082 = 3'h6 == tail ? 1'h0 : _GEN_3584; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4083 = 3'h7 == tail ? 1'h0 : _GEN_3585; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_4092 = _GEN_32729 | e_0_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4093 = _GEN_32730 | e_1_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4094 = _GEN_32731 | e_2_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4095 = _GEN_32732 | e_3_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4096 = _GEN_32733 | e_4_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4097 = _GEN_32734 | e_5_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4098 = _GEN_32735 | e_6_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_4099 = _GEN_32736 | e_7_active_vimu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_4100 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_3602; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4101 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_3603; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4102 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_3604; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4103 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_3605; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4104 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_3606; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4105 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_3607; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4106 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_3608; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_4107 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_3609; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_4108 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_1688; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4109 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_1689; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4110 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_1690; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4111 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_1691; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4112 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_1692; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4113 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_1693; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4114 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_1694; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_4115 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_1695; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4116 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_3836; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4117 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_3837; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4118 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_3838; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4119 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_3839; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4120 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_3840; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4121 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_3841; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4122 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_3842; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4123 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_3843; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4124 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_1696; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4125 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_1697; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4126 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_1698; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4127 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_1699; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4128 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_1700; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4129 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_1701; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4130 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_1702; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4131 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_1703; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4132 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_1704; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4133 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_1705; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4134 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_1706; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4135 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_1707; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4136 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_1708; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4137 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_1709; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4138 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_1710; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_4139 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_1711; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_4140 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_1712; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4141 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_1713; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4142 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_1714; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4143 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_1715; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4144 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_1716; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4145 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_1717; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4146 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_1718; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_4147 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_1719; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_4148 = io_op_bits_base_vp_valid ? _GEN_4108 : _GEN_1688; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4149 = io_op_bits_base_vp_valid ? _GEN_4109 : _GEN_1689; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4150 = io_op_bits_base_vp_valid ? _GEN_4110 : _GEN_1690; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4151 = io_op_bits_base_vp_valid ? _GEN_4111 : _GEN_1691; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4152 = io_op_bits_base_vp_valid ? _GEN_4112 : _GEN_1692; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4153 = io_op_bits_base_vp_valid ? _GEN_4113 : _GEN_1693; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4154 = io_op_bits_base_vp_valid ? _GEN_4114 : _GEN_1694; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_4155 = io_op_bits_base_vp_valid ? _GEN_4115 : _GEN_1695; // @[sequencer-master.scala 320:41]
  wire  _GEN_4156 = io_op_bits_base_vp_valid ? _GEN_4116 : _GEN_3836; // @[sequencer-master.scala 320:41]
  wire  _GEN_4157 = io_op_bits_base_vp_valid ? _GEN_4117 : _GEN_3837; // @[sequencer-master.scala 320:41]
  wire  _GEN_4158 = io_op_bits_base_vp_valid ? _GEN_4118 : _GEN_3838; // @[sequencer-master.scala 320:41]
  wire  _GEN_4159 = io_op_bits_base_vp_valid ? _GEN_4119 : _GEN_3839; // @[sequencer-master.scala 320:41]
  wire  _GEN_4160 = io_op_bits_base_vp_valid ? _GEN_4120 : _GEN_3840; // @[sequencer-master.scala 320:41]
  wire  _GEN_4161 = io_op_bits_base_vp_valid ? _GEN_4121 : _GEN_3841; // @[sequencer-master.scala 320:41]
  wire  _GEN_4162 = io_op_bits_base_vp_valid ? _GEN_4122 : _GEN_3842; // @[sequencer-master.scala 320:41]
  wire  _GEN_4163 = io_op_bits_base_vp_valid ? _GEN_4123 : _GEN_3843; // @[sequencer-master.scala 320:41]
  wire  _GEN_4164 = io_op_bits_base_vp_valid ? _GEN_4124 : _GEN_1696; // @[sequencer-master.scala 320:41]
  wire  _GEN_4165 = io_op_bits_base_vp_valid ? _GEN_4125 : _GEN_1697; // @[sequencer-master.scala 320:41]
  wire  _GEN_4166 = io_op_bits_base_vp_valid ? _GEN_4126 : _GEN_1698; // @[sequencer-master.scala 320:41]
  wire  _GEN_4167 = io_op_bits_base_vp_valid ? _GEN_4127 : _GEN_1699; // @[sequencer-master.scala 320:41]
  wire  _GEN_4168 = io_op_bits_base_vp_valid ? _GEN_4128 : _GEN_1700; // @[sequencer-master.scala 320:41]
  wire  _GEN_4169 = io_op_bits_base_vp_valid ? _GEN_4129 : _GEN_1701; // @[sequencer-master.scala 320:41]
  wire  _GEN_4170 = io_op_bits_base_vp_valid ? _GEN_4130 : _GEN_1702; // @[sequencer-master.scala 320:41]
  wire  _GEN_4171 = io_op_bits_base_vp_valid ? _GEN_4131 : _GEN_1703; // @[sequencer-master.scala 320:41]
  wire  _GEN_4172 = io_op_bits_base_vp_valid ? _GEN_4132 : _GEN_1704; // @[sequencer-master.scala 320:41]
  wire  _GEN_4173 = io_op_bits_base_vp_valid ? _GEN_4133 : _GEN_1705; // @[sequencer-master.scala 320:41]
  wire  _GEN_4174 = io_op_bits_base_vp_valid ? _GEN_4134 : _GEN_1706; // @[sequencer-master.scala 320:41]
  wire  _GEN_4175 = io_op_bits_base_vp_valid ? _GEN_4135 : _GEN_1707; // @[sequencer-master.scala 320:41]
  wire  _GEN_4176 = io_op_bits_base_vp_valid ? _GEN_4136 : _GEN_1708; // @[sequencer-master.scala 320:41]
  wire  _GEN_4177 = io_op_bits_base_vp_valid ? _GEN_4137 : _GEN_1709; // @[sequencer-master.scala 320:41]
  wire  _GEN_4178 = io_op_bits_base_vp_valid ? _GEN_4138 : _GEN_1710; // @[sequencer-master.scala 320:41]
  wire  _GEN_4179 = io_op_bits_base_vp_valid ? _GEN_4139 : _GEN_1711; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4180 = io_op_bits_base_vp_valid ? _GEN_4140 : _GEN_1712; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4181 = io_op_bits_base_vp_valid ? _GEN_4141 : _GEN_1713; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4182 = io_op_bits_base_vp_valid ? _GEN_4142 : _GEN_1714; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4183 = io_op_bits_base_vp_valid ? _GEN_4143 : _GEN_1715; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4184 = io_op_bits_base_vp_valid ? _GEN_4144 : _GEN_1716; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4185 = io_op_bits_base_vp_valid ? _GEN_4145 : _GEN_1717; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4186 = io_op_bits_base_vp_valid ? _GEN_4146 : _GEN_1718; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_4187 = io_op_bits_base_vp_valid ? _GEN_4147 : _GEN_1719; // @[sequencer-master.scala 320:41]
  wire  _GEN_4188 = _GEN_32729 | _GEN_3884; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4189 = _GEN_32730 | _GEN_3885; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4190 = _GEN_32731 | _GEN_3886; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4191 = _GEN_32732 | _GEN_3887; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4192 = _GEN_32733 | _GEN_3888; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4193 = _GEN_32734 | _GEN_3889; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4194 = _GEN_32735 | _GEN_3890; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4195 = _GEN_32736 | _GEN_3891; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4196 = _T_26 ? _GEN_4188 : _GEN_3884; // @[sequencer-master.scala 154:24]
  wire  _GEN_4197 = _T_26 ? _GEN_4189 : _GEN_3885; // @[sequencer-master.scala 154:24]
  wire  _GEN_4198 = _T_26 ? _GEN_4190 : _GEN_3886; // @[sequencer-master.scala 154:24]
  wire  _GEN_4199 = _T_26 ? _GEN_4191 : _GEN_3887; // @[sequencer-master.scala 154:24]
  wire  _GEN_4200 = _T_26 ? _GEN_4192 : _GEN_3888; // @[sequencer-master.scala 154:24]
  wire  _GEN_4201 = _T_26 ? _GEN_4193 : _GEN_3889; // @[sequencer-master.scala 154:24]
  wire  _GEN_4202 = _T_26 ? _GEN_4194 : _GEN_3890; // @[sequencer-master.scala 154:24]
  wire  _GEN_4203 = _T_26 ? _GEN_4195 : _GEN_3891; // @[sequencer-master.scala 154:24]
  wire  _GEN_4204 = _GEN_32729 | _GEN_3908; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4205 = _GEN_32730 | _GEN_3909; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4206 = _GEN_32731 | _GEN_3910; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4207 = _GEN_32732 | _GEN_3911; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4208 = _GEN_32733 | _GEN_3912; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4209 = _GEN_32734 | _GEN_3913; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4210 = _GEN_32735 | _GEN_3914; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4211 = _GEN_32736 | _GEN_3915; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4212 = _T_48 ? _GEN_4204 : _GEN_3908; // @[sequencer-master.scala 154:24]
  wire  _GEN_4213 = _T_48 ? _GEN_4205 : _GEN_3909; // @[sequencer-master.scala 154:24]
  wire  _GEN_4214 = _T_48 ? _GEN_4206 : _GEN_3910; // @[sequencer-master.scala 154:24]
  wire  _GEN_4215 = _T_48 ? _GEN_4207 : _GEN_3911; // @[sequencer-master.scala 154:24]
  wire  _GEN_4216 = _T_48 ? _GEN_4208 : _GEN_3912; // @[sequencer-master.scala 154:24]
  wire  _GEN_4217 = _T_48 ? _GEN_4209 : _GEN_3913; // @[sequencer-master.scala 154:24]
  wire  _GEN_4218 = _T_48 ? _GEN_4210 : _GEN_3914; // @[sequencer-master.scala 154:24]
  wire  _GEN_4219 = _T_48 ? _GEN_4211 : _GEN_3915; // @[sequencer-master.scala 154:24]
  wire  _GEN_4220 = _GEN_32729 | _GEN_3932; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4221 = _GEN_32730 | _GEN_3933; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4222 = _GEN_32731 | _GEN_3934; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4223 = _GEN_32732 | _GEN_3935; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4224 = _GEN_32733 | _GEN_3936; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4225 = _GEN_32734 | _GEN_3937; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4226 = _GEN_32735 | _GEN_3938; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4227 = _GEN_32736 | _GEN_3939; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4228 = _T_70 ? _GEN_4220 : _GEN_3932; // @[sequencer-master.scala 154:24]
  wire  _GEN_4229 = _T_70 ? _GEN_4221 : _GEN_3933; // @[sequencer-master.scala 154:24]
  wire  _GEN_4230 = _T_70 ? _GEN_4222 : _GEN_3934; // @[sequencer-master.scala 154:24]
  wire  _GEN_4231 = _T_70 ? _GEN_4223 : _GEN_3935; // @[sequencer-master.scala 154:24]
  wire  _GEN_4232 = _T_70 ? _GEN_4224 : _GEN_3936; // @[sequencer-master.scala 154:24]
  wire  _GEN_4233 = _T_70 ? _GEN_4225 : _GEN_3937; // @[sequencer-master.scala 154:24]
  wire  _GEN_4234 = _T_70 ? _GEN_4226 : _GEN_3938; // @[sequencer-master.scala 154:24]
  wire  _GEN_4235 = _T_70 ? _GEN_4227 : _GEN_3939; // @[sequencer-master.scala 154:24]
  wire  _GEN_4236 = _GEN_32729 | _GEN_3956; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4237 = _GEN_32730 | _GEN_3957; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4238 = _GEN_32731 | _GEN_3958; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4239 = _GEN_32732 | _GEN_3959; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4240 = _GEN_32733 | _GEN_3960; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4241 = _GEN_32734 | _GEN_3961; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4242 = _GEN_32735 | _GEN_3962; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4243 = _GEN_32736 | _GEN_3963; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4244 = _T_92 ? _GEN_4236 : _GEN_3956; // @[sequencer-master.scala 154:24]
  wire  _GEN_4245 = _T_92 ? _GEN_4237 : _GEN_3957; // @[sequencer-master.scala 154:24]
  wire  _GEN_4246 = _T_92 ? _GEN_4238 : _GEN_3958; // @[sequencer-master.scala 154:24]
  wire  _GEN_4247 = _T_92 ? _GEN_4239 : _GEN_3959; // @[sequencer-master.scala 154:24]
  wire  _GEN_4248 = _T_92 ? _GEN_4240 : _GEN_3960; // @[sequencer-master.scala 154:24]
  wire  _GEN_4249 = _T_92 ? _GEN_4241 : _GEN_3961; // @[sequencer-master.scala 154:24]
  wire  _GEN_4250 = _T_92 ? _GEN_4242 : _GEN_3962; // @[sequencer-master.scala 154:24]
  wire  _GEN_4251 = _T_92 ? _GEN_4243 : _GEN_3963; // @[sequencer-master.scala 154:24]
  wire  _GEN_4252 = _GEN_32729 | _GEN_3980; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4253 = _GEN_32730 | _GEN_3981; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4254 = _GEN_32731 | _GEN_3982; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4255 = _GEN_32732 | _GEN_3983; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4256 = _GEN_32733 | _GEN_3984; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4257 = _GEN_32734 | _GEN_3985; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4258 = _GEN_32735 | _GEN_3986; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4259 = _GEN_32736 | _GEN_3987; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4260 = _T_114 ? _GEN_4252 : _GEN_3980; // @[sequencer-master.scala 154:24]
  wire  _GEN_4261 = _T_114 ? _GEN_4253 : _GEN_3981; // @[sequencer-master.scala 154:24]
  wire  _GEN_4262 = _T_114 ? _GEN_4254 : _GEN_3982; // @[sequencer-master.scala 154:24]
  wire  _GEN_4263 = _T_114 ? _GEN_4255 : _GEN_3983; // @[sequencer-master.scala 154:24]
  wire  _GEN_4264 = _T_114 ? _GEN_4256 : _GEN_3984; // @[sequencer-master.scala 154:24]
  wire  _GEN_4265 = _T_114 ? _GEN_4257 : _GEN_3985; // @[sequencer-master.scala 154:24]
  wire  _GEN_4266 = _T_114 ? _GEN_4258 : _GEN_3986; // @[sequencer-master.scala 154:24]
  wire  _GEN_4267 = _T_114 ? _GEN_4259 : _GEN_3987; // @[sequencer-master.scala 154:24]
  wire  _GEN_4268 = _GEN_32729 | _GEN_4004; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4269 = _GEN_32730 | _GEN_4005; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4270 = _GEN_32731 | _GEN_4006; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4271 = _GEN_32732 | _GEN_4007; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4272 = _GEN_32733 | _GEN_4008; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4273 = _GEN_32734 | _GEN_4009; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4274 = _GEN_32735 | _GEN_4010; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4275 = _GEN_32736 | _GEN_4011; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4276 = _T_136 ? _GEN_4268 : _GEN_4004; // @[sequencer-master.scala 154:24]
  wire  _GEN_4277 = _T_136 ? _GEN_4269 : _GEN_4005; // @[sequencer-master.scala 154:24]
  wire  _GEN_4278 = _T_136 ? _GEN_4270 : _GEN_4006; // @[sequencer-master.scala 154:24]
  wire  _GEN_4279 = _T_136 ? _GEN_4271 : _GEN_4007; // @[sequencer-master.scala 154:24]
  wire  _GEN_4280 = _T_136 ? _GEN_4272 : _GEN_4008; // @[sequencer-master.scala 154:24]
  wire  _GEN_4281 = _T_136 ? _GEN_4273 : _GEN_4009; // @[sequencer-master.scala 154:24]
  wire  _GEN_4282 = _T_136 ? _GEN_4274 : _GEN_4010; // @[sequencer-master.scala 154:24]
  wire  _GEN_4283 = _T_136 ? _GEN_4275 : _GEN_4011; // @[sequencer-master.scala 154:24]
  wire  _GEN_4284 = _GEN_32729 | _GEN_4028; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4285 = _GEN_32730 | _GEN_4029; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4286 = _GEN_32731 | _GEN_4030; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4287 = _GEN_32732 | _GEN_4031; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4288 = _GEN_32733 | _GEN_4032; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4289 = _GEN_32734 | _GEN_4033; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4290 = _GEN_32735 | _GEN_4034; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4291 = _GEN_32736 | _GEN_4035; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4292 = _T_158 ? _GEN_4284 : _GEN_4028; // @[sequencer-master.scala 154:24]
  wire  _GEN_4293 = _T_158 ? _GEN_4285 : _GEN_4029; // @[sequencer-master.scala 154:24]
  wire  _GEN_4294 = _T_158 ? _GEN_4286 : _GEN_4030; // @[sequencer-master.scala 154:24]
  wire  _GEN_4295 = _T_158 ? _GEN_4287 : _GEN_4031; // @[sequencer-master.scala 154:24]
  wire  _GEN_4296 = _T_158 ? _GEN_4288 : _GEN_4032; // @[sequencer-master.scala 154:24]
  wire  _GEN_4297 = _T_158 ? _GEN_4289 : _GEN_4033; // @[sequencer-master.scala 154:24]
  wire  _GEN_4298 = _T_158 ? _GEN_4290 : _GEN_4034; // @[sequencer-master.scala 154:24]
  wire  _GEN_4299 = _T_158 ? _GEN_4291 : _GEN_4035; // @[sequencer-master.scala 154:24]
  wire  _GEN_4300 = _GEN_32729 | _GEN_4052; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4301 = _GEN_32730 | _GEN_4053; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4302 = _GEN_32731 | _GEN_4054; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4303 = _GEN_32732 | _GEN_4055; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4304 = _GEN_32733 | _GEN_4056; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4305 = _GEN_32734 | _GEN_4057; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4306 = _GEN_32735 | _GEN_4058; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4307 = _GEN_32736 | _GEN_4059; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4308 = _T_180 ? _GEN_4300 : _GEN_4052; // @[sequencer-master.scala 154:24]
  wire  _GEN_4309 = _T_180 ? _GEN_4301 : _GEN_4053; // @[sequencer-master.scala 154:24]
  wire  _GEN_4310 = _T_180 ? _GEN_4302 : _GEN_4054; // @[sequencer-master.scala 154:24]
  wire  _GEN_4311 = _T_180 ? _GEN_4303 : _GEN_4055; // @[sequencer-master.scala 154:24]
  wire  _GEN_4312 = _T_180 ? _GEN_4304 : _GEN_4056; // @[sequencer-master.scala 154:24]
  wire  _GEN_4313 = _T_180 ? _GEN_4305 : _GEN_4057; // @[sequencer-master.scala 154:24]
  wire  _GEN_4314 = _T_180 ? _GEN_4306 : _GEN_4058; // @[sequencer-master.scala 154:24]
  wire  _GEN_4315 = _T_180 ? _GEN_4307 : _GEN_4059; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_4316 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_3610; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4317 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_3611; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4318 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_3612; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4319 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_3613; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4320 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_3614; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4321 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_3615; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4322 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_3616; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4323 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_3617; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4324 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_3844; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4325 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_3845; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4326 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_3846; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4327 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_3847; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4328 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_3848; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4329 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_3849; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4330 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_3850; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4331 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_3851; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4332 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_3618; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4333 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_3619; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4334 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_3620; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4335 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_3621; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4336 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_3622; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4337 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_3623; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4338 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_3624; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4339 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_3625; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4340 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_3626; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4341 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_3627; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4342 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_3628; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4343 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_3629; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4344 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_3630; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4345 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_3631; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4346 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_3632; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4347 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_3633; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4348 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_3634; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4349 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_3635; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4350 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_3636; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4351 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_3637; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4352 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_3638; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4353 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_3639; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4354 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_3640; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4355 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_3641; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4356 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_3642; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4357 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_3643; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4358 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_3644; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4359 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_3645; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4360 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_3646; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4361 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_3647; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4362 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_3648; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4363 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_3649; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_4364 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_3650; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4365 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_3651; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4366 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_3652; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4367 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_3653; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4368 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_3654; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4369 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_3655; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4370 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_3656; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4371 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_3657; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4372 = _T_189 ? _GEN_4364 : _GEN_3650; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4373 = _T_189 ? _GEN_4365 : _GEN_3651; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4374 = _T_189 ? _GEN_4366 : _GEN_3652; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4375 = _T_189 ? _GEN_4367 : _GEN_3653; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4376 = _T_189 ? _GEN_4368 : _GEN_3654; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4377 = _T_189 ? _GEN_4369 : _GEN_3655; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4378 = _T_189 ? _GEN_4370 : _GEN_3656; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4379 = _T_189 ? _GEN_4371 : _GEN_3657; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_4380 = io_op_bits_base_vs1_valid ? _GEN_4316 : _GEN_3610; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4381 = io_op_bits_base_vs1_valid ? _GEN_4317 : _GEN_3611; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4382 = io_op_bits_base_vs1_valid ? _GEN_4318 : _GEN_3612; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4383 = io_op_bits_base_vs1_valid ? _GEN_4319 : _GEN_3613; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4384 = io_op_bits_base_vs1_valid ? _GEN_4320 : _GEN_3614; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4385 = io_op_bits_base_vs1_valid ? _GEN_4321 : _GEN_3615; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4386 = io_op_bits_base_vs1_valid ? _GEN_4322 : _GEN_3616; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4387 = io_op_bits_base_vs1_valid ? _GEN_4323 : _GEN_3617; // @[sequencer-master.scala 328:47]
  wire  _GEN_4388 = io_op_bits_base_vs1_valid ? _GEN_4324 : _GEN_3844; // @[sequencer-master.scala 328:47]
  wire  _GEN_4389 = io_op_bits_base_vs1_valid ? _GEN_4325 : _GEN_3845; // @[sequencer-master.scala 328:47]
  wire  _GEN_4390 = io_op_bits_base_vs1_valid ? _GEN_4326 : _GEN_3846; // @[sequencer-master.scala 328:47]
  wire  _GEN_4391 = io_op_bits_base_vs1_valid ? _GEN_4327 : _GEN_3847; // @[sequencer-master.scala 328:47]
  wire  _GEN_4392 = io_op_bits_base_vs1_valid ? _GEN_4328 : _GEN_3848; // @[sequencer-master.scala 328:47]
  wire  _GEN_4393 = io_op_bits_base_vs1_valid ? _GEN_4329 : _GEN_3849; // @[sequencer-master.scala 328:47]
  wire  _GEN_4394 = io_op_bits_base_vs1_valid ? _GEN_4330 : _GEN_3850; // @[sequencer-master.scala 328:47]
  wire  _GEN_4395 = io_op_bits_base_vs1_valid ? _GEN_4331 : _GEN_3851; // @[sequencer-master.scala 328:47]
  wire  _GEN_4396 = io_op_bits_base_vs1_valid ? _GEN_4332 : _GEN_3618; // @[sequencer-master.scala 328:47]
  wire  _GEN_4397 = io_op_bits_base_vs1_valid ? _GEN_4333 : _GEN_3619; // @[sequencer-master.scala 328:47]
  wire  _GEN_4398 = io_op_bits_base_vs1_valid ? _GEN_4334 : _GEN_3620; // @[sequencer-master.scala 328:47]
  wire  _GEN_4399 = io_op_bits_base_vs1_valid ? _GEN_4335 : _GEN_3621; // @[sequencer-master.scala 328:47]
  wire  _GEN_4400 = io_op_bits_base_vs1_valid ? _GEN_4336 : _GEN_3622; // @[sequencer-master.scala 328:47]
  wire  _GEN_4401 = io_op_bits_base_vs1_valid ? _GEN_4337 : _GEN_3623; // @[sequencer-master.scala 328:47]
  wire  _GEN_4402 = io_op_bits_base_vs1_valid ? _GEN_4338 : _GEN_3624; // @[sequencer-master.scala 328:47]
  wire  _GEN_4403 = io_op_bits_base_vs1_valid ? _GEN_4339 : _GEN_3625; // @[sequencer-master.scala 328:47]
  wire  _GEN_4404 = io_op_bits_base_vs1_valid ? _GEN_4340 : _GEN_3626; // @[sequencer-master.scala 328:47]
  wire  _GEN_4405 = io_op_bits_base_vs1_valid ? _GEN_4341 : _GEN_3627; // @[sequencer-master.scala 328:47]
  wire  _GEN_4406 = io_op_bits_base_vs1_valid ? _GEN_4342 : _GEN_3628; // @[sequencer-master.scala 328:47]
  wire  _GEN_4407 = io_op_bits_base_vs1_valid ? _GEN_4343 : _GEN_3629; // @[sequencer-master.scala 328:47]
  wire  _GEN_4408 = io_op_bits_base_vs1_valid ? _GEN_4344 : _GEN_3630; // @[sequencer-master.scala 328:47]
  wire  _GEN_4409 = io_op_bits_base_vs1_valid ? _GEN_4345 : _GEN_3631; // @[sequencer-master.scala 328:47]
  wire  _GEN_4410 = io_op_bits_base_vs1_valid ? _GEN_4346 : _GEN_3632; // @[sequencer-master.scala 328:47]
  wire  _GEN_4411 = io_op_bits_base_vs1_valid ? _GEN_4347 : _GEN_3633; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4412 = io_op_bits_base_vs1_valid ? _GEN_4348 : _GEN_3634; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4413 = io_op_bits_base_vs1_valid ? _GEN_4349 : _GEN_3635; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4414 = io_op_bits_base_vs1_valid ? _GEN_4350 : _GEN_3636; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4415 = io_op_bits_base_vs1_valid ? _GEN_4351 : _GEN_3637; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4416 = io_op_bits_base_vs1_valid ? _GEN_4352 : _GEN_3638; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4417 = io_op_bits_base_vs1_valid ? _GEN_4353 : _GEN_3639; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4418 = io_op_bits_base_vs1_valid ? _GEN_4354 : _GEN_3640; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4419 = io_op_bits_base_vs1_valid ? _GEN_4355 : _GEN_3641; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4420 = io_op_bits_base_vs1_valid ? _GEN_4356 : _GEN_3642; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4421 = io_op_bits_base_vs1_valid ? _GEN_4357 : _GEN_3643; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4422 = io_op_bits_base_vs1_valid ? _GEN_4358 : _GEN_3644; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4423 = io_op_bits_base_vs1_valid ? _GEN_4359 : _GEN_3645; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4424 = io_op_bits_base_vs1_valid ? _GEN_4360 : _GEN_3646; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4425 = io_op_bits_base_vs1_valid ? _GEN_4361 : _GEN_3647; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4426 = io_op_bits_base_vs1_valid ? _GEN_4362 : _GEN_3648; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4427 = io_op_bits_base_vs1_valid ? _GEN_4363 : _GEN_3649; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4428 = io_op_bits_base_vs1_valid ? _GEN_4372 : _GEN_3650; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4429 = io_op_bits_base_vs1_valid ? _GEN_4373 : _GEN_3651; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4430 = io_op_bits_base_vs1_valid ? _GEN_4374 : _GEN_3652; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4431 = io_op_bits_base_vs1_valid ? _GEN_4375 : _GEN_3653; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4432 = io_op_bits_base_vs1_valid ? _GEN_4376 : _GEN_3654; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4433 = io_op_bits_base_vs1_valid ? _GEN_4377 : _GEN_3655; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4434 = io_op_bits_base_vs1_valid ? _GEN_4378 : _GEN_3656; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4435 = io_op_bits_base_vs1_valid ? _GEN_4379 : _GEN_3657; // @[sequencer-master.scala 328:47]
  wire  _GEN_4436 = _GEN_32729 | _GEN_4196; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4437 = _GEN_32730 | _GEN_4197; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4438 = _GEN_32731 | _GEN_4198; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4439 = _GEN_32732 | _GEN_4199; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4440 = _GEN_32733 | _GEN_4200; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4441 = _GEN_32734 | _GEN_4201; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4442 = _GEN_32735 | _GEN_4202; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4443 = _GEN_32736 | _GEN_4203; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4444 = _T_203 ? _GEN_4436 : _GEN_4196; // @[sequencer-master.scala 154:24]
  wire  _GEN_4445 = _T_203 ? _GEN_4437 : _GEN_4197; // @[sequencer-master.scala 154:24]
  wire  _GEN_4446 = _T_203 ? _GEN_4438 : _GEN_4198; // @[sequencer-master.scala 154:24]
  wire  _GEN_4447 = _T_203 ? _GEN_4439 : _GEN_4199; // @[sequencer-master.scala 154:24]
  wire  _GEN_4448 = _T_203 ? _GEN_4440 : _GEN_4200; // @[sequencer-master.scala 154:24]
  wire  _GEN_4449 = _T_203 ? _GEN_4441 : _GEN_4201; // @[sequencer-master.scala 154:24]
  wire  _GEN_4450 = _T_203 ? _GEN_4442 : _GEN_4202; // @[sequencer-master.scala 154:24]
  wire  _GEN_4451 = _T_203 ? _GEN_4443 : _GEN_4203; // @[sequencer-master.scala 154:24]
  wire  _GEN_4452 = _GEN_32729 | _GEN_4212; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4453 = _GEN_32730 | _GEN_4213; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4454 = _GEN_32731 | _GEN_4214; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4455 = _GEN_32732 | _GEN_4215; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4456 = _GEN_32733 | _GEN_4216; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4457 = _GEN_32734 | _GEN_4217; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4458 = _GEN_32735 | _GEN_4218; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4459 = _GEN_32736 | _GEN_4219; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4460 = _T_225 ? _GEN_4452 : _GEN_4212; // @[sequencer-master.scala 154:24]
  wire  _GEN_4461 = _T_225 ? _GEN_4453 : _GEN_4213; // @[sequencer-master.scala 154:24]
  wire  _GEN_4462 = _T_225 ? _GEN_4454 : _GEN_4214; // @[sequencer-master.scala 154:24]
  wire  _GEN_4463 = _T_225 ? _GEN_4455 : _GEN_4215; // @[sequencer-master.scala 154:24]
  wire  _GEN_4464 = _T_225 ? _GEN_4456 : _GEN_4216; // @[sequencer-master.scala 154:24]
  wire  _GEN_4465 = _T_225 ? _GEN_4457 : _GEN_4217; // @[sequencer-master.scala 154:24]
  wire  _GEN_4466 = _T_225 ? _GEN_4458 : _GEN_4218; // @[sequencer-master.scala 154:24]
  wire  _GEN_4467 = _T_225 ? _GEN_4459 : _GEN_4219; // @[sequencer-master.scala 154:24]
  wire  _GEN_4468 = _GEN_32729 | _GEN_4228; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4469 = _GEN_32730 | _GEN_4229; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4470 = _GEN_32731 | _GEN_4230; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4471 = _GEN_32732 | _GEN_4231; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4472 = _GEN_32733 | _GEN_4232; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4473 = _GEN_32734 | _GEN_4233; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4474 = _GEN_32735 | _GEN_4234; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4475 = _GEN_32736 | _GEN_4235; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4476 = _T_247 ? _GEN_4468 : _GEN_4228; // @[sequencer-master.scala 154:24]
  wire  _GEN_4477 = _T_247 ? _GEN_4469 : _GEN_4229; // @[sequencer-master.scala 154:24]
  wire  _GEN_4478 = _T_247 ? _GEN_4470 : _GEN_4230; // @[sequencer-master.scala 154:24]
  wire  _GEN_4479 = _T_247 ? _GEN_4471 : _GEN_4231; // @[sequencer-master.scala 154:24]
  wire  _GEN_4480 = _T_247 ? _GEN_4472 : _GEN_4232; // @[sequencer-master.scala 154:24]
  wire  _GEN_4481 = _T_247 ? _GEN_4473 : _GEN_4233; // @[sequencer-master.scala 154:24]
  wire  _GEN_4482 = _T_247 ? _GEN_4474 : _GEN_4234; // @[sequencer-master.scala 154:24]
  wire  _GEN_4483 = _T_247 ? _GEN_4475 : _GEN_4235; // @[sequencer-master.scala 154:24]
  wire  _GEN_4484 = _GEN_32729 | _GEN_4244; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4485 = _GEN_32730 | _GEN_4245; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4486 = _GEN_32731 | _GEN_4246; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4487 = _GEN_32732 | _GEN_4247; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4488 = _GEN_32733 | _GEN_4248; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4489 = _GEN_32734 | _GEN_4249; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4490 = _GEN_32735 | _GEN_4250; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4491 = _GEN_32736 | _GEN_4251; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4492 = _T_269 ? _GEN_4484 : _GEN_4244; // @[sequencer-master.scala 154:24]
  wire  _GEN_4493 = _T_269 ? _GEN_4485 : _GEN_4245; // @[sequencer-master.scala 154:24]
  wire  _GEN_4494 = _T_269 ? _GEN_4486 : _GEN_4246; // @[sequencer-master.scala 154:24]
  wire  _GEN_4495 = _T_269 ? _GEN_4487 : _GEN_4247; // @[sequencer-master.scala 154:24]
  wire  _GEN_4496 = _T_269 ? _GEN_4488 : _GEN_4248; // @[sequencer-master.scala 154:24]
  wire  _GEN_4497 = _T_269 ? _GEN_4489 : _GEN_4249; // @[sequencer-master.scala 154:24]
  wire  _GEN_4498 = _T_269 ? _GEN_4490 : _GEN_4250; // @[sequencer-master.scala 154:24]
  wire  _GEN_4499 = _T_269 ? _GEN_4491 : _GEN_4251; // @[sequencer-master.scala 154:24]
  wire  _GEN_4500 = _GEN_32729 | _GEN_4260; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4501 = _GEN_32730 | _GEN_4261; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4502 = _GEN_32731 | _GEN_4262; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4503 = _GEN_32732 | _GEN_4263; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4504 = _GEN_32733 | _GEN_4264; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4505 = _GEN_32734 | _GEN_4265; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4506 = _GEN_32735 | _GEN_4266; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4507 = _GEN_32736 | _GEN_4267; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4508 = _T_291 ? _GEN_4500 : _GEN_4260; // @[sequencer-master.scala 154:24]
  wire  _GEN_4509 = _T_291 ? _GEN_4501 : _GEN_4261; // @[sequencer-master.scala 154:24]
  wire  _GEN_4510 = _T_291 ? _GEN_4502 : _GEN_4262; // @[sequencer-master.scala 154:24]
  wire  _GEN_4511 = _T_291 ? _GEN_4503 : _GEN_4263; // @[sequencer-master.scala 154:24]
  wire  _GEN_4512 = _T_291 ? _GEN_4504 : _GEN_4264; // @[sequencer-master.scala 154:24]
  wire  _GEN_4513 = _T_291 ? _GEN_4505 : _GEN_4265; // @[sequencer-master.scala 154:24]
  wire  _GEN_4514 = _T_291 ? _GEN_4506 : _GEN_4266; // @[sequencer-master.scala 154:24]
  wire  _GEN_4515 = _T_291 ? _GEN_4507 : _GEN_4267; // @[sequencer-master.scala 154:24]
  wire  _GEN_4516 = _GEN_32729 | _GEN_4276; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4517 = _GEN_32730 | _GEN_4277; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4518 = _GEN_32731 | _GEN_4278; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4519 = _GEN_32732 | _GEN_4279; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4520 = _GEN_32733 | _GEN_4280; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4521 = _GEN_32734 | _GEN_4281; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4522 = _GEN_32735 | _GEN_4282; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4523 = _GEN_32736 | _GEN_4283; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4524 = _T_313 ? _GEN_4516 : _GEN_4276; // @[sequencer-master.scala 154:24]
  wire  _GEN_4525 = _T_313 ? _GEN_4517 : _GEN_4277; // @[sequencer-master.scala 154:24]
  wire  _GEN_4526 = _T_313 ? _GEN_4518 : _GEN_4278; // @[sequencer-master.scala 154:24]
  wire  _GEN_4527 = _T_313 ? _GEN_4519 : _GEN_4279; // @[sequencer-master.scala 154:24]
  wire  _GEN_4528 = _T_313 ? _GEN_4520 : _GEN_4280; // @[sequencer-master.scala 154:24]
  wire  _GEN_4529 = _T_313 ? _GEN_4521 : _GEN_4281; // @[sequencer-master.scala 154:24]
  wire  _GEN_4530 = _T_313 ? _GEN_4522 : _GEN_4282; // @[sequencer-master.scala 154:24]
  wire  _GEN_4531 = _T_313 ? _GEN_4523 : _GEN_4283; // @[sequencer-master.scala 154:24]
  wire  _GEN_4532 = _GEN_32729 | _GEN_4292; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4533 = _GEN_32730 | _GEN_4293; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4534 = _GEN_32731 | _GEN_4294; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4535 = _GEN_32732 | _GEN_4295; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4536 = _GEN_32733 | _GEN_4296; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4537 = _GEN_32734 | _GEN_4297; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4538 = _GEN_32735 | _GEN_4298; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4539 = _GEN_32736 | _GEN_4299; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4540 = _T_335 ? _GEN_4532 : _GEN_4292; // @[sequencer-master.scala 154:24]
  wire  _GEN_4541 = _T_335 ? _GEN_4533 : _GEN_4293; // @[sequencer-master.scala 154:24]
  wire  _GEN_4542 = _T_335 ? _GEN_4534 : _GEN_4294; // @[sequencer-master.scala 154:24]
  wire  _GEN_4543 = _T_335 ? _GEN_4535 : _GEN_4295; // @[sequencer-master.scala 154:24]
  wire  _GEN_4544 = _T_335 ? _GEN_4536 : _GEN_4296; // @[sequencer-master.scala 154:24]
  wire  _GEN_4545 = _T_335 ? _GEN_4537 : _GEN_4297; // @[sequencer-master.scala 154:24]
  wire  _GEN_4546 = _T_335 ? _GEN_4538 : _GEN_4298; // @[sequencer-master.scala 154:24]
  wire  _GEN_4547 = _T_335 ? _GEN_4539 : _GEN_4299; // @[sequencer-master.scala 154:24]
  wire  _GEN_4548 = _GEN_32729 | _GEN_4308; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4549 = _GEN_32730 | _GEN_4309; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4550 = _GEN_32731 | _GEN_4310; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4551 = _GEN_32732 | _GEN_4311; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4552 = _GEN_32733 | _GEN_4312; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4553 = _GEN_32734 | _GEN_4313; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4554 = _GEN_32735 | _GEN_4314; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4555 = _GEN_32736 | _GEN_4315; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4556 = _T_357 ? _GEN_4548 : _GEN_4308; // @[sequencer-master.scala 154:24]
  wire  _GEN_4557 = _T_357 ? _GEN_4549 : _GEN_4309; // @[sequencer-master.scala 154:24]
  wire  _GEN_4558 = _T_357 ? _GEN_4550 : _GEN_4310; // @[sequencer-master.scala 154:24]
  wire  _GEN_4559 = _T_357 ? _GEN_4551 : _GEN_4311; // @[sequencer-master.scala 154:24]
  wire  _GEN_4560 = _T_357 ? _GEN_4552 : _GEN_4312; // @[sequencer-master.scala 154:24]
  wire  _GEN_4561 = _T_357 ? _GEN_4553 : _GEN_4313; // @[sequencer-master.scala 154:24]
  wire  _GEN_4562 = _T_357 ? _GEN_4554 : _GEN_4314; // @[sequencer-master.scala 154:24]
  wire  _GEN_4563 = _T_357 ? _GEN_4555 : _GEN_4315; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_4564 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_3658; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4565 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_3659; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4566 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_3660; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4567 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_3661; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4568 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_3662; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4569 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_3663; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4570 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_3664; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4571 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_3665; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4572 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_3852; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4573 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_3853; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4574 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_3854; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4575 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_3855; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4576 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_3856; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4577 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_3857; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4578 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_3858; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4579 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_3859; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4580 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_3666; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4581 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_3667; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4582 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_3668; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4583 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_3669; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4584 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_3670; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4585 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_3671; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4586 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_3672; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4587 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_3673; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4588 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_3674; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4589 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_3675; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4590 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_3676; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4591 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_3677; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4592 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_3678; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4593 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_3679; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4594 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_3680; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_4595 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_3681; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4596 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_3682; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4597 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_3683; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4598 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_3684; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4599 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_3685; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4600 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_3686; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4601 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_3687; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4602 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_3688; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_4603 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_3689; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_4604 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_3690; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4605 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_3691; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4606 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_3692; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4607 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_3693; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4608 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_3694; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4609 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_3695; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4610 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_3696; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_4611 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_3697; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_4612 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_3698; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4613 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_3699; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4614 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_3700; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4615 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_3701; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4616 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_3702; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4617 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_3703; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4618 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_3704; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4619 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_3705; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_4620 = _T_366 ? _GEN_4612 : _GEN_3698; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4621 = _T_366 ? _GEN_4613 : _GEN_3699; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4622 = _T_366 ? _GEN_4614 : _GEN_3700; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4623 = _T_366 ? _GEN_4615 : _GEN_3701; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4624 = _T_366 ? _GEN_4616 : _GEN_3702; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4625 = _T_366 ? _GEN_4617 : _GEN_3703; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4626 = _T_366 ? _GEN_4618 : _GEN_3704; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_4627 = _T_366 ? _GEN_4619 : _GEN_3705; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_4628 = io_op_bits_base_vs2_valid ? _GEN_4564 : _GEN_3658; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4629 = io_op_bits_base_vs2_valid ? _GEN_4565 : _GEN_3659; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4630 = io_op_bits_base_vs2_valid ? _GEN_4566 : _GEN_3660; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4631 = io_op_bits_base_vs2_valid ? _GEN_4567 : _GEN_3661; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4632 = io_op_bits_base_vs2_valid ? _GEN_4568 : _GEN_3662; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4633 = io_op_bits_base_vs2_valid ? _GEN_4569 : _GEN_3663; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4634 = io_op_bits_base_vs2_valid ? _GEN_4570 : _GEN_3664; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4635 = io_op_bits_base_vs2_valid ? _GEN_4571 : _GEN_3665; // @[sequencer-master.scala 328:47]
  wire  _GEN_4636 = io_op_bits_base_vs2_valid ? _GEN_4572 : _GEN_3852; // @[sequencer-master.scala 328:47]
  wire  _GEN_4637 = io_op_bits_base_vs2_valid ? _GEN_4573 : _GEN_3853; // @[sequencer-master.scala 328:47]
  wire  _GEN_4638 = io_op_bits_base_vs2_valid ? _GEN_4574 : _GEN_3854; // @[sequencer-master.scala 328:47]
  wire  _GEN_4639 = io_op_bits_base_vs2_valid ? _GEN_4575 : _GEN_3855; // @[sequencer-master.scala 328:47]
  wire  _GEN_4640 = io_op_bits_base_vs2_valid ? _GEN_4576 : _GEN_3856; // @[sequencer-master.scala 328:47]
  wire  _GEN_4641 = io_op_bits_base_vs2_valid ? _GEN_4577 : _GEN_3857; // @[sequencer-master.scala 328:47]
  wire  _GEN_4642 = io_op_bits_base_vs2_valid ? _GEN_4578 : _GEN_3858; // @[sequencer-master.scala 328:47]
  wire  _GEN_4643 = io_op_bits_base_vs2_valid ? _GEN_4579 : _GEN_3859; // @[sequencer-master.scala 328:47]
  wire  _GEN_4644 = io_op_bits_base_vs2_valid ? _GEN_4580 : _GEN_3666; // @[sequencer-master.scala 328:47]
  wire  _GEN_4645 = io_op_bits_base_vs2_valid ? _GEN_4581 : _GEN_3667; // @[sequencer-master.scala 328:47]
  wire  _GEN_4646 = io_op_bits_base_vs2_valid ? _GEN_4582 : _GEN_3668; // @[sequencer-master.scala 328:47]
  wire  _GEN_4647 = io_op_bits_base_vs2_valid ? _GEN_4583 : _GEN_3669; // @[sequencer-master.scala 328:47]
  wire  _GEN_4648 = io_op_bits_base_vs2_valid ? _GEN_4584 : _GEN_3670; // @[sequencer-master.scala 328:47]
  wire  _GEN_4649 = io_op_bits_base_vs2_valid ? _GEN_4585 : _GEN_3671; // @[sequencer-master.scala 328:47]
  wire  _GEN_4650 = io_op_bits_base_vs2_valid ? _GEN_4586 : _GEN_3672; // @[sequencer-master.scala 328:47]
  wire  _GEN_4651 = io_op_bits_base_vs2_valid ? _GEN_4587 : _GEN_3673; // @[sequencer-master.scala 328:47]
  wire  _GEN_4652 = io_op_bits_base_vs2_valid ? _GEN_4588 : _GEN_3674; // @[sequencer-master.scala 328:47]
  wire  _GEN_4653 = io_op_bits_base_vs2_valid ? _GEN_4589 : _GEN_3675; // @[sequencer-master.scala 328:47]
  wire  _GEN_4654 = io_op_bits_base_vs2_valid ? _GEN_4590 : _GEN_3676; // @[sequencer-master.scala 328:47]
  wire  _GEN_4655 = io_op_bits_base_vs2_valid ? _GEN_4591 : _GEN_3677; // @[sequencer-master.scala 328:47]
  wire  _GEN_4656 = io_op_bits_base_vs2_valid ? _GEN_4592 : _GEN_3678; // @[sequencer-master.scala 328:47]
  wire  _GEN_4657 = io_op_bits_base_vs2_valid ? _GEN_4593 : _GEN_3679; // @[sequencer-master.scala 328:47]
  wire  _GEN_4658 = io_op_bits_base_vs2_valid ? _GEN_4594 : _GEN_3680; // @[sequencer-master.scala 328:47]
  wire  _GEN_4659 = io_op_bits_base_vs2_valid ? _GEN_4595 : _GEN_3681; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4660 = io_op_bits_base_vs2_valid ? _GEN_4596 : _GEN_3682; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4661 = io_op_bits_base_vs2_valid ? _GEN_4597 : _GEN_3683; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4662 = io_op_bits_base_vs2_valid ? _GEN_4598 : _GEN_3684; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4663 = io_op_bits_base_vs2_valid ? _GEN_4599 : _GEN_3685; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4664 = io_op_bits_base_vs2_valid ? _GEN_4600 : _GEN_3686; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4665 = io_op_bits_base_vs2_valid ? _GEN_4601 : _GEN_3687; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4666 = io_op_bits_base_vs2_valid ? _GEN_4602 : _GEN_3688; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_4667 = io_op_bits_base_vs2_valid ? _GEN_4603 : _GEN_3689; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4668 = io_op_bits_base_vs2_valid ? _GEN_4604 : _GEN_3690; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4669 = io_op_bits_base_vs2_valid ? _GEN_4605 : _GEN_3691; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4670 = io_op_bits_base_vs2_valid ? _GEN_4606 : _GEN_3692; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4671 = io_op_bits_base_vs2_valid ? _GEN_4607 : _GEN_3693; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4672 = io_op_bits_base_vs2_valid ? _GEN_4608 : _GEN_3694; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4673 = io_op_bits_base_vs2_valid ? _GEN_4609 : _GEN_3695; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4674 = io_op_bits_base_vs2_valid ? _GEN_4610 : _GEN_3696; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_4675 = io_op_bits_base_vs2_valid ? _GEN_4611 : _GEN_3697; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4676 = io_op_bits_base_vs2_valid ? _GEN_4620 : _GEN_3698; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4677 = io_op_bits_base_vs2_valid ? _GEN_4621 : _GEN_3699; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4678 = io_op_bits_base_vs2_valid ? _GEN_4622 : _GEN_3700; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4679 = io_op_bits_base_vs2_valid ? _GEN_4623 : _GEN_3701; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4680 = io_op_bits_base_vs2_valid ? _GEN_4624 : _GEN_3702; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4681 = io_op_bits_base_vs2_valid ? _GEN_4625 : _GEN_3703; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4682 = io_op_bits_base_vs2_valid ? _GEN_4626 : _GEN_3704; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_4683 = io_op_bits_base_vs2_valid ? _GEN_4627 : _GEN_3705; // @[sequencer-master.scala 328:47]
  wire  _GEN_4684 = _GEN_32729 | _GEN_4444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4685 = _GEN_32730 | _GEN_4445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4686 = _GEN_32731 | _GEN_4446; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4687 = _GEN_32732 | _GEN_4447; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4688 = _GEN_32733 | _GEN_4448; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4689 = _GEN_32734 | _GEN_4449; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4690 = _GEN_32735 | _GEN_4450; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4691 = _GEN_32736 | _GEN_4451; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4692 = _T_380 ? _GEN_4684 : _GEN_4444; // @[sequencer-master.scala 154:24]
  wire  _GEN_4693 = _T_380 ? _GEN_4685 : _GEN_4445; // @[sequencer-master.scala 154:24]
  wire  _GEN_4694 = _T_380 ? _GEN_4686 : _GEN_4446; // @[sequencer-master.scala 154:24]
  wire  _GEN_4695 = _T_380 ? _GEN_4687 : _GEN_4447; // @[sequencer-master.scala 154:24]
  wire  _GEN_4696 = _T_380 ? _GEN_4688 : _GEN_4448; // @[sequencer-master.scala 154:24]
  wire  _GEN_4697 = _T_380 ? _GEN_4689 : _GEN_4449; // @[sequencer-master.scala 154:24]
  wire  _GEN_4698 = _T_380 ? _GEN_4690 : _GEN_4450; // @[sequencer-master.scala 154:24]
  wire  _GEN_4699 = _T_380 ? _GEN_4691 : _GEN_4451; // @[sequencer-master.scala 154:24]
  wire  _GEN_4700 = _GEN_32729 | _GEN_4460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4701 = _GEN_32730 | _GEN_4461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4702 = _GEN_32731 | _GEN_4462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4703 = _GEN_32732 | _GEN_4463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4704 = _GEN_32733 | _GEN_4464; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4705 = _GEN_32734 | _GEN_4465; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4706 = _GEN_32735 | _GEN_4466; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4707 = _GEN_32736 | _GEN_4467; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4708 = _T_402 ? _GEN_4700 : _GEN_4460; // @[sequencer-master.scala 154:24]
  wire  _GEN_4709 = _T_402 ? _GEN_4701 : _GEN_4461; // @[sequencer-master.scala 154:24]
  wire  _GEN_4710 = _T_402 ? _GEN_4702 : _GEN_4462; // @[sequencer-master.scala 154:24]
  wire  _GEN_4711 = _T_402 ? _GEN_4703 : _GEN_4463; // @[sequencer-master.scala 154:24]
  wire  _GEN_4712 = _T_402 ? _GEN_4704 : _GEN_4464; // @[sequencer-master.scala 154:24]
  wire  _GEN_4713 = _T_402 ? _GEN_4705 : _GEN_4465; // @[sequencer-master.scala 154:24]
  wire  _GEN_4714 = _T_402 ? _GEN_4706 : _GEN_4466; // @[sequencer-master.scala 154:24]
  wire  _GEN_4715 = _T_402 ? _GEN_4707 : _GEN_4467; // @[sequencer-master.scala 154:24]
  wire  _GEN_4716 = _GEN_32729 | _GEN_4476; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4717 = _GEN_32730 | _GEN_4477; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4718 = _GEN_32731 | _GEN_4478; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4719 = _GEN_32732 | _GEN_4479; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4720 = _GEN_32733 | _GEN_4480; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4721 = _GEN_32734 | _GEN_4481; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4722 = _GEN_32735 | _GEN_4482; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4723 = _GEN_32736 | _GEN_4483; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4724 = _T_424 ? _GEN_4716 : _GEN_4476; // @[sequencer-master.scala 154:24]
  wire  _GEN_4725 = _T_424 ? _GEN_4717 : _GEN_4477; // @[sequencer-master.scala 154:24]
  wire  _GEN_4726 = _T_424 ? _GEN_4718 : _GEN_4478; // @[sequencer-master.scala 154:24]
  wire  _GEN_4727 = _T_424 ? _GEN_4719 : _GEN_4479; // @[sequencer-master.scala 154:24]
  wire  _GEN_4728 = _T_424 ? _GEN_4720 : _GEN_4480; // @[sequencer-master.scala 154:24]
  wire  _GEN_4729 = _T_424 ? _GEN_4721 : _GEN_4481; // @[sequencer-master.scala 154:24]
  wire  _GEN_4730 = _T_424 ? _GEN_4722 : _GEN_4482; // @[sequencer-master.scala 154:24]
  wire  _GEN_4731 = _T_424 ? _GEN_4723 : _GEN_4483; // @[sequencer-master.scala 154:24]
  wire  _GEN_4732 = _GEN_32729 | _GEN_4492; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4733 = _GEN_32730 | _GEN_4493; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4734 = _GEN_32731 | _GEN_4494; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4735 = _GEN_32732 | _GEN_4495; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4736 = _GEN_32733 | _GEN_4496; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4737 = _GEN_32734 | _GEN_4497; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4738 = _GEN_32735 | _GEN_4498; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4739 = _GEN_32736 | _GEN_4499; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4740 = _T_446 ? _GEN_4732 : _GEN_4492; // @[sequencer-master.scala 154:24]
  wire  _GEN_4741 = _T_446 ? _GEN_4733 : _GEN_4493; // @[sequencer-master.scala 154:24]
  wire  _GEN_4742 = _T_446 ? _GEN_4734 : _GEN_4494; // @[sequencer-master.scala 154:24]
  wire  _GEN_4743 = _T_446 ? _GEN_4735 : _GEN_4495; // @[sequencer-master.scala 154:24]
  wire  _GEN_4744 = _T_446 ? _GEN_4736 : _GEN_4496; // @[sequencer-master.scala 154:24]
  wire  _GEN_4745 = _T_446 ? _GEN_4737 : _GEN_4497; // @[sequencer-master.scala 154:24]
  wire  _GEN_4746 = _T_446 ? _GEN_4738 : _GEN_4498; // @[sequencer-master.scala 154:24]
  wire  _GEN_4747 = _T_446 ? _GEN_4739 : _GEN_4499; // @[sequencer-master.scala 154:24]
  wire  _GEN_4748 = _GEN_32729 | _GEN_4508; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4749 = _GEN_32730 | _GEN_4509; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4750 = _GEN_32731 | _GEN_4510; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4751 = _GEN_32732 | _GEN_4511; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4752 = _GEN_32733 | _GEN_4512; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4753 = _GEN_32734 | _GEN_4513; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4754 = _GEN_32735 | _GEN_4514; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4755 = _GEN_32736 | _GEN_4515; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4756 = _T_468 ? _GEN_4748 : _GEN_4508; // @[sequencer-master.scala 154:24]
  wire  _GEN_4757 = _T_468 ? _GEN_4749 : _GEN_4509; // @[sequencer-master.scala 154:24]
  wire  _GEN_4758 = _T_468 ? _GEN_4750 : _GEN_4510; // @[sequencer-master.scala 154:24]
  wire  _GEN_4759 = _T_468 ? _GEN_4751 : _GEN_4511; // @[sequencer-master.scala 154:24]
  wire  _GEN_4760 = _T_468 ? _GEN_4752 : _GEN_4512; // @[sequencer-master.scala 154:24]
  wire  _GEN_4761 = _T_468 ? _GEN_4753 : _GEN_4513; // @[sequencer-master.scala 154:24]
  wire  _GEN_4762 = _T_468 ? _GEN_4754 : _GEN_4514; // @[sequencer-master.scala 154:24]
  wire  _GEN_4763 = _T_468 ? _GEN_4755 : _GEN_4515; // @[sequencer-master.scala 154:24]
  wire  _GEN_4764 = _GEN_32729 | _GEN_4524; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4765 = _GEN_32730 | _GEN_4525; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4766 = _GEN_32731 | _GEN_4526; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4767 = _GEN_32732 | _GEN_4527; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4768 = _GEN_32733 | _GEN_4528; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4769 = _GEN_32734 | _GEN_4529; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4770 = _GEN_32735 | _GEN_4530; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4771 = _GEN_32736 | _GEN_4531; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4772 = _T_490 ? _GEN_4764 : _GEN_4524; // @[sequencer-master.scala 154:24]
  wire  _GEN_4773 = _T_490 ? _GEN_4765 : _GEN_4525; // @[sequencer-master.scala 154:24]
  wire  _GEN_4774 = _T_490 ? _GEN_4766 : _GEN_4526; // @[sequencer-master.scala 154:24]
  wire  _GEN_4775 = _T_490 ? _GEN_4767 : _GEN_4527; // @[sequencer-master.scala 154:24]
  wire  _GEN_4776 = _T_490 ? _GEN_4768 : _GEN_4528; // @[sequencer-master.scala 154:24]
  wire  _GEN_4777 = _T_490 ? _GEN_4769 : _GEN_4529; // @[sequencer-master.scala 154:24]
  wire  _GEN_4778 = _T_490 ? _GEN_4770 : _GEN_4530; // @[sequencer-master.scala 154:24]
  wire  _GEN_4779 = _T_490 ? _GEN_4771 : _GEN_4531; // @[sequencer-master.scala 154:24]
  wire  _GEN_4780 = _GEN_32729 | _GEN_4540; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4781 = _GEN_32730 | _GEN_4541; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4782 = _GEN_32731 | _GEN_4542; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4783 = _GEN_32732 | _GEN_4543; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4784 = _GEN_32733 | _GEN_4544; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4785 = _GEN_32734 | _GEN_4545; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4786 = _GEN_32735 | _GEN_4546; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4787 = _GEN_32736 | _GEN_4547; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4788 = _T_512 ? _GEN_4780 : _GEN_4540; // @[sequencer-master.scala 154:24]
  wire  _GEN_4789 = _T_512 ? _GEN_4781 : _GEN_4541; // @[sequencer-master.scala 154:24]
  wire  _GEN_4790 = _T_512 ? _GEN_4782 : _GEN_4542; // @[sequencer-master.scala 154:24]
  wire  _GEN_4791 = _T_512 ? _GEN_4783 : _GEN_4543; // @[sequencer-master.scala 154:24]
  wire  _GEN_4792 = _T_512 ? _GEN_4784 : _GEN_4544; // @[sequencer-master.scala 154:24]
  wire  _GEN_4793 = _T_512 ? _GEN_4785 : _GEN_4545; // @[sequencer-master.scala 154:24]
  wire  _GEN_4794 = _T_512 ? _GEN_4786 : _GEN_4546; // @[sequencer-master.scala 154:24]
  wire  _GEN_4795 = _T_512 ? _GEN_4787 : _GEN_4547; // @[sequencer-master.scala 154:24]
  wire  _GEN_4796 = _GEN_32729 | _GEN_4556; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4797 = _GEN_32730 | _GEN_4557; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4798 = _GEN_32731 | _GEN_4558; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4799 = _GEN_32732 | _GEN_4559; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4800 = _GEN_32733 | _GEN_4560; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4801 = _GEN_32734 | _GEN_4561; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4802 = _GEN_32735 | _GEN_4562; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4803 = _GEN_32736 | _GEN_4563; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_4804 = _T_534 ? _GEN_4796 : _GEN_4556; // @[sequencer-master.scala 154:24]
  wire  _GEN_4805 = _T_534 ? _GEN_4797 : _GEN_4557; // @[sequencer-master.scala 154:24]
  wire  _GEN_4806 = _T_534 ? _GEN_4798 : _GEN_4558; // @[sequencer-master.scala 154:24]
  wire  _GEN_4807 = _T_534 ? _GEN_4799 : _GEN_4559; // @[sequencer-master.scala 154:24]
  wire  _GEN_4808 = _T_534 ? _GEN_4800 : _GEN_4560; // @[sequencer-master.scala 154:24]
  wire  _GEN_4809 = _T_534 ? _GEN_4801 : _GEN_4561; // @[sequencer-master.scala 154:24]
  wire  _GEN_4810 = _T_534 ? _GEN_4802 : _GEN_4562; // @[sequencer-master.scala 154:24]
  wire  _GEN_4811 = _T_534 ? _GEN_4803 : _GEN_4563; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_4812 = 3'h0 == tail ? io_op_bits_base_vd_id : _GEN_3754; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4813 = 3'h1 == tail ? io_op_bits_base_vd_id : _GEN_3755; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4814 = 3'h2 == tail ? io_op_bits_base_vd_id : _GEN_3756; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4815 = 3'h3 == tail ? io_op_bits_base_vd_id : _GEN_3757; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4816 = 3'h4 == tail ? io_op_bits_base_vd_id : _GEN_3758; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4817 = 3'h5 == tail ? io_op_bits_base_vd_id : _GEN_3759; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4818 = 3'h6 == tail ? io_op_bits_base_vd_id : _GEN_3760; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4819 = 3'h7 == tail ? io_op_bits_base_vd_id : _GEN_3761; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4820 = 3'h0 == tail ? io_op_bits_base_vd_valid : _GEN_3868; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4821 = 3'h1 == tail ? io_op_bits_base_vd_valid : _GEN_3869; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4822 = 3'h2 == tail ? io_op_bits_base_vd_valid : _GEN_3870; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4823 = 3'h3 == tail ? io_op_bits_base_vd_valid : _GEN_3871; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4824 = 3'h4 == tail ? io_op_bits_base_vd_valid : _GEN_3872; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4825 = 3'h5 == tail ? io_op_bits_base_vd_valid : _GEN_3873; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4826 = 3'h6 == tail ? io_op_bits_base_vd_valid : _GEN_3874; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4827 = 3'h7 == tail ? io_op_bits_base_vd_valid : _GEN_3875; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4828 = 3'h0 == tail ? io_op_bits_base_vd_scalar : _GEN_3762; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4829 = 3'h1 == tail ? io_op_bits_base_vd_scalar : _GEN_3763; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4830 = 3'h2 == tail ? io_op_bits_base_vd_scalar : _GEN_3764; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4831 = 3'h3 == tail ? io_op_bits_base_vd_scalar : _GEN_3765; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4832 = 3'h4 == tail ? io_op_bits_base_vd_scalar : _GEN_3766; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4833 = 3'h5 == tail ? io_op_bits_base_vd_scalar : _GEN_3767; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4834 = 3'h6 == tail ? io_op_bits_base_vd_scalar : _GEN_3768; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4835 = 3'h7 == tail ? io_op_bits_base_vd_scalar : _GEN_3769; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4836 = 3'h0 == tail ? io_op_bits_base_vd_pred : _GEN_3770; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4837 = 3'h1 == tail ? io_op_bits_base_vd_pred : _GEN_3771; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4838 = 3'h2 == tail ? io_op_bits_base_vd_pred : _GEN_3772; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4839 = 3'h3 == tail ? io_op_bits_base_vd_pred : _GEN_3773; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4840 = 3'h4 == tail ? io_op_bits_base_vd_pred : _GEN_3774; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4841 = 3'h5 == tail ? io_op_bits_base_vd_pred : _GEN_3775; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4842 = 3'h6 == tail ? io_op_bits_base_vd_pred : _GEN_3776; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_4843 = 3'h7 == tail ? io_op_bits_base_vd_pred : _GEN_3777; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4844 = 3'h0 == tail ? io_op_bits_base_vd_prec : _GEN_3778; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4845 = 3'h1 == tail ? io_op_bits_base_vd_prec : _GEN_3779; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4846 = 3'h2 == tail ? io_op_bits_base_vd_prec : _GEN_3780; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4847 = 3'h3 == tail ? io_op_bits_base_vd_prec : _GEN_3781; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4848 = 3'h4 == tail ? io_op_bits_base_vd_prec : _GEN_3782; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4849 = 3'h5 == tail ? io_op_bits_base_vd_prec : _GEN_3783; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4850 = 3'h6 == tail ? io_op_bits_base_vd_prec : _GEN_3784; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_4851 = 3'h7 == tail ? io_op_bits_base_vd_prec : _GEN_3785; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_4852 = 3'h0 == tail ? io_op_bits_reg_vd_id : _GEN_3786; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4853 = 3'h1 == tail ? io_op_bits_reg_vd_id : _GEN_3787; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4854 = 3'h2 == tail ? io_op_bits_reg_vd_id : _GEN_3788; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4855 = 3'h3 == tail ? io_op_bits_reg_vd_id : _GEN_3789; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4856 = 3'h4 == tail ? io_op_bits_reg_vd_id : _GEN_3790; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4857 = 3'h5 == tail ? io_op_bits_reg_vd_id : _GEN_3791; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4858 = 3'h6 == tail ? io_op_bits_reg_vd_id : _GEN_3792; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4859 = 3'h7 == tail ? io_op_bits_reg_vd_id : _GEN_3793; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_4860 = io_op_bits_base_vd_valid ? _GEN_4812 : _GEN_3754; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4861 = io_op_bits_base_vd_valid ? _GEN_4813 : _GEN_3755; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4862 = io_op_bits_base_vd_valid ? _GEN_4814 : _GEN_3756; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4863 = io_op_bits_base_vd_valid ? _GEN_4815 : _GEN_3757; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4864 = io_op_bits_base_vd_valid ? _GEN_4816 : _GEN_3758; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4865 = io_op_bits_base_vd_valid ? _GEN_4817 : _GEN_3759; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4866 = io_op_bits_base_vd_valid ? _GEN_4818 : _GEN_3760; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4867 = io_op_bits_base_vd_valid ? _GEN_4819 : _GEN_3761; // @[sequencer-master.scala 362:41]
  wire  _GEN_4868 = io_op_bits_base_vd_valid ? _GEN_4820 : _GEN_3868; // @[sequencer-master.scala 362:41]
  wire  _GEN_4869 = io_op_bits_base_vd_valid ? _GEN_4821 : _GEN_3869; // @[sequencer-master.scala 362:41]
  wire  _GEN_4870 = io_op_bits_base_vd_valid ? _GEN_4822 : _GEN_3870; // @[sequencer-master.scala 362:41]
  wire  _GEN_4871 = io_op_bits_base_vd_valid ? _GEN_4823 : _GEN_3871; // @[sequencer-master.scala 362:41]
  wire  _GEN_4872 = io_op_bits_base_vd_valid ? _GEN_4824 : _GEN_3872; // @[sequencer-master.scala 362:41]
  wire  _GEN_4873 = io_op_bits_base_vd_valid ? _GEN_4825 : _GEN_3873; // @[sequencer-master.scala 362:41]
  wire  _GEN_4874 = io_op_bits_base_vd_valid ? _GEN_4826 : _GEN_3874; // @[sequencer-master.scala 362:41]
  wire  _GEN_4875 = io_op_bits_base_vd_valid ? _GEN_4827 : _GEN_3875; // @[sequencer-master.scala 362:41]
  wire  _GEN_4876 = io_op_bits_base_vd_valid ? _GEN_4828 : _GEN_3762; // @[sequencer-master.scala 362:41]
  wire  _GEN_4877 = io_op_bits_base_vd_valid ? _GEN_4829 : _GEN_3763; // @[sequencer-master.scala 362:41]
  wire  _GEN_4878 = io_op_bits_base_vd_valid ? _GEN_4830 : _GEN_3764; // @[sequencer-master.scala 362:41]
  wire  _GEN_4879 = io_op_bits_base_vd_valid ? _GEN_4831 : _GEN_3765; // @[sequencer-master.scala 362:41]
  wire  _GEN_4880 = io_op_bits_base_vd_valid ? _GEN_4832 : _GEN_3766; // @[sequencer-master.scala 362:41]
  wire  _GEN_4881 = io_op_bits_base_vd_valid ? _GEN_4833 : _GEN_3767; // @[sequencer-master.scala 362:41]
  wire  _GEN_4882 = io_op_bits_base_vd_valid ? _GEN_4834 : _GEN_3768; // @[sequencer-master.scala 362:41]
  wire  _GEN_4883 = io_op_bits_base_vd_valid ? _GEN_4835 : _GEN_3769; // @[sequencer-master.scala 362:41]
  wire  _GEN_4884 = io_op_bits_base_vd_valid ? _GEN_4836 : _GEN_3770; // @[sequencer-master.scala 362:41]
  wire  _GEN_4885 = io_op_bits_base_vd_valid ? _GEN_4837 : _GEN_3771; // @[sequencer-master.scala 362:41]
  wire  _GEN_4886 = io_op_bits_base_vd_valid ? _GEN_4838 : _GEN_3772; // @[sequencer-master.scala 362:41]
  wire  _GEN_4887 = io_op_bits_base_vd_valid ? _GEN_4839 : _GEN_3773; // @[sequencer-master.scala 362:41]
  wire  _GEN_4888 = io_op_bits_base_vd_valid ? _GEN_4840 : _GEN_3774; // @[sequencer-master.scala 362:41]
  wire  _GEN_4889 = io_op_bits_base_vd_valid ? _GEN_4841 : _GEN_3775; // @[sequencer-master.scala 362:41]
  wire  _GEN_4890 = io_op_bits_base_vd_valid ? _GEN_4842 : _GEN_3776; // @[sequencer-master.scala 362:41]
  wire  _GEN_4891 = io_op_bits_base_vd_valid ? _GEN_4843 : _GEN_3777; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4892 = io_op_bits_base_vd_valid ? _GEN_4844 : _GEN_3778; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4893 = io_op_bits_base_vd_valid ? _GEN_4845 : _GEN_3779; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4894 = io_op_bits_base_vd_valid ? _GEN_4846 : _GEN_3780; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4895 = io_op_bits_base_vd_valid ? _GEN_4847 : _GEN_3781; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4896 = io_op_bits_base_vd_valid ? _GEN_4848 : _GEN_3782; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4897 = io_op_bits_base_vd_valid ? _GEN_4849 : _GEN_3783; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4898 = io_op_bits_base_vd_valid ? _GEN_4850 : _GEN_3784; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_4899 = io_op_bits_base_vd_valid ? _GEN_4851 : _GEN_3785; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4900 = io_op_bits_base_vd_valid ? _GEN_4852 : _GEN_3786; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4901 = io_op_bits_base_vd_valid ? _GEN_4853 : _GEN_3787; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4902 = io_op_bits_base_vd_valid ? _GEN_4854 : _GEN_3788; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4903 = io_op_bits_base_vd_valid ? _GEN_4855 : _GEN_3789; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4904 = io_op_bits_base_vd_valid ? _GEN_4856 : _GEN_3790; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4905 = io_op_bits_base_vd_valid ? _GEN_4857 : _GEN_3791; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4906 = io_op_bits_base_vd_valid ? _GEN_4858 : _GEN_3792; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_4907 = io_op_bits_base_vd_valid ? _GEN_4859 : _GEN_3793; // @[sequencer-master.scala 362:41]
  wire  _GEN_4908 = _GEN_32729 | _GEN_3892; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4909 = _GEN_32730 | _GEN_3893; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4910 = _GEN_32731 | _GEN_3894; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4911 = _GEN_32732 | _GEN_3895; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4912 = _GEN_32733 | _GEN_3896; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4913 = _GEN_32734 | _GEN_3897; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4914 = _GEN_32735 | _GEN_3898; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4915 = _GEN_32736 | _GEN_3899; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4916 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4908 : _GEN_3892; // @[sequencer-master.scala 161:86]
  wire  _GEN_4917 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4909 : _GEN_3893; // @[sequencer-master.scala 161:86]
  wire  _GEN_4918 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4910 : _GEN_3894; // @[sequencer-master.scala 161:86]
  wire  _GEN_4919 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4911 : _GEN_3895; // @[sequencer-master.scala 161:86]
  wire  _GEN_4920 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4912 : _GEN_3896; // @[sequencer-master.scala 161:86]
  wire  _GEN_4921 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4913 : _GEN_3897; // @[sequencer-master.scala 161:86]
  wire  _GEN_4922 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4914 : _GEN_3898; // @[sequencer-master.scala 161:86]
  wire  _GEN_4923 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_4915 : _GEN_3899; // @[sequencer-master.scala 161:86]
  wire  _GEN_4924 = _GEN_32729 | _GEN_3916; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4925 = _GEN_32730 | _GEN_3917; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4926 = _GEN_32731 | _GEN_3918; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4927 = _GEN_32732 | _GEN_3919; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4928 = _GEN_32733 | _GEN_3920; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4929 = _GEN_32734 | _GEN_3921; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4930 = _GEN_32735 | _GEN_3922; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4931 = _GEN_32736 | _GEN_3923; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4932 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4924 : _GEN_3916; // @[sequencer-master.scala 161:86]
  wire  _GEN_4933 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4925 : _GEN_3917; // @[sequencer-master.scala 161:86]
  wire  _GEN_4934 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4926 : _GEN_3918; // @[sequencer-master.scala 161:86]
  wire  _GEN_4935 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4927 : _GEN_3919; // @[sequencer-master.scala 161:86]
  wire  _GEN_4936 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4928 : _GEN_3920; // @[sequencer-master.scala 161:86]
  wire  _GEN_4937 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4929 : _GEN_3921; // @[sequencer-master.scala 161:86]
  wire  _GEN_4938 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4930 : _GEN_3922; // @[sequencer-master.scala 161:86]
  wire  _GEN_4939 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_4931 : _GEN_3923; // @[sequencer-master.scala 161:86]
  wire  _GEN_4940 = _GEN_32729 | _GEN_3940; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4941 = _GEN_32730 | _GEN_3941; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4942 = _GEN_32731 | _GEN_3942; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4943 = _GEN_32732 | _GEN_3943; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4944 = _GEN_32733 | _GEN_3944; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4945 = _GEN_32734 | _GEN_3945; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4946 = _GEN_32735 | _GEN_3946; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4947 = _GEN_32736 | _GEN_3947; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4948 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4940 : _GEN_3940; // @[sequencer-master.scala 161:86]
  wire  _GEN_4949 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4941 : _GEN_3941; // @[sequencer-master.scala 161:86]
  wire  _GEN_4950 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4942 : _GEN_3942; // @[sequencer-master.scala 161:86]
  wire  _GEN_4951 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4943 : _GEN_3943; // @[sequencer-master.scala 161:86]
  wire  _GEN_4952 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4944 : _GEN_3944; // @[sequencer-master.scala 161:86]
  wire  _GEN_4953 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4945 : _GEN_3945; // @[sequencer-master.scala 161:86]
  wire  _GEN_4954 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4946 : _GEN_3946; // @[sequencer-master.scala 161:86]
  wire  _GEN_4955 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_4947 : _GEN_3947; // @[sequencer-master.scala 161:86]
  wire  _GEN_4956 = _GEN_32729 | _GEN_3964; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4957 = _GEN_32730 | _GEN_3965; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4958 = _GEN_32731 | _GEN_3966; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4959 = _GEN_32732 | _GEN_3967; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4960 = _GEN_32733 | _GEN_3968; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4961 = _GEN_32734 | _GEN_3969; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4962 = _GEN_32735 | _GEN_3970; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4963 = _GEN_32736 | _GEN_3971; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4964 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4956 : _GEN_3964; // @[sequencer-master.scala 161:86]
  wire  _GEN_4965 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4957 : _GEN_3965; // @[sequencer-master.scala 161:86]
  wire  _GEN_4966 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4958 : _GEN_3966; // @[sequencer-master.scala 161:86]
  wire  _GEN_4967 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4959 : _GEN_3967; // @[sequencer-master.scala 161:86]
  wire  _GEN_4968 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4960 : _GEN_3968; // @[sequencer-master.scala 161:86]
  wire  _GEN_4969 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4961 : _GEN_3969; // @[sequencer-master.scala 161:86]
  wire  _GEN_4970 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4962 : _GEN_3970; // @[sequencer-master.scala 161:86]
  wire  _GEN_4971 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_4963 : _GEN_3971; // @[sequencer-master.scala 161:86]
  wire  _GEN_4972 = _GEN_32729 | _GEN_3988; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4973 = _GEN_32730 | _GEN_3989; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4974 = _GEN_32731 | _GEN_3990; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4975 = _GEN_32732 | _GEN_3991; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4976 = _GEN_32733 | _GEN_3992; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4977 = _GEN_32734 | _GEN_3993; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4978 = _GEN_32735 | _GEN_3994; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4979 = _GEN_32736 | _GEN_3995; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4980 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4972 : _GEN_3988; // @[sequencer-master.scala 161:86]
  wire  _GEN_4981 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4973 : _GEN_3989; // @[sequencer-master.scala 161:86]
  wire  _GEN_4982 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4974 : _GEN_3990; // @[sequencer-master.scala 161:86]
  wire  _GEN_4983 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4975 : _GEN_3991; // @[sequencer-master.scala 161:86]
  wire  _GEN_4984 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4976 : _GEN_3992; // @[sequencer-master.scala 161:86]
  wire  _GEN_4985 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4977 : _GEN_3993; // @[sequencer-master.scala 161:86]
  wire  _GEN_4986 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4978 : _GEN_3994; // @[sequencer-master.scala 161:86]
  wire  _GEN_4987 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_4979 : _GEN_3995; // @[sequencer-master.scala 161:86]
  wire  _GEN_4988 = _GEN_32729 | _GEN_4012; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4989 = _GEN_32730 | _GEN_4013; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4990 = _GEN_32731 | _GEN_4014; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4991 = _GEN_32732 | _GEN_4015; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4992 = _GEN_32733 | _GEN_4016; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4993 = _GEN_32734 | _GEN_4017; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4994 = _GEN_32735 | _GEN_4018; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4995 = _GEN_32736 | _GEN_4019; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_4996 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4988 : _GEN_4012; // @[sequencer-master.scala 161:86]
  wire  _GEN_4997 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4989 : _GEN_4013; // @[sequencer-master.scala 161:86]
  wire  _GEN_4998 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4990 : _GEN_4014; // @[sequencer-master.scala 161:86]
  wire  _GEN_4999 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4991 : _GEN_4015; // @[sequencer-master.scala 161:86]
  wire  _GEN_5000 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4992 : _GEN_4016; // @[sequencer-master.scala 161:86]
  wire  _GEN_5001 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4993 : _GEN_4017; // @[sequencer-master.scala 161:86]
  wire  _GEN_5002 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4994 : _GEN_4018; // @[sequencer-master.scala 161:86]
  wire  _GEN_5003 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_4995 : _GEN_4019; // @[sequencer-master.scala 161:86]
  wire  _GEN_5004 = _GEN_32729 | _GEN_4036; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5005 = _GEN_32730 | _GEN_4037; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5006 = _GEN_32731 | _GEN_4038; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5007 = _GEN_32732 | _GEN_4039; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5008 = _GEN_32733 | _GEN_4040; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5009 = _GEN_32734 | _GEN_4041; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5010 = _GEN_32735 | _GEN_4042; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5011 = _GEN_32736 | _GEN_4043; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5012 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5004 : _GEN_4036; // @[sequencer-master.scala 161:86]
  wire  _GEN_5013 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5005 : _GEN_4037; // @[sequencer-master.scala 161:86]
  wire  _GEN_5014 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5006 : _GEN_4038; // @[sequencer-master.scala 161:86]
  wire  _GEN_5015 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5007 : _GEN_4039; // @[sequencer-master.scala 161:86]
  wire  _GEN_5016 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5008 : _GEN_4040; // @[sequencer-master.scala 161:86]
  wire  _GEN_5017 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5009 : _GEN_4041; // @[sequencer-master.scala 161:86]
  wire  _GEN_5018 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5010 : _GEN_4042; // @[sequencer-master.scala 161:86]
  wire  _GEN_5019 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_5011 : _GEN_4043; // @[sequencer-master.scala 161:86]
  wire  _GEN_5020 = _GEN_32729 | _GEN_4060; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5021 = _GEN_32730 | _GEN_4061; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5022 = _GEN_32731 | _GEN_4062; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5023 = _GEN_32732 | _GEN_4063; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5024 = _GEN_32733 | _GEN_4064; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5025 = _GEN_32734 | _GEN_4065; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5026 = _GEN_32735 | _GEN_4066; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5027 = _GEN_32736 | _GEN_4067; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_5028 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5020 : _GEN_4060; // @[sequencer-master.scala 161:86]
  wire  _GEN_5029 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5021 : _GEN_4061; // @[sequencer-master.scala 161:86]
  wire  _GEN_5030 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5022 : _GEN_4062; // @[sequencer-master.scala 161:86]
  wire  _GEN_5031 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5023 : _GEN_4063; // @[sequencer-master.scala 161:86]
  wire  _GEN_5032 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5024 : _GEN_4064; // @[sequencer-master.scala 161:86]
  wire  _GEN_5033 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5025 : _GEN_4065; // @[sequencer-master.scala 161:86]
  wire  _GEN_5034 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5026 : _GEN_4066; // @[sequencer-master.scala 161:86]
  wire  _GEN_5035 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_5027 : _GEN_4067; // @[sequencer-master.scala 161:86]
  wire  _GEN_5036 = _GEN_32729 | _GEN_3900; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5037 = _GEN_32730 | _GEN_3901; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5038 = _GEN_32731 | _GEN_3902; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5039 = _GEN_32732 | _GEN_3903; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5040 = _GEN_32733 | _GEN_3904; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5041 = _GEN_32734 | _GEN_3905; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5042 = _GEN_32735 | _GEN_3906; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5043 = _GEN_32736 | _GEN_3907; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5044 = _T_1442 ? _GEN_5036 : _GEN_3900; // @[sequencer-master.scala 168:32]
  wire  _GEN_5045 = _T_1442 ? _GEN_5037 : _GEN_3901; // @[sequencer-master.scala 168:32]
  wire  _GEN_5046 = _T_1442 ? _GEN_5038 : _GEN_3902; // @[sequencer-master.scala 168:32]
  wire  _GEN_5047 = _T_1442 ? _GEN_5039 : _GEN_3903; // @[sequencer-master.scala 168:32]
  wire  _GEN_5048 = _T_1442 ? _GEN_5040 : _GEN_3904; // @[sequencer-master.scala 168:32]
  wire  _GEN_5049 = _T_1442 ? _GEN_5041 : _GEN_3905; // @[sequencer-master.scala 168:32]
  wire  _GEN_5050 = _T_1442 ? _GEN_5042 : _GEN_3906; // @[sequencer-master.scala 168:32]
  wire  _GEN_5051 = _T_1442 ? _GEN_5043 : _GEN_3907; // @[sequencer-master.scala 168:32]
  wire  _GEN_5052 = _GEN_32729 | _GEN_3924; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5053 = _GEN_32730 | _GEN_3925; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5054 = _GEN_32731 | _GEN_3926; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5055 = _GEN_32732 | _GEN_3927; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5056 = _GEN_32733 | _GEN_3928; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5057 = _GEN_32734 | _GEN_3929; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5058 = _GEN_32735 | _GEN_3930; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5059 = _GEN_32736 | _GEN_3931; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5060 = _T_1464 ? _GEN_5052 : _GEN_3924; // @[sequencer-master.scala 168:32]
  wire  _GEN_5061 = _T_1464 ? _GEN_5053 : _GEN_3925; // @[sequencer-master.scala 168:32]
  wire  _GEN_5062 = _T_1464 ? _GEN_5054 : _GEN_3926; // @[sequencer-master.scala 168:32]
  wire  _GEN_5063 = _T_1464 ? _GEN_5055 : _GEN_3927; // @[sequencer-master.scala 168:32]
  wire  _GEN_5064 = _T_1464 ? _GEN_5056 : _GEN_3928; // @[sequencer-master.scala 168:32]
  wire  _GEN_5065 = _T_1464 ? _GEN_5057 : _GEN_3929; // @[sequencer-master.scala 168:32]
  wire  _GEN_5066 = _T_1464 ? _GEN_5058 : _GEN_3930; // @[sequencer-master.scala 168:32]
  wire  _GEN_5067 = _T_1464 ? _GEN_5059 : _GEN_3931; // @[sequencer-master.scala 168:32]
  wire  _GEN_5068 = _GEN_32729 | _GEN_3948; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5069 = _GEN_32730 | _GEN_3949; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5070 = _GEN_32731 | _GEN_3950; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5071 = _GEN_32732 | _GEN_3951; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5072 = _GEN_32733 | _GEN_3952; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5073 = _GEN_32734 | _GEN_3953; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5074 = _GEN_32735 | _GEN_3954; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5075 = _GEN_32736 | _GEN_3955; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5076 = _T_1486 ? _GEN_5068 : _GEN_3948; // @[sequencer-master.scala 168:32]
  wire  _GEN_5077 = _T_1486 ? _GEN_5069 : _GEN_3949; // @[sequencer-master.scala 168:32]
  wire  _GEN_5078 = _T_1486 ? _GEN_5070 : _GEN_3950; // @[sequencer-master.scala 168:32]
  wire  _GEN_5079 = _T_1486 ? _GEN_5071 : _GEN_3951; // @[sequencer-master.scala 168:32]
  wire  _GEN_5080 = _T_1486 ? _GEN_5072 : _GEN_3952; // @[sequencer-master.scala 168:32]
  wire  _GEN_5081 = _T_1486 ? _GEN_5073 : _GEN_3953; // @[sequencer-master.scala 168:32]
  wire  _GEN_5082 = _T_1486 ? _GEN_5074 : _GEN_3954; // @[sequencer-master.scala 168:32]
  wire  _GEN_5083 = _T_1486 ? _GEN_5075 : _GEN_3955; // @[sequencer-master.scala 168:32]
  wire  _GEN_5084 = _GEN_32729 | _GEN_3972; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5085 = _GEN_32730 | _GEN_3973; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5086 = _GEN_32731 | _GEN_3974; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5087 = _GEN_32732 | _GEN_3975; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5088 = _GEN_32733 | _GEN_3976; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5089 = _GEN_32734 | _GEN_3977; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5090 = _GEN_32735 | _GEN_3978; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5091 = _GEN_32736 | _GEN_3979; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5092 = _T_1508 ? _GEN_5084 : _GEN_3972; // @[sequencer-master.scala 168:32]
  wire  _GEN_5093 = _T_1508 ? _GEN_5085 : _GEN_3973; // @[sequencer-master.scala 168:32]
  wire  _GEN_5094 = _T_1508 ? _GEN_5086 : _GEN_3974; // @[sequencer-master.scala 168:32]
  wire  _GEN_5095 = _T_1508 ? _GEN_5087 : _GEN_3975; // @[sequencer-master.scala 168:32]
  wire  _GEN_5096 = _T_1508 ? _GEN_5088 : _GEN_3976; // @[sequencer-master.scala 168:32]
  wire  _GEN_5097 = _T_1508 ? _GEN_5089 : _GEN_3977; // @[sequencer-master.scala 168:32]
  wire  _GEN_5098 = _T_1508 ? _GEN_5090 : _GEN_3978; // @[sequencer-master.scala 168:32]
  wire  _GEN_5099 = _T_1508 ? _GEN_5091 : _GEN_3979; // @[sequencer-master.scala 168:32]
  wire  _GEN_5100 = _GEN_32729 | _GEN_3996; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5101 = _GEN_32730 | _GEN_3997; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5102 = _GEN_32731 | _GEN_3998; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5103 = _GEN_32732 | _GEN_3999; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5104 = _GEN_32733 | _GEN_4000; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5105 = _GEN_32734 | _GEN_4001; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5106 = _GEN_32735 | _GEN_4002; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5107 = _GEN_32736 | _GEN_4003; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5108 = _T_1530 ? _GEN_5100 : _GEN_3996; // @[sequencer-master.scala 168:32]
  wire  _GEN_5109 = _T_1530 ? _GEN_5101 : _GEN_3997; // @[sequencer-master.scala 168:32]
  wire  _GEN_5110 = _T_1530 ? _GEN_5102 : _GEN_3998; // @[sequencer-master.scala 168:32]
  wire  _GEN_5111 = _T_1530 ? _GEN_5103 : _GEN_3999; // @[sequencer-master.scala 168:32]
  wire  _GEN_5112 = _T_1530 ? _GEN_5104 : _GEN_4000; // @[sequencer-master.scala 168:32]
  wire  _GEN_5113 = _T_1530 ? _GEN_5105 : _GEN_4001; // @[sequencer-master.scala 168:32]
  wire  _GEN_5114 = _T_1530 ? _GEN_5106 : _GEN_4002; // @[sequencer-master.scala 168:32]
  wire  _GEN_5115 = _T_1530 ? _GEN_5107 : _GEN_4003; // @[sequencer-master.scala 168:32]
  wire  _GEN_5116 = _GEN_32729 | _GEN_4020; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5117 = _GEN_32730 | _GEN_4021; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5118 = _GEN_32731 | _GEN_4022; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5119 = _GEN_32732 | _GEN_4023; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5120 = _GEN_32733 | _GEN_4024; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5121 = _GEN_32734 | _GEN_4025; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5122 = _GEN_32735 | _GEN_4026; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5123 = _GEN_32736 | _GEN_4027; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5124 = _T_1552 ? _GEN_5116 : _GEN_4020; // @[sequencer-master.scala 168:32]
  wire  _GEN_5125 = _T_1552 ? _GEN_5117 : _GEN_4021; // @[sequencer-master.scala 168:32]
  wire  _GEN_5126 = _T_1552 ? _GEN_5118 : _GEN_4022; // @[sequencer-master.scala 168:32]
  wire  _GEN_5127 = _T_1552 ? _GEN_5119 : _GEN_4023; // @[sequencer-master.scala 168:32]
  wire  _GEN_5128 = _T_1552 ? _GEN_5120 : _GEN_4024; // @[sequencer-master.scala 168:32]
  wire  _GEN_5129 = _T_1552 ? _GEN_5121 : _GEN_4025; // @[sequencer-master.scala 168:32]
  wire  _GEN_5130 = _T_1552 ? _GEN_5122 : _GEN_4026; // @[sequencer-master.scala 168:32]
  wire  _GEN_5131 = _T_1552 ? _GEN_5123 : _GEN_4027; // @[sequencer-master.scala 168:32]
  wire  _GEN_5132 = _GEN_32729 | _GEN_4044; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5133 = _GEN_32730 | _GEN_4045; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5134 = _GEN_32731 | _GEN_4046; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5135 = _GEN_32732 | _GEN_4047; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5136 = _GEN_32733 | _GEN_4048; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5137 = _GEN_32734 | _GEN_4049; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5138 = _GEN_32735 | _GEN_4050; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5139 = _GEN_32736 | _GEN_4051; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5140 = _T_1574 ? _GEN_5132 : _GEN_4044; // @[sequencer-master.scala 168:32]
  wire  _GEN_5141 = _T_1574 ? _GEN_5133 : _GEN_4045; // @[sequencer-master.scala 168:32]
  wire  _GEN_5142 = _T_1574 ? _GEN_5134 : _GEN_4046; // @[sequencer-master.scala 168:32]
  wire  _GEN_5143 = _T_1574 ? _GEN_5135 : _GEN_4047; // @[sequencer-master.scala 168:32]
  wire  _GEN_5144 = _T_1574 ? _GEN_5136 : _GEN_4048; // @[sequencer-master.scala 168:32]
  wire  _GEN_5145 = _T_1574 ? _GEN_5137 : _GEN_4049; // @[sequencer-master.scala 168:32]
  wire  _GEN_5146 = _T_1574 ? _GEN_5138 : _GEN_4050; // @[sequencer-master.scala 168:32]
  wire  _GEN_5147 = _T_1574 ? _GEN_5139 : _GEN_4051; // @[sequencer-master.scala 168:32]
  wire  _GEN_5148 = _GEN_32729 | _GEN_4068; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5149 = _GEN_32730 | _GEN_4069; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5150 = _GEN_32731 | _GEN_4070; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5151 = _GEN_32732 | _GEN_4071; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5152 = _GEN_32733 | _GEN_4072; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5153 = _GEN_32734 | _GEN_4073; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5154 = _GEN_32735 | _GEN_4074; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5155 = _GEN_32736 | _GEN_4075; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_5156 = _T_1596 ? _GEN_5148 : _GEN_4068; // @[sequencer-master.scala 168:32]
  wire  _GEN_5157 = _T_1596 ? _GEN_5149 : _GEN_4069; // @[sequencer-master.scala 168:32]
  wire  _GEN_5158 = _T_1596 ? _GEN_5150 : _GEN_4070; // @[sequencer-master.scala 168:32]
  wire  _GEN_5159 = _T_1596 ? _GEN_5151 : _GEN_4071; // @[sequencer-master.scala 168:32]
  wire  _GEN_5160 = _T_1596 ? _GEN_5152 : _GEN_4072; // @[sequencer-master.scala 168:32]
  wire  _GEN_5161 = _T_1596 ? _GEN_5153 : _GEN_4073; // @[sequencer-master.scala 168:32]
  wire  _GEN_5162 = _T_1596 ? _GEN_5154 : _GEN_4074; // @[sequencer-master.scala 168:32]
  wire  _GEN_5163 = _T_1596 ? _GEN_5155 : _GEN_4075; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_5164 = 3'h0 == tail ? _T_1615[1:0] : _GEN_3794; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5165 = 3'h1 == tail ? _T_1615[1:0] : _GEN_3795; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5166 = 3'h2 == tail ? _T_1615[1:0] : _GEN_3796; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5167 = 3'h3 == tail ? _T_1615[1:0] : _GEN_3797; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5168 = 3'h4 == tail ? _T_1615[1:0] : _GEN_3798; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5169 = 3'h5 == tail ? _T_1615[1:0] : _GEN_3799; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5170 = 3'h6 == tail ? _T_1615[1:0] : _GEN_3800; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_5171 = 3'h7 == tail ? _T_1615[1:0] : _GEN_3801; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_5172 = 3'h0 == tail ? 4'h0 : _GEN_3802; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5173 = 3'h1 == tail ? 4'h0 : _GEN_3803; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5174 = 3'h2 == tail ? 4'h0 : _GEN_3804; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5175 = 3'h3 == tail ? 4'h0 : _GEN_3805; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5176 = 3'h4 == tail ? 4'h0 : _GEN_3806; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5177 = 3'h5 == tail ? 4'h0 : _GEN_3807; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5178 = 3'h6 == tail ? 4'h0 : _GEN_3808; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_5179 = 3'h7 == tail ? 4'h0 : _GEN_3809; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_5180 = 3'h0 == tail ? 3'h0 : _GEN_3810; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5181 = 3'h1 == tail ? 3'h0 : _GEN_3811; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5182 = 3'h2 == tail ? 3'h0 : _GEN_3812; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5183 = 3'h3 == tail ? 3'h0 : _GEN_3813; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5184 = 3'h4 == tail ? 3'h0 : _GEN_3814; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5185 = 3'h5 == tail ? 3'h0 : _GEN_3815; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5186 = 3'h6 == tail ? 3'h0 : _GEN_3816; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_5187 = 3'h7 == tail ? 3'h0 : _GEN_3817; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [3:0] _T_1880 = _T_1789[3:0] + 4'h4; // @[sequencer-master.scala 247:56]
  wire [3:0] _GEN_5188 = 3'h0 == tail ? _T_1880 : _GEN_5172; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5189 = 3'h1 == tail ? _T_1880 : _GEN_5173; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5190 = 3'h2 == tail ? _T_1880 : _GEN_5174; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5191 = 3'h3 == tail ? _T_1880 : _GEN_5175; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5192 = 3'h4 == tail ? _T_1880 : _GEN_5176; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5193 = 3'h5 == tail ? _T_1880 : _GEN_5177; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5194 = 3'h6 == tail ? _T_1880 : _GEN_5178; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5195 = 3'h7 == tail ? _T_1880 : _GEN_5179; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_5196 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5188 : _GEN_5172; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5197 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5189 : _GEN_5173; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5198 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5190 : _GEN_5174; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5199 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5191 : _GEN_5175; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5200 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5192 : _GEN_5176; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5201 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5193 : _GEN_5177; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5202 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5194 : _GEN_5178; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_5203 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_5195 : _GEN_5179; // @[sequencer-master.scala 235:47]
  wire [2:0] _GEN_5204 = 3'h0 == tail ? _T_1880[2:0] : _GEN_5180; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5205 = 3'h1 == tail ? _T_1880[2:0] : _GEN_5181; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5206 = 3'h2 == tail ? _T_1880[2:0] : _GEN_5182; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5207 = 3'h3 == tail ? _T_1880[2:0] : _GEN_5183; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5208 = 3'h4 == tail ? _T_1880[2:0] : _GEN_5184; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5209 = 3'h5 == tail ? _T_1880[2:0] : _GEN_5185; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5210 = 3'h6 == tail ? _T_1880[2:0] : _GEN_5186; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5211 = 3'h7 == tail ? _T_1880[2:0] : _GEN_5187; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_5212 = io_op_bits_base_vd_pred ? _GEN_5204 : _GEN_5180; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5213 = io_op_bits_base_vd_pred ? _GEN_5205 : _GEN_5181; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5214 = io_op_bits_base_vd_pred ? _GEN_5206 : _GEN_5182; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5215 = io_op_bits_base_vd_pred ? _GEN_5207 : _GEN_5183; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5216 = io_op_bits_base_vd_pred ? _GEN_5208 : _GEN_5184; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5217 = io_op_bits_base_vd_pred ? _GEN_5209 : _GEN_5185; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5218 = io_op_bits_base_vd_pred ? _GEN_5210 : _GEN_5186; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_5219 = io_op_bits_base_vd_pred ? _GEN_5211 : _GEN_5187; // @[sequencer-master.scala 236:45]
  wire  _GEN_5220 = io_op_bits_active_vimul ? _GEN_3820 : _GEN_3322; // @[sequencer-master.scala 642:40]
  wire  _GEN_5221 = io_op_bits_active_vimul ? _GEN_3821 : _GEN_3323; // @[sequencer-master.scala 642:40]
  wire  _GEN_5222 = io_op_bits_active_vimul ? _GEN_3822 : _GEN_3324; // @[sequencer-master.scala 642:40]
  wire  _GEN_5223 = io_op_bits_active_vimul ? _GEN_3823 : _GEN_3325; // @[sequencer-master.scala 642:40]
  wire  _GEN_5224 = io_op_bits_active_vimul ? _GEN_3824 : _GEN_3326; // @[sequencer-master.scala 642:40]
  wire  _GEN_5225 = io_op_bits_active_vimul ? _GEN_3825 : _GEN_3327; // @[sequencer-master.scala 642:40]
  wire  _GEN_5226 = io_op_bits_active_vimul ? _GEN_3826 : _GEN_3328; // @[sequencer-master.scala 642:40]
  wire  _GEN_5227 = io_op_bits_active_vimul ? _GEN_3827 : _GEN_3329; // @[sequencer-master.scala 642:40]
  wire  _GEN_5236 = io_op_bits_active_vimul ? _GEN_4156 : _GEN_3338; // @[sequencer-master.scala 642:40]
  wire  _GEN_5237 = io_op_bits_active_vimul ? _GEN_4157 : _GEN_3339; // @[sequencer-master.scala 642:40]
  wire  _GEN_5238 = io_op_bits_active_vimul ? _GEN_4158 : _GEN_3340; // @[sequencer-master.scala 642:40]
  wire  _GEN_5239 = io_op_bits_active_vimul ? _GEN_4159 : _GEN_3341; // @[sequencer-master.scala 642:40]
  wire  _GEN_5240 = io_op_bits_active_vimul ? _GEN_4160 : _GEN_3342; // @[sequencer-master.scala 642:40]
  wire  _GEN_5241 = io_op_bits_active_vimul ? _GEN_4161 : _GEN_3343; // @[sequencer-master.scala 642:40]
  wire  _GEN_5242 = io_op_bits_active_vimul ? _GEN_4162 : _GEN_3344; // @[sequencer-master.scala 642:40]
  wire  _GEN_5243 = io_op_bits_active_vimul ? _GEN_4163 : _GEN_3345; // @[sequencer-master.scala 642:40]
  wire  _GEN_5244 = io_op_bits_active_vimul ? _GEN_4388 : _GEN_3346; // @[sequencer-master.scala 642:40]
  wire  _GEN_5245 = io_op_bits_active_vimul ? _GEN_4389 : _GEN_3347; // @[sequencer-master.scala 642:40]
  wire  _GEN_5246 = io_op_bits_active_vimul ? _GEN_4390 : _GEN_3348; // @[sequencer-master.scala 642:40]
  wire  _GEN_5247 = io_op_bits_active_vimul ? _GEN_4391 : _GEN_3349; // @[sequencer-master.scala 642:40]
  wire  _GEN_5248 = io_op_bits_active_vimul ? _GEN_4392 : _GEN_3350; // @[sequencer-master.scala 642:40]
  wire  _GEN_5249 = io_op_bits_active_vimul ? _GEN_4393 : _GEN_3351; // @[sequencer-master.scala 642:40]
  wire  _GEN_5250 = io_op_bits_active_vimul ? _GEN_4394 : _GEN_3352; // @[sequencer-master.scala 642:40]
  wire  _GEN_5251 = io_op_bits_active_vimul ? _GEN_4395 : _GEN_3353; // @[sequencer-master.scala 642:40]
  wire  _GEN_5252 = io_op_bits_active_vimul ? _GEN_4636 : _GEN_3354; // @[sequencer-master.scala 642:40]
  wire  _GEN_5253 = io_op_bits_active_vimul ? _GEN_4637 : _GEN_3355; // @[sequencer-master.scala 642:40]
  wire  _GEN_5254 = io_op_bits_active_vimul ? _GEN_4638 : _GEN_3356; // @[sequencer-master.scala 642:40]
  wire  _GEN_5255 = io_op_bits_active_vimul ? _GEN_4639 : _GEN_3357; // @[sequencer-master.scala 642:40]
  wire  _GEN_5256 = io_op_bits_active_vimul ? _GEN_4640 : _GEN_3358; // @[sequencer-master.scala 642:40]
  wire  _GEN_5257 = io_op_bits_active_vimul ? _GEN_4641 : _GEN_3359; // @[sequencer-master.scala 642:40]
  wire  _GEN_5258 = io_op_bits_active_vimul ? _GEN_4642 : _GEN_3360; // @[sequencer-master.scala 642:40]
  wire  _GEN_5259 = io_op_bits_active_vimul ? _GEN_4643 : _GEN_3361; // @[sequencer-master.scala 642:40]
  wire  _GEN_5260 = io_op_bits_active_vimul ? _GEN_3860 : _GEN_3362; // @[sequencer-master.scala 642:40]
  wire  _GEN_5261 = io_op_bits_active_vimul ? _GEN_3861 : _GEN_3363; // @[sequencer-master.scala 642:40]
  wire  _GEN_5262 = io_op_bits_active_vimul ? _GEN_3862 : _GEN_3364; // @[sequencer-master.scala 642:40]
  wire  _GEN_5263 = io_op_bits_active_vimul ? _GEN_3863 : _GEN_3365; // @[sequencer-master.scala 642:40]
  wire  _GEN_5264 = io_op_bits_active_vimul ? _GEN_3864 : _GEN_3366; // @[sequencer-master.scala 642:40]
  wire  _GEN_5265 = io_op_bits_active_vimul ? _GEN_3865 : _GEN_3367; // @[sequencer-master.scala 642:40]
  wire  _GEN_5266 = io_op_bits_active_vimul ? _GEN_3866 : _GEN_3368; // @[sequencer-master.scala 642:40]
  wire  _GEN_5267 = io_op_bits_active_vimul ? _GEN_3867 : _GEN_3369; // @[sequencer-master.scala 642:40]
  wire  _GEN_5268 = io_op_bits_active_vimul ? _GEN_4868 : _GEN_3370; // @[sequencer-master.scala 642:40]
  wire  _GEN_5269 = io_op_bits_active_vimul ? _GEN_4869 : _GEN_3371; // @[sequencer-master.scala 642:40]
  wire  _GEN_5270 = io_op_bits_active_vimul ? _GEN_4870 : _GEN_3372; // @[sequencer-master.scala 642:40]
  wire  _GEN_5271 = io_op_bits_active_vimul ? _GEN_4871 : _GEN_3373; // @[sequencer-master.scala 642:40]
  wire  _GEN_5272 = io_op_bits_active_vimul ? _GEN_4872 : _GEN_3374; // @[sequencer-master.scala 642:40]
  wire  _GEN_5273 = io_op_bits_active_vimul ? _GEN_4873 : _GEN_3375; // @[sequencer-master.scala 642:40]
  wire  _GEN_5274 = io_op_bits_active_vimul ? _GEN_4874 : _GEN_3376; // @[sequencer-master.scala 642:40]
  wire  _GEN_5275 = io_op_bits_active_vimul ? _GEN_4875 : _GEN_3377; // @[sequencer-master.scala 642:40]
  wire  _GEN_5276 = io_op_bits_active_vimul ? _GEN_3876 : _GEN_3378; // @[sequencer-master.scala 642:40]
  wire  _GEN_5277 = io_op_bits_active_vimul ? _GEN_3877 : _GEN_3379; // @[sequencer-master.scala 642:40]
  wire  _GEN_5278 = io_op_bits_active_vimul ? _GEN_3878 : _GEN_3380; // @[sequencer-master.scala 642:40]
  wire  _GEN_5279 = io_op_bits_active_vimul ? _GEN_3879 : _GEN_3381; // @[sequencer-master.scala 642:40]
  wire  _GEN_5280 = io_op_bits_active_vimul ? _GEN_3880 : _GEN_3382; // @[sequencer-master.scala 642:40]
  wire  _GEN_5281 = io_op_bits_active_vimul ? _GEN_3881 : _GEN_3383; // @[sequencer-master.scala 642:40]
  wire  _GEN_5282 = io_op_bits_active_vimul ? _GEN_3882 : _GEN_3384; // @[sequencer-master.scala 642:40]
  wire  _GEN_5283 = io_op_bits_active_vimul ? _GEN_3883 : _GEN_3385; // @[sequencer-master.scala 642:40]
  wire  _GEN_5284 = io_op_bits_active_vimul ? _GEN_4692 : _GEN_3386; // @[sequencer-master.scala 642:40]
  wire  _GEN_5285 = io_op_bits_active_vimul ? _GEN_4693 : _GEN_3387; // @[sequencer-master.scala 642:40]
  wire  _GEN_5286 = io_op_bits_active_vimul ? _GEN_4694 : _GEN_3388; // @[sequencer-master.scala 642:40]
  wire  _GEN_5287 = io_op_bits_active_vimul ? _GEN_4695 : _GEN_3389; // @[sequencer-master.scala 642:40]
  wire  _GEN_5288 = io_op_bits_active_vimul ? _GEN_4696 : _GEN_3390; // @[sequencer-master.scala 642:40]
  wire  _GEN_5289 = io_op_bits_active_vimul ? _GEN_4697 : _GEN_3391; // @[sequencer-master.scala 642:40]
  wire  _GEN_5290 = io_op_bits_active_vimul ? _GEN_4698 : _GEN_3392; // @[sequencer-master.scala 642:40]
  wire  _GEN_5291 = io_op_bits_active_vimul ? _GEN_4699 : _GEN_3393; // @[sequencer-master.scala 642:40]
  wire  _GEN_5292 = io_op_bits_active_vimul ? _GEN_4916 : _GEN_3394; // @[sequencer-master.scala 642:40]
  wire  _GEN_5293 = io_op_bits_active_vimul ? _GEN_4917 : _GEN_3395; // @[sequencer-master.scala 642:40]
  wire  _GEN_5294 = io_op_bits_active_vimul ? _GEN_4918 : _GEN_3396; // @[sequencer-master.scala 642:40]
  wire  _GEN_5295 = io_op_bits_active_vimul ? _GEN_4919 : _GEN_3397; // @[sequencer-master.scala 642:40]
  wire  _GEN_5296 = io_op_bits_active_vimul ? _GEN_4920 : _GEN_3398; // @[sequencer-master.scala 642:40]
  wire  _GEN_5297 = io_op_bits_active_vimul ? _GEN_4921 : _GEN_3399; // @[sequencer-master.scala 642:40]
  wire  _GEN_5298 = io_op_bits_active_vimul ? _GEN_4922 : _GEN_3400; // @[sequencer-master.scala 642:40]
  wire  _GEN_5299 = io_op_bits_active_vimul ? _GEN_4923 : _GEN_3401; // @[sequencer-master.scala 642:40]
  wire  _GEN_5300 = io_op_bits_active_vimul ? _GEN_5044 : _GEN_3402; // @[sequencer-master.scala 642:40]
  wire  _GEN_5301 = io_op_bits_active_vimul ? _GEN_5045 : _GEN_3403; // @[sequencer-master.scala 642:40]
  wire  _GEN_5302 = io_op_bits_active_vimul ? _GEN_5046 : _GEN_3404; // @[sequencer-master.scala 642:40]
  wire  _GEN_5303 = io_op_bits_active_vimul ? _GEN_5047 : _GEN_3405; // @[sequencer-master.scala 642:40]
  wire  _GEN_5304 = io_op_bits_active_vimul ? _GEN_5048 : _GEN_3406; // @[sequencer-master.scala 642:40]
  wire  _GEN_5305 = io_op_bits_active_vimul ? _GEN_5049 : _GEN_3407; // @[sequencer-master.scala 642:40]
  wire  _GEN_5306 = io_op_bits_active_vimul ? _GEN_5050 : _GEN_3408; // @[sequencer-master.scala 642:40]
  wire  _GEN_5307 = io_op_bits_active_vimul ? _GEN_5051 : _GEN_3409; // @[sequencer-master.scala 642:40]
  wire  _GEN_5308 = io_op_bits_active_vimul ? _GEN_4708 : _GEN_3410; // @[sequencer-master.scala 642:40]
  wire  _GEN_5309 = io_op_bits_active_vimul ? _GEN_4709 : _GEN_3411; // @[sequencer-master.scala 642:40]
  wire  _GEN_5310 = io_op_bits_active_vimul ? _GEN_4710 : _GEN_3412; // @[sequencer-master.scala 642:40]
  wire  _GEN_5311 = io_op_bits_active_vimul ? _GEN_4711 : _GEN_3413; // @[sequencer-master.scala 642:40]
  wire  _GEN_5312 = io_op_bits_active_vimul ? _GEN_4712 : _GEN_3414; // @[sequencer-master.scala 642:40]
  wire  _GEN_5313 = io_op_bits_active_vimul ? _GEN_4713 : _GEN_3415; // @[sequencer-master.scala 642:40]
  wire  _GEN_5314 = io_op_bits_active_vimul ? _GEN_4714 : _GEN_3416; // @[sequencer-master.scala 642:40]
  wire  _GEN_5315 = io_op_bits_active_vimul ? _GEN_4715 : _GEN_3417; // @[sequencer-master.scala 642:40]
  wire  _GEN_5316 = io_op_bits_active_vimul ? _GEN_4932 : _GEN_3418; // @[sequencer-master.scala 642:40]
  wire  _GEN_5317 = io_op_bits_active_vimul ? _GEN_4933 : _GEN_3419; // @[sequencer-master.scala 642:40]
  wire  _GEN_5318 = io_op_bits_active_vimul ? _GEN_4934 : _GEN_3420; // @[sequencer-master.scala 642:40]
  wire  _GEN_5319 = io_op_bits_active_vimul ? _GEN_4935 : _GEN_3421; // @[sequencer-master.scala 642:40]
  wire  _GEN_5320 = io_op_bits_active_vimul ? _GEN_4936 : _GEN_3422; // @[sequencer-master.scala 642:40]
  wire  _GEN_5321 = io_op_bits_active_vimul ? _GEN_4937 : _GEN_3423; // @[sequencer-master.scala 642:40]
  wire  _GEN_5322 = io_op_bits_active_vimul ? _GEN_4938 : _GEN_3424; // @[sequencer-master.scala 642:40]
  wire  _GEN_5323 = io_op_bits_active_vimul ? _GEN_4939 : _GEN_3425; // @[sequencer-master.scala 642:40]
  wire  _GEN_5324 = io_op_bits_active_vimul ? _GEN_5060 : _GEN_3426; // @[sequencer-master.scala 642:40]
  wire  _GEN_5325 = io_op_bits_active_vimul ? _GEN_5061 : _GEN_3427; // @[sequencer-master.scala 642:40]
  wire  _GEN_5326 = io_op_bits_active_vimul ? _GEN_5062 : _GEN_3428; // @[sequencer-master.scala 642:40]
  wire  _GEN_5327 = io_op_bits_active_vimul ? _GEN_5063 : _GEN_3429; // @[sequencer-master.scala 642:40]
  wire  _GEN_5328 = io_op_bits_active_vimul ? _GEN_5064 : _GEN_3430; // @[sequencer-master.scala 642:40]
  wire  _GEN_5329 = io_op_bits_active_vimul ? _GEN_5065 : _GEN_3431; // @[sequencer-master.scala 642:40]
  wire  _GEN_5330 = io_op_bits_active_vimul ? _GEN_5066 : _GEN_3432; // @[sequencer-master.scala 642:40]
  wire  _GEN_5331 = io_op_bits_active_vimul ? _GEN_5067 : _GEN_3433; // @[sequencer-master.scala 642:40]
  wire  _GEN_5332 = io_op_bits_active_vimul ? _GEN_4724 : _GEN_3434; // @[sequencer-master.scala 642:40]
  wire  _GEN_5333 = io_op_bits_active_vimul ? _GEN_4725 : _GEN_3435; // @[sequencer-master.scala 642:40]
  wire  _GEN_5334 = io_op_bits_active_vimul ? _GEN_4726 : _GEN_3436; // @[sequencer-master.scala 642:40]
  wire  _GEN_5335 = io_op_bits_active_vimul ? _GEN_4727 : _GEN_3437; // @[sequencer-master.scala 642:40]
  wire  _GEN_5336 = io_op_bits_active_vimul ? _GEN_4728 : _GEN_3438; // @[sequencer-master.scala 642:40]
  wire  _GEN_5337 = io_op_bits_active_vimul ? _GEN_4729 : _GEN_3439; // @[sequencer-master.scala 642:40]
  wire  _GEN_5338 = io_op_bits_active_vimul ? _GEN_4730 : _GEN_3440; // @[sequencer-master.scala 642:40]
  wire  _GEN_5339 = io_op_bits_active_vimul ? _GEN_4731 : _GEN_3441; // @[sequencer-master.scala 642:40]
  wire  _GEN_5340 = io_op_bits_active_vimul ? _GEN_4948 : _GEN_3442; // @[sequencer-master.scala 642:40]
  wire  _GEN_5341 = io_op_bits_active_vimul ? _GEN_4949 : _GEN_3443; // @[sequencer-master.scala 642:40]
  wire  _GEN_5342 = io_op_bits_active_vimul ? _GEN_4950 : _GEN_3444; // @[sequencer-master.scala 642:40]
  wire  _GEN_5343 = io_op_bits_active_vimul ? _GEN_4951 : _GEN_3445; // @[sequencer-master.scala 642:40]
  wire  _GEN_5344 = io_op_bits_active_vimul ? _GEN_4952 : _GEN_3446; // @[sequencer-master.scala 642:40]
  wire  _GEN_5345 = io_op_bits_active_vimul ? _GEN_4953 : _GEN_3447; // @[sequencer-master.scala 642:40]
  wire  _GEN_5346 = io_op_bits_active_vimul ? _GEN_4954 : _GEN_3448; // @[sequencer-master.scala 642:40]
  wire  _GEN_5347 = io_op_bits_active_vimul ? _GEN_4955 : _GEN_3449; // @[sequencer-master.scala 642:40]
  wire  _GEN_5348 = io_op_bits_active_vimul ? _GEN_5076 : _GEN_3450; // @[sequencer-master.scala 642:40]
  wire  _GEN_5349 = io_op_bits_active_vimul ? _GEN_5077 : _GEN_3451; // @[sequencer-master.scala 642:40]
  wire  _GEN_5350 = io_op_bits_active_vimul ? _GEN_5078 : _GEN_3452; // @[sequencer-master.scala 642:40]
  wire  _GEN_5351 = io_op_bits_active_vimul ? _GEN_5079 : _GEN_3453; // @[sequencer-master.scala 642:40]
  wire  _GEN_5352 = io_op_bits_active_vimul ? _GEN_5080 : _GEN_3454; // @[sequencer-master.scala 642:40]
  wire  _GEN_5353 = io_op_bits_active_vimul ? _GEN_5081 : _GEN_3455; // @[sequencer-master.scala 642:40]
  wire  _GEN_5354 = io_op_bits_active_vimul ? _GEN_5082 : _GEN_3456; // @[sequencer-master.scala 642:40]
  wire  _GEN_5355 = io_op_bits_active_vimul ? _GEN_5083 : _GEN_3457; // @[sequencer-master.scala 642:40]
  wire  _GEN_5356 = io_op_bits_active_vimul ? _GEN_4740 : _GEN_3458; // @[sequencer-master.scala 642:40]
  wire  _GEN_5357 = io_op_bits_active_vimul ? _GEN_4741 : _GEN_3459; // @[sequencer-master.scala 642:40]
  wire  _GEN_5358 = io_op_bits_active_vimul ? _GEN_4742 : _GEN_3460; // @[sequencer-master.scala 642:40]
  wire  _GEN_5359 = io_op_bits_active_vimul ? _GEN_4743 : _GEN_3461; // @[sequencer-master.scala 642:40]
  wire  _GEN_5360 = io_op_bits_active_vimul ? _GEN_4744 : _GEN_3462; // @[sequencer-master.scala 642:40]
  wire  _GEN_5361 = io_op_bits_active_vimul ? _GEN_4745 : _GEN_3463; // @[sequencer-master.scala 642:40]
  wire  _GEN_5362 = io_op_bits_active_vimul ? _GEN_4746 : _GEN_3464; // @[sequencer-master.scala 642:40]
  wire  _GEN_5363 = io_op_bits_active_vimul ? _GEN_4747 : _GEN_3465; // @[sequencer-master.scala 642:40]
  wire  _GEN_5364 = io_op_bits_active_vimul ? _GEN_4964 : _GEN_3466; // @[sequencer-master.scala 642:40]
  wire  _GEN_5365 = io_op_bits_active_vimul ? _GEN_4965 : _GEN_3467; // @[sequencer-master.scala 642:40]
  wire  _GEN_5366 = io_op_bits_active_vimul ? _GEN_4966 : _GEN_3468; // @[sequencer-master.scala 642:40]
  wire  _GEN_5367 = io_op_bits_active_vimul ? _GEN_4967 : _GEN_3469; // @[sequencer-master.scala 642:40]
  wire  _GEN_5368 = io_op_bits_active_vimul ? _GEN_4968 : _GEN_3470; // @[sequencer-master.scala 642:40]
  wire  _GEN_5369 = io_op_bits_active_vimul ? _GEN_4969 : _GEN_3471; // @[sequencer-master.scala 642:40]
  wire  _GEN_5370 = io_op_bits_active_vimul ? _GEN_4970 : _GEN_3472; // @[sequencer-master.scala 642:40]
  wire  _GEN_5371 = io_op_bits_active_vimul ? _GEN_4971 : _GEN_3473; // @[sequencer-master.scala 642:40]
  wire  _GEN_5372 = io_op_bits_active_vimul ? _GEN_5092 : _GEN_3474; // @[sequencer-master.scala 642:40]
  wire  _GEN_5373 = io_op_bits_active_vimul ? _GEN_5093 : _GEN_3475; // @[sequencer-master.scala 642:40]
  wire  _GEN_5374 = io_op_bits_active_vimul ? _GEN_5094 : _GEN_3476; // @[sequencer-master.scala 642:40]
  wire  _GEN_5375 = io_op_bits_active_vimul ? _GEN_5095 : _GEN_3477; // @[sequencer-master.scala 642:40]
  wire  _GEN_5376 = io_op_bits_active_vimul ? _GEN_5096 : _GEN_3478; // @[sequencer-master.scala 642:40]
  wire  _GEN_5377 = io_op_bits_active_vimul ? _GEN_5097 : _GEN_3479; // @[sequencer-master.scala 642:40]
  wire  _GEN_5378 = io_op_bits_active_vimul ? _GEN_5098 : _GEN_3480; // @[sequencer-master.scala 642:40]
  wire  _GEN_5379 = io_op_bits_active_vimul ? _GEN_5099 : _GEN_3481; // @[sequencer-master.scala 642:40]
  wire  _GEN_5380 = io_op_bits_active_vimul ? _GEN_4756 : _GEN_3482; // @[sequencer-master.scala 642:40]
  wire  _GEN_5381 = io_op_bits_active_vimul ? _GEN_4757 : _GEN_3483; // @[sequencer-master.scala 642:40]
  wire  _GEN_5382 = io_op_bits_active_vimul ? _GEN_4758 : _GEN_3484; // @[sequencer-master.scala 642:40]
  wire  _GEN_5383 = io_op_bits_active_vimul ? _GEN_4759 : _GEN_3485; // @[sequencer-master.scala 642:40]
  wire  _GEN_5384 = io_op_bits_active_vimul ? _GEN_4760 : _GEN_3486; // @[sequencer-master.scala 642:40]
  wire  _GEN_5385 = io_op_bits_active_vimul ? _GEN_4761 : _GEN_3487; // @[sequencer-master.scala 642:40]
  wire  _GEN_5386 = io_op_bits_active_vimul ? _GEN_4762 : _GEN_3488; // @[sequencer-master.scala 642:40]
  wire  _GEN_5387 = io_op_bits_active_vimul ? _GEN_4763 : _GEN_3489; // @[sequencer-master.scala 642:40]
  wire  _GEN_5388 = io_op_bits_active_vimul ? _GEN_4980 : _GEN_3490; // @[sequencer-master.scala 642:40]
  wire  _GEN_5389 = io_op_bits_active_vimul ? _GEN_4981 : _GEN_3491; // @[sequencer-master.scala 642:40]
  wire  _GEN_5390 = io_op_bits_active_vimul ? _GEN_4982 : _GEN_3492; // @[sequencer-master.scala 642:40]
  wire  _GEN_5391 = io_op_bits_active_vimul ? _GEN_4983 : _GEN_3493; // @[sequencer-master.scala 642:40]
  wire  _GEN_5392 = io_op_bits_active_vimul ? _GEN_4984 : _GEN_3494; // @[sequencer-master.scala 642:40]
  wire  _GEN_5393 = io_op_bits_active_vimul ? _GEN_4985 : _GEN_3495; // @[sequencer-master.scala 642:40]
  wire  _GEN_5394 = io_op_bits_active_vimul ? _GEN_4986 : _GEN_3496; // @[sequencer-master.scala 642:40]
  wire  _GEN_5395 = io_op_bits_active_vimul ? _GEN_4987 : _GEN_3497; // @[sequencer-master.scala 642:40]
  wire  _GEN_5396 = io_op_bits_active_vimul ? _GEN_5108 : _GEN_3498; // @[sequencer-master.scala 642:40]
  wire  _GEN_5397 = io_op_bits_active_vimul ? _GEN_5109 : _GEN_3499; // @[sequencer-master.scala 642:40]
  wire  _GEN_5398 = io_op_bits_active_vimul ? _GEN_5110 : _GEN_3500; // @[sequencer-master.scala 642:40]
  wire  _GEN_5399 = io_op_bits_active_vimul ? _GEN_5111 : _GEN_3501; // @[sequencer-master.scala 642:40]
  wire  _GEN_5400 = io_op_bits_active_vimul ? _GEN_5112 : _GEN_3502; // @[sequencer-master.scala 642:40]
  wire  _GEN_5401 = io_op_bits_active_vimul ? _GEN_5113 : _GEN_3503; // @[sequencer-master.scala 642:40]
  wire  _GEN_5402 = io_op_bits_active_vimul ? _GEN_5114 : _GEN_3504; // @[sequencer-master.scala 642:40]
  wire  _GEN_5403 = io_op_bits_active_vimul ? _GEN_5115 : _GEN_3505; // @[sequencer-master.scala 642:40]
  wire  _GEN_5404 = io_op_bits_active_vimul ? _GEN_4772 : _GEN_3506; // @[sequencer-master.scala 642:40]
  wire  _GEN_5405 = io_op_bits_active_vimul ? _GEN_4773 : _GEN_3507; // @[sequencer-master.scala 642:40]
  wire  _GEN_5406 = io_op_bits_active_vimul ? _GEN_4774 : _GEN_3508; // @[sequencer-master.scala 642:40]
  wire  _GEN_5407 = io_op_bits_active_vimul ? _GEN_4775 : _GEN_3509; // @[sequencer-master.scala 642:40]
  wire  _GEN_5408 = io_op_bits_active_vimul ? _GEN_4776 : _GEN_3510; // @[sequencer-master.scala 642:40]
  wire  _GEN_5409 = io_op_bits_active_vimul ? _GEN_4777 : _GEN_3511; // @[sequencer-master.scala 642:40]
  wire  _GEN_5410 = io_op_bits_active_vimul ? _GEN_4778 : _GEN_3512; // @[sequencer-master.scala 642:40]
  wire  _GEN_5411 = io_op_bits_active_vimul ? _GEN_4779 : _GEN_3513; // @[sequencer-master.scala 642:40]
  wire  _GEN_5412 = io_op_bits_active_vimul ? _GEN_4996 : _GEN_3514; // @[sequencer-master.scala 642:40]
  wire  _GEN_5413 = io_op_bits_active_vimul ? _GEN_4997 : _GEN_3515; // @[sequencer-master.scala 642:40]
  wire  _GEN_5414 = io_op_bits_active_vimul ? _GEN_4998 : _GEN_3516; // @[sequencer-master.scala 642:40]
  wire  _GEN_5415 = io_op_bits_active_vimul ? _GEN_4999 : _GEN_3517; // @[sequencer-master.scala 642:40]
  wire  _GEN_5416 = io_op_bits_active_vimul ? _GEN_5000 : _GEN_3518; // @[sequencer-master.scala 642:40]
  wire  _GEN_5417 = io_op_bits_active_vimul ? _GEN_5001 : _GEN_3519; // @[sequencer-master.scala 642:40]
  wire  _GEN_5418 = io_op_bits_active_vimul ? _GEN_5002 : _GEN_3520; // @[sequencer-master.scala 642:40]
  wire  _GEN_5419 = io_op_bits_active_vimul ? _GEN_5003 : _GEN_3521; // @[sequencer-master.scala 642:40]
  wire  _GEN_5420 = io_op_bits_active_vimul ? _GEN_5124 : _GEN_3522; // @[sequencer-master.scala 642:40]
  wire  _GEN_5421 = io_op_bits_active_vimul ? _GEN_5125 : _GEN_3523; // @[sequencer-master.scala 642:40]
  wire  _GEN_5422 = io_op_bits_active_vimul ? _GEN_5126 : _GEN_3524; // @[sequencer-master.scala 642:40]
  wire  _GEN_5423 = io_op_bits_active_vimul ? _GEN_5127 : _GEN_3525; // @[sequencer-master.scala 642:40]
  wire  _GEN_5424 = io_op_bits_active_vimul ? _GEN_5128 : _GEN_3526; // @[sequencer-master.scala 642:40]
  wire  _GEN_5425 = io_op_bits_active_vimul ? _GEN_5129 : _GEN_3527; // @[sequencer-master.scala 642:40]
  wire  _GEN_5426 = io_op_bits_active_vimul ? _GEN_5130 : _GEN_3528; // @[sequencer-master.scala 642:40]
  wire  _GEN_5427 = io_op_bits_active_vimul ? _GEN_5131 : _GEN_3529; // @[sequencer-master.scala 642:40]
  wire  _GEN_5428 = io_op_bits_active_vimul ? _GEN_4788 : _GEN_3530; // @[sequencer-master.scala 642:40]
  wire  _GEN_5429 = io_op_bits_active_vimul ? _GEN_4789 : _GEN_3531; // @[sequencer-master.scala 642:40]
  wire  _GEN_5430 = io_op_bits_active_vimul ? _GEN_4790 : _GEN_3532; // @[sequencer-master.scala 642:40]
  wire  _GEN_5431 = io_op_bits_active_vimul ? _GEN_4791 : _GEN_3533; // @[sequencer-master.scala 642:40]
  wire  _GEN_5432 = io_op_bits_active_vimul ? _GEN_4792 : _GEN_3534; // @[sequencer-master.scala 642:40]
  wire  _GEN_5433 = io_op_bits_active_vimul ? _GEN_4793 : _GEN_3535; // @[sequencer-master.scala 642:40]
  wire  _GEN_5434 = io_op_bits_active_vimul ? _GEN_4794 : _GEN_3536; // @[sequencer-master.scala 642:40]
  wire  _GEN_5435 = io_op_bits_active_vimul ? _GEN_4795 : _GEN_3537; // @[sequencer-master.scala 642:40]
  wire  _GEN_5436 = io_op_bits_active_vimul ? _GEN_5012 : _GEN_3538; // @[sequencer-master.scala 642:40]
  wire  _GEN_5437 = io_op_bits_active_vimul ? _GEN_5013 : _GEN_3539; // @[sequencer-master.scala 642:40]
  wire  _GEN_5438 = io_op_bits_active_vimul ? _GEN_5014 : _GEN_3540; // @[sequencer-master.scala 642:40]
  wire  _GEN_5439 = io_op_bits_active_vimul ? _GEN_5015 : _GEN_3541; // @[sequencer-master.scala 642:40]
  wire  _GEN_5440 = io_op_bits_active_vimul ? _GEN_5016 : _GEN_3542; // @[sequencer-master.scala 642:40]
  wire  _GEN_5441 = io_op_bits_active_vimul ? _GEN_5017 : _GEN_3543; // @[sequencer-master.scala 642:40]
  wire  _GEN_5442 = io_op_bits_active_vimul ? _GEN_5018 : _GEN_3544; // @[sequencer-master.scala 642:40]
  wire  _GEN_5443 = io_op_bits_active_vimul ? _GEN_5019 : _GEN_3545; // @[sequencer-master.scala 642:40]
  wire  _GEN_5444 = io_op_bits_active_vimul ? _GEN_5140 : _GEN_3546; // @[sequencer-master.scala 642:40]
  wire  _GEN_5445 = io_op_bits_active_vimul ? _GEN_5141 : _GEN_3547; // @[sequencer-master.scala 642:40]
  wire  _GEN_5446 = io_op_bits_active_vimul ? _GEN_5142 : _GEN_3548; // @[sequencer-master.scala 642:40]
  wire  _GEN_5447 = io_op_bits_active_vimul ? _GEN_5143 : _GEN_3549; // @[sequencer-master.scala 642:40]
  wire  _GEN_5448 = io_op_bits_active_vimul ? _GEN_5144 : _GEN_3550; // @[sequencer-master.scala 642:40]
  wire  _GEN_5449 = io_op_bits_active_vimul ? _GEN_5145 : _GEN_3551; // @[sequencer-master.scala 642:40]
  wire  _GEN_5450 = io_op_bits_active_vimul ? _GEN_5146 : _GEN_3552; // @[sequencer-master.scala 642:40]
  wire  _GEN_5451 = io_op_bits_active_vimul ? _GEN_5147 : _GEN_3553; // @[sequencer-master.scala 642:40]
  wire  _GEN_5452 = io_op_bits_active_vimul ? _GEN_4804 : _GEN_3554; // @[sequencer-master.scala 642:40]
  wire  _GEN_5453 = io_op_bits_active_vimul ? _GEN_4805 : _GEN_3555; // @[sequencer-master.scala 642:40]
  wire  _GEN_5454 = io_op_bits_active_vimul ? _GEN_4806 : _GEN_3556; // @[sequencer-master.scala 642:40]
  wire  _GEN_5455 = io_op_bits_active_vimul ? _GEN_4807 : _GEN_3557; // @[sequencer-master.scala 642:40]
  wire  _GEN_5456 = io_op_bits_active_vimul ? _GEN_4808 : _GEN_3558; // @[sequencer-master.scala 642:40]
  wire  _GEN_5457 = io_op_bits_active_vimul ? _GEN_4809 : _GEN_3559; // @[sequencer-master.scala 642:40]
  wire  _GEN_5458 = io_op_bits_active_vimul ? _GEN_4810 : _GEN_3560; // @[sequencer-master.scala 642:40]
  wire  _GEN_5459 = io_op_bits_active_vimul ? _GEN_4811 : _GEN_3561; // @[sequencer-master.scala 642:40]
  wire  _GEN_5460 = io_op_bits_active_vimul ? _GEN_5028 : _GEN_3562; // @[sequencer-master.scala 642:40]
  wire  _GEN_5461 = io_op_bits_active_vimul ? _GEN_5029 : _GEN_3563; // @[sequencer-master.scala 642:40]
  wire  _GEN_5462 = io_op_bits_active_vimul ? _GEN_5030 : _GEN_3564; // @[sequencer-master.scala 642:40]
  wire  _GEN_5463 = io_op_bits_active_vimul ? _GEN_5031 : _GEN_3565; // @[sequencer-master.scala 642:40]
  wire  _GEN_5464 = io_op_bits_active_vimul ? _GEN_5032 : _GEN_3566; // @[sequencer-master.scala 642:40]
  wire  _GEN_5465 = io_op_bits_active_vimul ? _GEN_5033 : _GEN_3567; // @[sequencer-master.scala 642:40]
  wire  _GEN_5466 = io_op_bits_active_vimul ? _GEN_5034 : _GEN_3568; // @[sequencer-master.scala 642:40]
  wire  _GEN_5467 = io_op_bits_active_vimul ? _GEN_5035 : _GEN_3569; // @[sequencer-master.scala 642:40]
  wire  _GEN_5468 = io_op_bits_active_vimul ? _GEN_5156 : _GEN_3570; // @[sequencer-master.scala 642:40]
  wire  _GEN_5469 = io_op_bits_active_vimul ? _GEN_5157 : _GEN_3571; // @[sequencer-master.scala 642:40]
  wire  _GEN_5470 = io_op_bits_active_vimul ? _GEN_5158 : _GEN_3572; // @[sequencer-master.scala 642:40]
  wire  _GEN_5471 = io_op_bits_active_vimul ? _GEN_5159 : _GEN_3573; // @[sequencer-master.scala 642:40]
  wire  _GEN_5472 = io_op_bits_active_vimul ? _GEN_5160 : _GEN_3574; // @[sequencer-master.scala 642:40]
  wire  _GEN_5473 = io_op_bits_active_vimul ? _GEN_5161 : _GEN_3575; // @[sequencer-master.scala 642:40]
  wire  _GEN_5474 = io_op_bits_active_vimul ? _GEN_5162 : _GEN_3576; // @[sequencer-master.scala 642:40]
  wire  _GEN_5475 = io_op_bits_active_vimul ? _GEN_5163 : _GEN_3577; // @[sequencer-master.scala 642:40]
  wire  _GEN_5476 = io_op_bits_active_vimul ? _GEN_4076 : _GEN_3578; // @[sequencer-master.scala 642:40]
  wire  _GEN_5477 = io_op_bits_active_vimul ? _GEN_4077 : _GEN_3579; // @[sequencer-master.scala 642:40]
  wire  _GEN_5478 = io_op_bits_active_vimul ? _GEN_4078 : _GEN_3580; // @[sequencer-master.scala 642:40]
  wire  _GEN_5479 = io_op_bits_active_vimul ? _GEN_4079 : _GEN_3581; // @[sequencer-master.scala 642:40]
  wire  _GEN_5480 = io_op_bits_active_vimul ? _GEN_4080 : _GEN_3582; // @[sequencer-master.scala 642:40]
  wire  _GEN_5481 = io_op_bits_active_vimul ? _GEN_4081 : _GEN_3583; // @[sequencer-master.scala 642:40]
  wire  _GEN_5482 = io_op_bits_active_vimul ? _GEN_4082 : _GEN_3584; // @[sequencer-master.scala 642:40]
  wire  _GEN_5483 = io_op_bits_active_vimul ? _GEN_4083 : _GEN_3585; // @[sequencer-master.scala 642:40]
  wire  _GEN_5492 = io_op_bits_active_vimul ? _GEN_4092 : e_0_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5493 = io_op_bits_active_vimul ? _GEN_4093 : e_1_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5494 = io_op_bits_active_vimul ? _GEN_4094 : e_2_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5495 = io_op_bits_active_vimul ? _GEN_4095 : e_3_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5496 = io_op_bits_active_vimul ? _GEN_4096 : e_4_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5497 = io_op_bits_active_vimul ? _GEN_4097 : e_5_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5498 = io_op_bits_active_vimul ? _GEN_4098 : e_6_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire  _GEN_5499 = io_op_bits_active_vimul ? _GEN_4099 : e_7_active_vimu; // @[sequencer-master.scala 642:40 sequencer-master.scala 109:14]
  wire [9:0] _GEN_5500 = io_op_bits_active_vimul ? _GEN_4100 : _GEN_3602; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5501 = io_op_bits_active_vimul ? _GEN_4101 : _GEN_3603; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5502 = io_op_bits_active_vimul ? _GEN_4102 : _GEN_3604; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5503 = io_op_bits_active_vimul ? _GEN_4103 : _GEN_3605; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5504 = io_op_bits_active_vimul ? _GEN_4104 : _GEN_3606; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5505 = io_op_bits_active_vimul ? _GEN_4105 : _GEN_3607; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5506 = io_op_bits_active_vimul ? _GEN_4106 : _GEN_3608; // @[sequencer-master.scala 642:40]
  wire [9:0] _GEN_5507 = io_op_bits_active_vimul ? _GEN_4107 : _GEN_3609; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5508 = io_op_bits_active_vimul ? _GEN_4148 : _GEN_1688; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5509 = io_op_bits_active_vimul ? _GEN_4149 : _GEN_1689; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5510 = io_op_bits_active_vimul ? _GEN_4150 : _GEN_1690; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5511 = io_op_bits_active_vimul ? _GEN_4151 : _GEN_1691; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5512 = io_op_bits_active_vimul ? _GEN_4152 : _GEN_1692; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5513 = io_op_bits_active_vimul ? _GEN_4153 : _GEN_1693; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5514 = io_op_bits_active_vimul ? _GEN_4154 : _GEN_1694; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5515 = io_op_bits_active_vimul ? _GEN_4155 : _GEN_1695; // @[sequencer-master.scala 642:40]
  wire  _GEN_5516 = io_op_bits_active_vimul ? _GEN_4164 : _GEN_1696; // @[sequencer-master.scala 642:40]
  wire  _GEN_5517 = io_op_bits_active_vimul ? _GEN_4165 : _GEN_1697; // @[sequencer-master.scala 642:40]
  wire  _GEN_5518 = io_op_bits_active_vimul ? _GEN_4166 : _GEN_1698; // @[sequencer-master.scala 642:40]
  wire  _GEN_5519 = io_op_bits_active_vimul ? _GEN_4167 : _GEN_1699; // @[sequencer-master.scala 642:40]
  wire  _GEN_5520 = io_op_bits_active_vimul ? _GEN_4168 : _GEN_1700; // @[sequencer-master.scala 642:40]
  wire  _GEN_5521 = io_op_bits_active_vimul ? _GEN_4169 : _GEN_1701; // @[sequencer-master.scala 642:40]
  wire  _GEN_5522 = io_op_bits_active_vimul ? _GEN_4170 : _GEN_1702; // @[sequencer-master.scala 642:40]
  wire  _GEN_5523 = io_op_bits_active_vimul ? _GEN_4171 : _GEN_1703; // @[sequencer-master.scala 642:40]
  wire  _GEN_5524 = io_op_bits_active_vimul ? _GEN_4172 : _GEN_1704; // @[sequencer-master.scala 642:40]
  wire  _GEN_5525 = io_op_bits_active_vimul ? _GEN_4173 : _GEN_1705; // @[sequencer-master.scala 642:40]
  wire  _GEN_5526 = io_op_bits_active_vimul ? _GEN_4174 : _GEN_1706; // @[sequencer-master.scala 642:40]
  wire  _GEN_5527 = io_op_bits_active_vimul ? _GEN_4175 : _GEN_1707; // @[sequencer-master.scala 642:40]
  wire  _GEN_5528 = io_op_bits_active_vimul ? _GEN_4176 : _GEN_1708; // @[sequencer-master.scala 642:40]
  wire  _GEN_5529 = io_op_bits_active_vimul ? _GEN_4177 : _GEN_1709; // @[sequencer-master.scala 642:40]
  wire  _GEN_5530 = io_op_bits_active_vimul ? _GEN_4178 : _GEN_1710; // @[sequencer-master.scala 642:40]
  wire  _GEN_5531 = io_op_bits_active_vimul ? _GEN_4179 : _GEN_1711; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5532 = io_op_bits_active_vimul ? _GEN_4180 : _GEN_1712; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5533 = io_op_bits_active_vimul ? _GEN_4181 : _GEN_1713; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5534 = io_op_bits_active_vimul ? _GEN_4182 : _GEN_1714; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5535 = io_op_bits_active_vimul ? _GEN_4183 : _GEN_1715; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5536 = io_op_bits_active_vimul ? _GEN_4184 : _GEN_1716; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5537 = io_op_bits_active_vimul ? _GEN_4185 : _GEN_1717; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5538 = io_op_bits_active_vimul ? _GEN_4186 : _GEN_1718; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5539 = io_op_bits_active_vimul ? _GEN_4187 : _GEN_1719; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5540 = io_op_bits_active_vimul ? _GEN_4380 : _GEN_3610; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5541 = io_op_bits_active_vimul ? _GEN_4381 : _GEN_3611; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5542 = io_op_bits_active_vimul ? _GEN_4382 : _GEN_3612; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5543 = io_op_bits_active_vimul ? _GEN_4383 : _GEN_3613; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5544 = io_op_bits_active_vimul ? _GEN_4384 : _GEN_3614; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5545 = io_op_bits_active_vimul ? _GEN_4385 : _GEN_3615; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5546 = io_op_bits_active_vimul ? _GEN_4386 : _GEN_3616; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5547 = io_op_bits_active_vimul ? _GEN_4387 : _GEN_3617; // @[sequencer-master.scala 642:40]
  wire  _GEN_5548 = io_op_bits_active_vimul ? _GEN_4396 : _GEN_3618; // @[sequencer-master.scala 642:40]
  wire  _GEN_5549 = io_op_bits_active_vimul ? _GEN_4397 : _GEN_3619; // @[sequencer-master.scala 642:40]
  wire  _GEN_5550 = io_op_bits_active_vimul ? _GEN_4398 : _GEN_3620; // @[sequencer-master.scala 642:40]
  wire  _GEN_5551 = io_op_bits_active_vimul ? _GEN_4399 : _GEN_3621; // @[sequencer-master.scala 642:40]
  wire  _GEN_5552 = io_op_bits_active_vimul ? _GEN_4400 : _GEN_3622; // @[sequencer-master.scala 642:40]
  wire  _GEN_5553 = io_op_bits_active_vimul ? _GEN_4401 : _GEN_3623; // @[sequencer-master.scala 642:40]
  wire  _GEN_5554 = io_op_bits_active_vimul ? _GEN_4402 : _GEN_3624; // @[sequencer-master.scala 642:40]
  wire  _GEN_5555 = io_op_bits_active_vimul ? _GEN_4403 : _GEN_3625; // @[sequencer-master.scala 642:40]
  wire  _GEN_5556 = io_op_bits_active_vimul ? _GEN_4404 : _GEN_3626; // @[sequencer-master.scala 642:40]
  wire  _GEN_5557 = io_op_bits_active_vimul ? _GEN_4405 : _GEN_3627; // @[sequencer-master.scala 642:40]
  wire  _GEN_5558 = io_op_bits_active_vimul ? _GEN_4406 : _GEN_3628; // @[sequencer-master.scala 642:40]
  wire  _GEN_5559 = io_op_bits_active_vimul ? _GEN_4407 : _GEN_3629; // @[sequencer-master.scala 642:40]
  wire  _GEN_5560 = io_op_bits_active_vimul ? _GEN_4408 : _GEN_3630; // @[sequencer-master.scala 642:40]
  wire  _GEN_5561 = io_op_bits_active_vimul ? _GEN_4409 : _GEN_3631; // @[sequencer-master.scala 642:40]
  wire  _GEN_5562 = io_op_bits_active_vimul ? _GEN_4410 : _GEN_3632; // @[sequencer-master.scala 642:40]
  wire  _GEN_5563 = io_op_bits_active_vimul ? _GEN_4411 : _GEN_3633; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5564 = io_op_bits_active_vimul ? _GEN_4412 : _GEN_3634; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5565 = io_op_bits_active_vimul ? _GEN_4413 : _GEN_3635; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5566 = io_op_bits_active_vimul ? _GEN_4414 : _GEN_3636; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5567 = io_op_bits_active_vimul ? _GEN_4415 : _GEN_3637; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5568 = io_op_bits_active_vimul ? _GEN_4416 : _GEN_3638; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5569 = io_op_bits_active_vimul ? _GEN_4417 : _GEN_3639; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5570 = io_op_bits_active_vimul ? _GEN_4418 : _GEN_3640; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5571 = io_op_bits_active_vimul ? _GEN_4419 : _GEN_3641; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5572 = io_op_bits_active_vimul ? _GEN_4420 : _GEN_3642; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5573 = io_op_bits_active_vimul ? _GEN_4421 : _GEN_3643; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5574 = io_op_bits_active_vimul ? _GEN_4422 : _GEN_3644; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5575 = io_op_bits_active_vimul ? _GEN_4423 : _GEN_3645; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5576 = io_op_bits_active_vimul ? _GEN_4424 : _GEN_3646; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5577 = io_op_bits_active_vimul ? _GEN_4425 : _GEN_3647; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5578 = io_op_bits_active_vimul ? _GEN_4426 : _GEN_3648; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5579 = io_op_bits_active_vimul ? _GEN_4427 : _GEN_3649; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5580 = io_op_bits_active_vimul ? _GEN_4428 : _GEN_3650; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5581 = io_op_bits_active_vimul ? _GEN_4429 : _GEN_3651; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5582 = io_op_bits_active_vimul ? _GEN_4430 : _GEN_3652; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5583 = io_op_bits_active_vimul ? _GEN_4431 : _GEN_3653; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5584 = io_op_bits_active_vimul ? _GEN_4432 : _GEN_3654; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5585 = io_op_bits_active_vimul ? _GEN_4433 : _GEN_3655; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5586 = io_op_bits_active_vimul ? _GEN_4434 : _GEN_3656; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5587 = io_op_bits_active_vimul ? _GEN_4435 : _GEN_3657; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5588 = io_op_bits_active_vimul ? _GEN_4628 : _GEN_3658; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5589 = io_op_bits_active_vimul ? _GEN_4629 : _GEN_3659; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5590 = io_op_bits_active_vimul ? _GEN_4630 : _GEN_3660; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5591 = io_op_bits_active_vimul ? _GEN_4631 : _GEN_3661; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5592 = io_op_bits_active_vimul ? _GEN_4632 : _GEN_3662; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5593 = io_op_bits_active_vimul ? _GEN_4633 : _GEN_3663; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5594 = io_op_bits_active_vimul ? _GEN_4634 : _GEN_3664; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5595 = io_op_bits_active_vimul ? _GEN_4635 : _GEN_3665; // @[sequencer-master.scala 642:40]
  wire  _GEN_5596 = io_op_bits_active_vimul ? _GEN_4644 : _GEN_3666; // @[sequencer-master.scala 642:40]
  wire  _GEN_5597 = io_op_bits_active_vimul ? _GEN_4645 : _GEN_3667; // @[sequencer-master.scala 642:40]
  wire  _GEN_5598 = io_op_bits_active_vimul ? _GEN_4646 : _GEN_3668; // @[sequencer-master.scala 642:40]
  wire  _GEN_5599 = io_op_bits_active_vimul ? _GEN_4647 : _GEN_3669; // @[sequencer-master.scala 642:40]
  wire  _GEN_5600 = io_op_bits_active_vimul ? _GEN_4648 : _GEN_3670; // @[sequencer-master.scala 642:40]
  wire  _GEN_5601 = io_op_bits_active_vimul ? _GEN_4649 : _GEN_3671; // @[sequencer-master.scala 642:40]
  wire  _GEN_5602 = io_op_bits_active_vimul ? _GEN_4650 : _GEN_3672; // @[sequencer-master.scala 642:40]
  wire  _GEN_5603 = io_op_bits_active_vimul ? _GEN_4651 : _GEN_3673; // @[sequencer-master.scala 642:40]
  wire  _GEN_5604 = io_op_bits_active_vimul ? _GEN_4652 : _GEN_3674; // @[sequencer-master.scala 642:40]
  wire  _GEN_5605 = io_op_bits_active_vimul ? _GEN_4653 : _GEN_3675; // @[sequencer-master.scala 642:40]
  wire  _GEN_5606 = io_op_bits_active_vimul ? _GEN_4654 : _GEN_3676; // @[sequencer-master.scala 642:40]
  wire  _GEN_5607 = io_op_bits_active_vimul ? _GEN_4655 : _GEN_3677; // @[sequencer-master.scala 642:40]
  wire  _GEN_5608 = io_op_bits_active_vimul ? _GEN_4656 : _GEN_3678; // @[sequencer-master.scala 642:40]
  wire  _GEN_5609 = io_op_bits_active_vimul ? _GEN_4657 : _GEN_3679; // @[sequencer-master.scala 642:40]
  wire  _GEN_5610 = io_op_bits_active_vimul ? _GEN_4658 : _GEN_3680; // @[sequencer-master.scala 642:40]
  wire  _GEN_5611 = io_op_bits_active_vimul ? _GEN_4659 : _GEN_3681; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5612 = io_op_bits_active_vimul ? _GEN_4660 : _GEN_3682; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5613 = io_op_bits_active_vimul ? _GEN_4661 : _GEN_3683; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5614 = io_op_bits_active_vimul ? _GEN_4662 : _GEN_3684; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5615 = io_op_bits_active_vimul ? _GEN_4663 : _GEN_3685; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5616 = io_op_bits_active_vimul ? _GEN_4664 : _GEN_3686; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5617 = io_op_bits_active_vimul ? _GEN_4665 : _GEN_3687; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5618 = io_op_bits_active_vimul ? _GEN_4666 : _GEN_3688; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5619 = io_op_bits_active_vimul ? _GEN_4667 : _GEN_3689; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5620 = io_op_bits_active_vimul ? _GEN_4668 : _GEN_3690; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5621 = io_op_bits_active_vimul ? _GEN_4669 : _GEN_3691; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5622 = io_op_bits_active_vimul ? _GEN_4670 : _GEN_3692; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5623 = io_op_bits_active_vimul ? _GEN_4671 : _GEN_3693; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5624 = io_op_bits_active_vimul ? _GEN_4672 : _GEN_3694; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5625 = io_op_bits_active_vimul ? _GEN_4673 : _GEN_3695; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5626 = io_op_bits_active_vimul ? _GEN_4674 : _GEN_3696; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5627 = io_op_bits_active_vimul ? _GEN_4675 : _GEN_3697; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5628 = io_op_bits_active_vimul ? _GEN_4676 : _GEN_3698; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5629 = io_op_bits_active_vimul ? _GEN_4677 : _GEN_3699; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5630 = io_op_bits_active_vimul ? _GEN_4678 : _GEN_3700; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5631 = io_op_bits_active_vimul ? _GEN_4679 : _GEN_3701; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5632 = io_op_bits_active_vimul ? _GEN_4680 : _GEN_3702; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5633 = io_op_bits_active_vimul ? _GEN_4681 : _GEN_3703; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5634 = io_op_bits_active_vimul ? _GEN_4682 : _GEN_3704; // @[sequencer-master.scala 642:40]
  wire [63:0] _GEN_5635 = io_op_bits_active_vimul ? _GEN_4683 : _GEN_3705; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5636 = io_op_bits_active_vimul ? _GEN_4860 : _GEN_3754; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5637 = io_op_bits_active_vimul ? _GEN_4861 : _GEN_3755; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5638 = io_op_bits_active_vimul ? _GEN_4862 : _GEN_3756; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5639 = io_op_bits_active_vimul ? _GEN_4863 : _GEN_3757; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5640 = io_op_bits_active_vimul ? _GEN_4864 : _GEN_3758; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5641 = io_op_bits_active_vimul ? _GEN_4865 : _GEN_3759; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5642 = io_op_bits_active_vimul ? _GEN_4866 : _GEN_3760; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5643 = io_op_bits_active_vimul ? _GEN_4867 : _GEN_3761; // @[sequencer-master.scala 642:40]
  wire  _GEN_5644 = io_op_bits_active_vimul ? _GEN_4876 : _GEN_3762; // @[sequencer-master.scala 642:40]
  wire  _GEN_5645 = io_op_bits_active_vimul ? _GEN_4877 : _GEN_3763; // @[sequencer-master.scala 642:40]
  wire  _GEN_5646 = io_op_bits_active_vimul ? _GEN_4878 : _GEN_3764; // @[sequencer-master.scala 642:40]
  wire  _GEN_5647 = io_op_bits_active_vimul ? _GEN_4879 : _GEN_3765; // @[sequencer-master.scala 642:40]
  wire  _GEN_5648 = io_op_bits_active_vimul ? _GEN_4880 : _GEN_3766; // @[sequencer-master.scala 642:40]
  wire  _GEN_5649 = io_op_bits_active_vimul ? _GEN_4881 : _GEN_3767; // @[sequencer-master.scala 642:40]
  wire  _GEN_5650 = io_op_bits_active_vimul ? _GEN_4882 : _GEN_3768; // @[sequencer-master.scala 642:40]
  wire  _GEN_5651 = io_op_bits_active_vimul ? _GEN_4883 : _GEN_3769; // @[sequencer-master.scala 642:40]
  wire  _GEN_5652 = io_op_bits_active_vimul ? _GEN_4884 : _GEN_3770; // @[sequencer-master.scala 642:40]
  wire  _GEN_5653 = io_op_bits_active_vimul ? _GEN_4885 : _GEN_3771; // @[sequencer-master.scala 642:40]
  wire  _GEN_5654 = io_op_bits_active_vimul ? _GEN_4886 : _GEN_3772; // @[sequencer-master.scala 642:40]
  wire  _GEN_5655 = io_op_bits_active_vimul ? _GEN_4887 : _GEN_3773; // @[sequencer-master.scala 642:40]
  wire  _GEN_5656 = io_op_bits_active_vimul ? _GEN_4888 : _GEN_3774; // @[sequencer-master.scala 642:40]
  wire  _GEN_5657 = io_op_bits_active_vimul ? _GEN_4889 : _GEN_3775; // @[sequencer-master.scala 642:40]
  wire  _GEN_5658 = io_op_bits_active_vimul ? _GEN_4890 : _GEN_3776; // @[sequencer-master.scala 642:40]
  wire  _GEN_5659 = io_op_bits_active_vimul ? _GEN_4891 : _GEN_3777; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5660 = io_op_bits_active_vimul ? _GEN_4892 : _GEN_3778; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5661 = io_op_bits_active_vimul ? _GEN_4893 : _GEN_3779; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5662 = io_op_bits_active_vimul ? _GEN_4894 : _GEN_3780; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5663 = io_op_bits_active_vimul ? _GEN_4895 : _GEN_3781; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5664 = io_op_bits_active_vimul ? _GEN_4896 : _GEN_3782; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5665 = io_op_bits_active_vimul ? _GEN_4897 : _GEN_3783; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5666 = io_op_bits_active_vimul ? _GEN_4898 : _GEN_3784; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5667 = io_op_bits_active_vimul ? _GEN_4899 : _GEN_3785; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5668 = io_op_bits_active_vimul ? _GEN_4900 : _GEN_3786; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5669 = io_op_bits_active_vimul ? _GEN_4901 : _GEN_3787; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5670 = io_op_bits_active_vimul ? _GEN_4902 : _GEN_3788; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5671 = io_op_bits_active_vimul ? _GEN_4903 : _GEN_3789; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5672 = io_op_bits_active_vimul ? _GEN_4904 : _GEN_3790; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5673 = io_op_bits_active_vimul ? _GEN_4905 : _GEN_3791; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5674 = io_op_bits_active_vimul ? _GEN_4906 : _GEN_3792; // @[sequencer-master.scala 642:40]
  wire [7:0] _GEN_5675 = io_op_bits_active_vimul ? _GEN_4907 : _GEN_3793; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5676 = io_op_bits_active_vimul ? _GEN_5164 : _GEN_3794; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5677 = io_op_bits_active_vimul ? _GEN_5165 : _GEN_3795; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5678 = io_op_bits_active_vimul ? _GEN_5166 : _GEN_3796; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5679 = io_op_bits_active_vimul ? _GEN_5167 : _GEN_3797; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5680 = io_op_bits_active_vimul ? _GEN_5168 : _GEN_3798; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5681 = io_op_bits_active_vimul ? _GEN_5169 : _GEN_3799; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5682 = io_op_bits_active_vimul ? _GEN_5170 : _GEN_3800; // @[sequencer-master.scala 642:40]
  wire [1:0] _GEN_5683 = io_op_bits_active_vimul ? _GEN_5171 : _GEN_3801; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5684 = io_op_bits_active_vimul ? _GEN_5196 : _GEN_3802; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5685 = io_op_bits_active_vimul ? _GEN_5197 : _GEN_3803; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5686 = io_op_bits_active_vimul ? _GEN_5198 : _GEN_3804; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5687 = io_op_bits_active_vimul ? _GEN_5199 : _GEN_3805; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5688 = io_op_bits_active_vimul ? _GEN_5200 : _GEN_3806; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5689 = io_op_bits_active_vimul ? _GEN_5201 : _GEN_3807; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5690 = io_op_bits_active_vimul ? _GEN_5202 : _GEN_3808; // @[sequencer-master.scala 642:40]
  wire [3:0] _GEN_5691 = io_op_bits_active_vimul ? _GEN_5203 : _GEN_3809; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5692 = io_op_bits_active_vimul ? _GEN_5212 : _GEN_3810; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5693 = io_op_bits_active_vimul ? _GEN_5213 : _GEN_3811; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5694 = io_op_bits_active_vimul ? _GEN_5214 : _GEN_3812; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5695 = io_op_bits_active_vimul ? _GEN_5215 : _GEN_3813; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5696 = io_op_bits_active_vimul ? _GEN_5216 : _GEN_3814; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5697 = io_op_bits_active_vimul ? _GEN_5217 : _GEN_3815; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5698 = io_op_bits_active_vimul ? _GEN_5218 : _GEN_3816; // @[sequencer-master.scala 642:40]
  wire [2:0] _GEN_5699 = io_op_bits_active_vimul ? _GEN_5219 : _GEN_3817; // @[sequencer-master.scala 642:40]
  wire  _GEN_5700 = io_op_bits_active_vimul | _GEN_3818; // @[sequencer-master.scala 642:40 sequencer-master.scala 265:41]
  wire [2:0] _GEN_5701 = io_op_bits_active_vimul ? _T_1645 : _GEN_3819; // @[sequencer-master.scala 642:40 sequencer-master.scala 265:66]
  wire  _GEN_5718 = 3'h0 == tail ? 1'h0 : _GEN_5236; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5719 = 3'h1 == tail ? 1'h0 : _GEN_5237; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5720 = 3'h2 == tail ? 1'h0 : _GEN_5238; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5721 = 3'h3 == tail ? 1'h0 : _GEN_5239; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5722 = 3'h4 == tail ? 1'h0 : _GEN_5240; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5723 = 3'h5 == tail ? 1'h0 : _GEN_5241; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5724 = 3'h6 == tail ? 1'h0 : _GEN_5242; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5725 = 3'h7 == tail ? 1'h0 : _GEN_5243; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_5726 = 3'h0 == tail ? 1'h0 : _GEN_5244; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5727 = 3'h1 == tail ? 1'h0 : _GEN_5245; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5728 = 3'h2 == tail ? 1'h0 : _GEN_5246; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5729 = 3'h3 == tail ? 1'h0 : _GEN_5247; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5730 = 3'h4 == tail ? 1'h0 : _GEN_5248; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5731 = 3'h5 == tail ? 1'h0 : _GEN_5249; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5732 = 3'h6 == tail ? 1'h0 : _GEN_5250; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5733 = 3'h7 == tail ? 1'h0 : _GEN_5251; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_5734 = 3'h0 == tail ? 1'h0 : _GEN_5252; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5735 = 3'h1 == tail ? 1'h0 : _GEN_5253; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5736 = 3'h2 == tail ? 1'h0 : _GEN_5254; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5737 = 3'h3 == tail ? 1'h0 : _GEN_5255; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5738 = 3'h4 == tail ? 1'h0 : _GEN_5256; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5739 = 3'h5 == tail ? 1'h0 : _GEN_5257; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5740 = 3'h6 == tail ? 1'h0 : _GEN_5258; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5741 = 3'h7 == tail ? 1'h0 : _GEN_5259; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_5742 = 3'h0 == tail ? 1'h0 : _GEN_5260; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5743 = 3'h1 == tail ? 1'h0 : _GEN_5261; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5744 = 3'h2 == tail ? 1'h0 : _GEN_5262; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5745 = 3'h3 == tail ? 1'h0 : _GEN_5263; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5746 = 3'h4 == tail ? 1'h0 : _GEN_5264; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5747 = 3'h5 == tail ? 1'h0 : _GEN_5265; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5748 = 3'h6 == tail ? 1'h0 : _GEN_5266; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5749 = 3'h7 == tail ? 1'h0 : _GEN_5267; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_5750 = 3'h0 == tail ? 1'h0 : _GEN_5268; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5751 = 3'h1 == tail ? 1'h0 : _GEN_5269; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5752 = 3'h2 == tail ? 1'h0 : _GEN_5270; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5753 = 3'h3 == tail ? 1'h0 : _GEN_5271; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5754 = 3'h4 == tail ? 1'h0 : _GEN_5272; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5755 = 3'h5 == tail ? 1'h0 : _GEN_5273; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5756 = 3'h6 == tail ? 1'h0 : _GEN_5274; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5757 = 3'h7 == tail ? 1'h0 : _GEN_5275; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_5766 = 3'h0 == tail ? 1'h0 : _GEN_5284; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5767 = 3'h1 == tail ? 1'h0 : _GEN_5285; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5768 = 3'h2 == tail ? 1'h0 : _GEN_5286; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5769 = 3'h3 == tail ? 1'h0 : _GEN_5287; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5770 = 3'h4 == tail ? 1'h0 : _GEN_5288; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5771 = 3'h5 == tail ? 1'h0 : _GEN_5289; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5772 = 3'h6 == tail ? 1'h0 : _GEN_5290; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5773 = 3'h7 == tail ? 1'h0 : _GEN_5291; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5774 = 3'h0 == tail ? 1'h0 : _GEN_5292; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5775 = 3'h1 == tail ? 1'h0 : _GEN_5293; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5776 = 3'h2 == tail ? 1'h0 : _GEN_5294; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5777 = 3'h3 == tail ? 1'h0 : _GEN_5295; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5778 = 3'h4 == tail ? 1'h0 : _GEN_5296; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5779 = 3'h5 == tail ? 1'h0 : _GEN_5297; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5780 = 3'h6 == tail ? 1'h0 : _GEN_5298; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5781 = 3'h7 == tail ? 1'h0 : _GEN_5299; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5782 = 3'h0 == tail ? 1'h0 : _GEN_5300; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5783 = 3'h1 == tail ? 1'h0 : _GEN_5301; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5784 = 3'h2 == tail ? 1'h0 : _GEN_5302; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5785 = 3'h3 == tail ? 1'h0 : _GEN_5303; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5786 = 3'h4 == tail ? 1'h0 : _GEN_5304; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5787 = 3'h5 == tail ? 1'h0 : _GEN_5305; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5788 = 3'h6 == tail ? 1'h0 : _GEN_5306; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5789 = 3'h7 == tail ? 1'h0 : _GEN_5307; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5790 = 3'h0 == tail ? 1'h0 : _GEN_5308; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5791 = 3'h1 == tail ? 1'h0 : _GEN_5309; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5792 = 3'h2 == tail ? 1'h0 : _GEN_5310; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5793 = 3'h3 == tail ? 1'h0 : _GEN_5311; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5794 = 3'h4 == tail ? 1'h0 : _GEN_5312; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5795 = 3'h5 == tail ? 1'h0 : _GEN_5313; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5796 = 3'h6 == tail ? 1'h0 : _GEN_5314; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5797 = 3'h7 == tail ? 1'h0 : _GEN_5315; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5798 = 3'h0 == tail ? 1'h0 : _GEN_5316; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5799 = 3'h1 == tail ? 1'h0 : _GEN_5317; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5800 = 3'h2 == tail ? 1'h0 : _GEN_5318; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5801 = 3'h3 == tail ? 1'h0 : _GEN_5319; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5802 = 3'h4 == tail ? 1'h0 : _GEN_5320; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5803 = 3'h5 == tail ? 1'h0 : _GEN_5321; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5804 = 3'h6 == tail ? 1'h0 : _GEN_5322; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5805 = 3'h7 == tail ? 1'h0 : _GEN_5323; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5806 = 3'h0 == tail ? 1'h0 : _GEN_5324; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5807 = 3'h1 == tail ? 1'h0 : _GEN_5325; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5808 = 3'h2 == tail ? 1'h0 : _GEN_5326; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5809 = 3'h3 == tail ? 1'h0 : _GEN_5327; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5810 = 3'h4 == tail ? 1'h0 : _GEN_5328; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5811 = 3'h5 == tail ? 1'h0 : _GEN_5329; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5812 = 3'h6 == tail ? 1'h0 : _GEN_5330; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5813 = 3'h7 == tail ? 1'h0 : _GEN_5331; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5814 = 3'h0 == tail ? 1'h0 : _GEN_5332; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5815 = 3'h1 == tail ? 1'h0 : _GEN_5333; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5816 = 3'h2 == tail ? 1'h0 : _GEN_5334; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5817 = 3'h3 == tail ? 1'h0 : _GEN_5335; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5818 = 3'h4 == tail ? 1'h0 : _GEN_5336; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5819 = 3'h5 == tail ? 1'h0 : _GEN_5337; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5820 = 3'h6 == tail ? 1'h0 : _GEN_5338; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5821 = 3'h7 == tail ? 1'h0 : _GEN_5339; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5822 = 3'h0 == tail ? 1'h0 : _GEN_5340; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5823 = 3'h1 == tail ? 1'h0 : _GEN_5341; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5824 = 3'h2 == tail ? 1'h0 : _GEN_5342; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5825 = 3'h3 == tail ? 1'h0 : _GEN_5343; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5826 = 3'h4 == tail ? 1'h0 : _GEN_5344; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5827 = 3'h5 == tail ? 1'h0 : _GEN_5345; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5828 = 3'h6 == tail ? 1'h0 : _GEN_5346; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5829 = 3'h7 == tail ? 1'h0 : _GEN_5347; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5830 = 3'h0 == tail ? 1'h0 : _GEN_5348; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5831 = 3'h1 == tail ? 1'h0 : _GEN_5349; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5832 = 3'h2 == tail ? 1'h0 : _GEN_5350; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5833 = 3'h3 == tail ? 1'h0 : _GEN_5351; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5834 = 3'h4 == tail ? 1'h0 : _GEN_5352; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5835 = 3'h5 == tail ? 1'h0 : _GEN_5353; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5836 = 3'h6 == tail ? 1'h0 : _GEN_5354; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5837 = 3'h7 == tail ? 1'h0 : _GEN_5355; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5838 = 3'h0 == tail ? 1'h0 : _GEN_5356; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5839 = 3'h1 == tail ? 1'h0 : _GEN_5357; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5840 = 3'h2 == tail ? 1'h0 : _GEN_5358; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5841 = 3'h3 == tail ? 1'h0 : _GEN_5359; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5842 = 3'h4 == tail ? 1'h0 : _GEN_5360; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5843 = 3'h5 == tail ? 1'h0 : _GEN_5361; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5844 = 3'h6 == tail ? 1'h0 : _GEN_5362; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5845 = 3'h7 == tail ? 1'h0 : _GEN_5363; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5846 = 3'h0 == tail ? 1'h0 : _GEN_5364; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5847 = 3'h1 == tail ? 1'h0 : _GEN_5365; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5848 = 3'h2 == tail ? 1'h0 : _GEN_5366; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5849 = 3'h3 == tail ? 1'h0 : _GEN_5367; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5850 = 3'h4 == tail ? 1'h0 : _GEN_5368; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5851 = 3'h5 == tail ? 1'h0 : _GEN_5369; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5852 = 3'h6 == tail ? 1'h0 : _GEN_5370; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5853 = 3'h7 == tail ? 1'h0 : _GEN_5371; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5854 = 3'h0 == tail ? 1'h0 : _GEN_5372; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5855 = 3'h1 == tail ? 1'h0 : _GEN_5373; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5856 = 3'h2 == tail ? 1'h0 : _GEN_5374; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5857 = 3'h3 == tail ? 1'h0 : _GEN_5375; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5858 = 3'h4 == tail ? 1'h0 : _GEN_5376; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5859 = 3'h5 == tail ? 1'h0 : _GEN_5377; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5860 = 3'h6 == tail ? 1'h0 : _GEN_5378; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5861 = 3'h7 == tail ? 1'h0 : _GEN_5379; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5862 = 3'h0 == tail ? 1'h0 : _GEN_5380; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5863 = 3'h1 == tail ? 1'h0 : _GEN_5381; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5864 = 3'h2 == tail ? 1'h0 : _GEN_5382; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5865 = 3'h3 == tail ? 1'h0 : _GEN_5383; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5866 = 3'h4 == tail ? 1'h0 : _GEN_5384; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5867 = 3'h5 == tail ? 1'h0 : _GEN_5385; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5868 = 3'h6 == tail ? 1'h0 : _GEN_5386; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5869 = 3'h7 == tail ? 1'h0 : _GEN_5387; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5870 = 3'h0 == tail ? 1'h0 : _GEN_5388; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5871 = 3'h1 == tail ? 1'h0 : _GEN_5389; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5872 = 3'h2 == tail ? 1'h0 : _GEN_5390; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5873 = 3'h3 == tail ? 1'h0 : _GEN_5391; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5874 = 3'h4 == tail ? 1'h0 : _GEN_5392; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5875 = 3'h5 == tail ? 1'h0 : _GEN_5393; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5876 = 3'h6 == tail ? 1'h0 : _GEN_5394; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5877 = 3'h7 == tail ? 1'h0 : _GEN_5395; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5878 = 3'h0 == tail ? 1'h0 : _GEN_5396; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5879 = 3'h1 == tail ? 1'h0 : _GEN_5397; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5880 = 3'h2 == tail ? 1'h0 : _GEN_5398; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5881 = 3'h3 == tail ? 1'h0 : _GEN_5399; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5882 = 3'h4 == tail ? 1'h0 : _GEN_5400; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5883 = 3'h5 == tail ? 1'h0 : _GEN_5401; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5884 = 3'h6 == tail ? 1'h0 : _GEN_5402; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5885 = 3'h7 == tail ? 1'h0 : _GEN_5403; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5886 = 3'h0 == tail ? 1'h0 : _GEN_5404; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5887 = 3'h1 == tail ? 1'h0 : _GEN_5405; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5888 = 3'h2 == tail ? 1'h0 : _GEN_5406; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5889 = 3'h3 == tail ? 1'h0 : _GEN_5407; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5890 = 3'h4 == tail ? 1'h0 : _GEN_5408; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5891 = 3'h5 == tail ? 1'h0 : _GEN_5409; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5892 = 3'h6 == tail ? 1'h0 : _GEN_5410; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5893 = 3'h7 == tail ? 1'h0 : _GEN_5411; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5894 = 3'h0 == tail ? 1'h0 : _GEN_5412; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5895 = 3'h1 == tail ? 1'h0 : _GEN_5413; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5896 = 3'h2 == tail ? 1'h0 : _GEN_5414; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5897 = 3'h3 == tail ? 1'h0 : _GEN_5415; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5898 = 3'h4 == tail ? 1'h0 : _GEN_5416; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5899 = 3'h5 == tail ? 1'h0 : _GEN_5417; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5900 = 3'h6 == tail ? 1'h0 : _GEN_5418; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5901 = 3'h7 == tail ? 1'h0 : _GEN_5419; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5902 = 3'h0 == tail ? 1'h0 : _GEN_5420; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5903 = 3'h1 == tail ? 1'h0 : _GEN_5421; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5904 = 3'h2 == tail ? 1'h0 : _GEN_5422; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5905 = 3'h3 == tail ? 1'h0 : _GEN_5423; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5906 = 3'h4 == tail ? 1'h0 : _GEN_5424; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5907 = 3'h5 == tail ? 1'h0 : _GEN_5425; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5908 = 3'h6 == tail ? 1'h0 : _GEN_5426; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5909 = 3'h7 == tail ? 1'h0 : _GEN_5427; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5910 = 3'h0 == tail ? 1'h0 : _GEN_5428; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5911 = 3'h1 == tail ? 1'h0 : _GEN_5429; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5912 = 3'h2 == tail ? 1'h0 : _GEN_5430; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5913 = 3'h3 == tail ? 1'h0 : _GEN_5431; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5914 = 3'h4 == tail ? 1'h0 : _GEN_5432; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5915 = 3'h5 == tail ? 1'h0 : _GEN_5433; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5916 = 3'h6 == tail ? 1'h0 : _GEN_5434; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5917 = 3'h7 == tail ? 1'h0 : _GEN_5435; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5918 = 3'h0 == tail ? 1'h0 : _GEN_5436; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5919 = 3'h1 == tail ? 1'h0 : _GEN_5437; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5920 = 3'h2 == tail ? 1'h0 : _GEN_5438; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5921 = 3'h3 == tail ? 1'h0 : _GEN_5439; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5922 = 3'h4 == tail ? 1'h0 : _GEN_5440; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5923 = 3'h5 == tail ? 1'h0 : _GEN_5441; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5924 = 3'h6 == tail ? 1'h0 : _GEN_5442; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5925 = 3'h7 == tail ? 1'h0 : _GEN_5443; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5926 = 3'h0 == tail ? 1'h0 : _GEN_5444; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5927 = 3'h1 == tail ? 1'h0 : _GEN_5445; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5928 = 3'h2 == tail ? 1'h0 : _GEN_5446; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5929 = 3'h3 == tail ? 1'h0 : _GEN_5447; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5930 = 3'h4 == tail ? 1'h0 : _GEN_5448; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5931 = 3'h5 == tail ? 1'h0 : _GEN_5449; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5932 = 3'h6 == tail ? 1'h0 : _GEN_5450; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5933 = 3'h7 == tail ? 1'h0 : _GEN_5451; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5934 = 3'h0 == tail ? 1'h0 : _GEN_5452; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5935 = 3'h1 == tail ? 1'h0 : _GEN_5453; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5936 = 3'h2 == tail ? 1'h0 : _GEN_5454; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5937 = 3'h3 == tail ? 1'h0 : _GEN_5455; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5938 = 3'h4 == tail ? 1'h0 : _GEN_5456; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5939 = 3'h5 == tail ? 1'h0 : _GEN_5457; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5940 = 3'h6 == tail ? 1'h0 : _GEN_5458; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5941 = 3'h7 == tail ? 1'h0 : _GEN_5459; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_5942 = 3'h0 == tail ? 1'h0 : _GEN_5460; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5943 = 3'h1 == tail ? 1'h0 : _GEN_5461; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5944 = 3'h2 == tail ? 1'h0 : _GEN_5462; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5945 = 3'h3 == tail ? 1'h0 : _GEN_5463; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5946 = 3'h4 == tail ? 1'h0 : _GEN_5464; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5947 = 3'h5 == tail ? 1'h0 : _GEN_5465; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5948 = 3'h6 == tail ? 1'h0 : _GEN_5466; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5949 = 3'h7 == tail ? 1'h0 : _GEN_5467; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_5950 = 3'h0 == tail ? 1'h0 : _GEN_5468; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5951 = 3'h1 == tail ? 1'h0 : _GEN_5469; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5952 = 3'h2 == tail ? 1'h0 : _GEN_5470; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5953 = 3'h3 == tail ? 1'h0 : _GEN_5471; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5954 = 3'h4 == tail ? 1'h0 : _GEN_5472; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5955 = 3'h5 == tail ? 1'h0 : _GEN_5473; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5956 = 3'h6 == tail ? 1'h0 : _GEN_5474; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5957 = 3'h7 == tail ? 1'h0 : _GEN_5475; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_5958 = 3'h0 == tail ? 1'h0 : _GEN_5476; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5959 = 3'h1 == tail ? 1'h0 : _GEN_5477; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5960 = 3'h2 == tail ? 1'h0 : _GEN_5478; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5961 = 3'h3 == tail ? 1'h0 : _GEN_5479; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5962 = 3'h4 == tail ? 1'h0 : _GEN_5480; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5963 = 3'h5 == tail ? 1'h0 : _GEN_5481; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5964 = 3'h6 == tail ? 1'h0 : _GEN_5482; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5965 = 3'h7 == tail ? 1'h0 : _GEN_5483; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_5974 = _GEN_32729 | e_0_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5975 = _GEN_32730 | e_1_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5976 = _GEN_32731 | e_2_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5977 = _GEN_32732 | e_3_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5978 = _GEN_32733 | e_4_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5979 = _GEN_32734 | e_5_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5980 = _GEN_32735 | e_6_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_5981 = _GEN_32736 | e_7_active_vqu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _T_1884 = io_op_bits_active_vidiv | io_op_bits_active_vfdiv; // @[sequencer-master.scala 298:31]
  wire  _T_1895 = ~io_op_bits_fn_union[0]; // @[types-vxu.scala 54:51]
  wire  _T_1897 = io_op_bits_active_vidiv | io_op_bits_active_vfdiv & _T_1895; // @[sequencer-master.scala 300:28]
  wire  _T_1899 = _T_1884 | io_op_bits_active_vrfirst; // @[sequencer-master.scala 301:46]
  wire [1:0] _T_1900 = {_T_1897,_T_1899}; // @[Cat.scala 30:58]
  wire [9:0] _e_tail_fn_union_2 = {{8'd0}, _T_1900}; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5982 = 3'h0 == tail ? _e_tail_fn_union_2 : _GEN_5500; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5983 = 3'h1 == tail ? _e_tail_fn_union_2 : _GEN_5501; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5984 = 3'h2 == tail ? _e_tail_fn_union_2 : _GEN_5502; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5985 = 3'h3 == tail ? _e_tail_fn_union_2 : _GEN_5503; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5986 = 3'h4 == tail ? _e_tail_fn_union_2 : _GEN_5504; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5987 = 3'h5 == tail ? _e_tail_fn_union_2 : _GEN_5505; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5988 = 3'h6 == tail ? _e_tail_fn_union_2 : _GEN_5506; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_5989 = 3'h7 == tail ? _e_tail_fn_union_2 : _GEN_5507; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_5990 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_5508; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5991 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_5509; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5992 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_5510; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5993 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_5511; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5994 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_5512; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5995 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_5513; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5996 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_5514; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_5997 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_5515; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_5998 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_5718; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_5999 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_5719; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6000 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_5720; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6001 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_5721; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6002 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_5722; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6003 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_5723; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6004 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_5724; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6005 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_5725; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6006 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_5516; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6007 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_5517; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6008 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_5518; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6009 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_5519; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6010 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_5520; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6011 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_5521; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6012 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_5522; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6013 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_5523; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6014 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_5524; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6015 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_5525; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6016 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_5526; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6017 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_5527; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6018 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_5528; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6019 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_5529; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6020 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_5530; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_6021 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_5531; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_6022 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_5532; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6023 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_5533; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6024 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_5534; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6025 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_5535; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6026 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_5536; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6027 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_5537; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6028 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_5538; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_6029 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_5539; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_6030 = io_op_bits_base_vp_valid ? _GEN_5990 : _GEN_5508; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6031 = io_op_bits_base_vp_valid ? _GEN_5991 : _GEN_5509; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6032 = io_op_bits_base_vp_valid ? _GEN_5992 : _GEN_5510; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6033 = io_op_bits_base_vp_valid ? _GEN_5993 : _GEN_5511; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6034 = io_op_bits_base_vp_valid ? _GEN_5994 : _GEN_5512; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6035 = io_op_bits_base_vp_valid ? _GEN_5995 : _GEN_5513; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6036 = io_op_bits_base_vp_valid ? _GEN_5996 : _GEN_5514; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_6037 = io_op_bits_base_vp_valid ? _GEN_5997 : _GEN_5515; // @[sequencer-master.scala 320:41]
  wire  _GEN_6038 = io_op_bits_base_vp_valid ? _GEN_5998 : _GEN_5718; // @[sequencer-master.scala 320:41]
  wire  _GEN_6039 = io_op_bits_base_vp_valid ? _GEN_5999 : _GEN_5719; // @[sequencer-master.scala 320:41]
  wire  _GEN_6040 = io_op_bits_base_vp_valid ? _GEN_6000 : _GEN_5720; // @[sequencer-master.scala 320:41]
  wire  _GEN_6041 = io_op_bits_base_vp_valid ? _GEN_6001 : _GEN_5721; // @[sequencer-master.scala 320:41]
  wire  _GEN_6042 = io_op_bits_base_vp_valid ? _GEN_6002 : _GEN_5722; // @[sequencer-master.scala 320:41]
  wire  _GEN_6043 = io_op_bits_base_vp_valid ? _GEN_6003 : _GEN_5723; // @[sequencer-master.scala 320:41]
  wire  _GEN_6044 = io_op_bits_base_vp_valid ? _GEN_6004 : _GEN_5724; // @[sequencer-master.scala 320:41]
  wire  _GEN_6045 = io_op_bits_base_vp_valid ? _GEN_6005 : _GEN_5725; // @[sequencer-master.scala 320:41]
  wire  _GEN_6046 = io_op_bits_base_vp_valid ? _GEN_6006 : _GEN_5516; // @[sequencer-master.scala 320:41]
  wire  _GEN_6047 = io_op_bits_base_vp_valid ? _GEN_6007 : _GEN_5517; // @[sequencer-master.scala 320:41]
  wire  _GEN_6048 = io_op_bits_base_vp_valid ? _GEN_6008 : _GEN_5518; // @[sequencer-master.scala 320:41]
  wire  _GEN_6049 = io_op_bits_base_vp_valid ? _GEN_6009 : _GEN_5519; // @[sequencer-master.scala 320:41]
  wire  _GEN_6050 = io_op_bits_base_vp_valid ? _GEN_6010 : _GEN_5520; // @[sequencer-master.scala 320:41]
  wire  _GEN_6051 = io_op_bits_base_vp_valid ? _GEN_6011 : _GEN_5521; // @[sequencer-master.scala 320:41]
  wire  _GEN_6052 = io_op_bits_base_vp_valid ? _GEN_6012 : _GEN_5522; // @[sequencer-master.scala 320:41]
  wire  _GEN_6053 = io_op_bits_base_vp_valid ? _GEN_6013 : _GEN_5523; // @[sequencer-master.scala 320:41]
  wire  _GEN_6054 = io_op_bits_base_vp_valid ? _GEN_6014 : _GEN_5524; // @[sequencer-master.scala 320:41]
  wire  _GEN_6055 = io_op_bits_base_vp_valid ? _GEN_6015 : _GEN_5525; // @[sequencer-master.scala 320:41]
  wire  _GEN_6056 = io_op_bits_base_vp_valid ? _GEN_6016 : _GEN_5526; // @[sequencer-master.scala 320:41]
  wire  _GEN_6057 = io_op_bits_base_vp_valid ? _GEN_6017 : _GEN_5527; // @[sequencer-master.scala 320:41]
  wire  _GEN_6058 = io_op_bits_base_vp_valid ? _GEN_6018 : _GEN_5528; // @[sequencer-master.scala 320:41]
  wire  _GEN_6059 = io_op_bits_base_vp_valid ? _GEN_6019 : _GEN_5529; // @[sequencer-master.scala 320:41]
  wire  _GEN_6060 = io_op_bits_base_vp_valid ? _GEN_6020 : _GEN_5530; // @[sequencer-master.scala 320:41]
  wire  _GEN_6061 = io_op_bits_base_vp_valid ? _GEN_6021 : _GEN_5531; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6062 = io_op_bits_base_vp_valid ? _GEN_6022 : _GEN_5532; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6063 = io_op_bits_base_vp_valid ? _GEN_6023 : _GEN_5533; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6064 = io_op_bits_base_vp_valid ? _GEN_6024 : _GEN_5534; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6065 = io_op_bits_base_vp_valid ? _GEN_6025 : _GEN_5535; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6066 = io_op_bits_base_vp_valid ? _GEN_6026 : _GEN_5536; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6067 = io_op_bits_base_vp_valid ? _GEN_6027 : _GEN_5537; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6068 = io_op_bits_base_vp_valid ? _GEN_6028 : _GEN_5538; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_6069 = io_op_bits_base_vp_valid ? _GEN_6029 : _GEN_5539; // @[sequencer-master.scala 320:41]
  wire  _GEN_6070 = _GEN_32729 | _GEN_5766; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6071 = _GEN_32730 | _GEN_5767; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6072 = _GEN_32731 | _GEN_5768; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6073 = _GEN_32732 | _GEN_5769; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6074 = _GEN_32733 | _GEN_5770; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6075 = _GEN_32734 | _GEN_5771; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6076 = _GEN_32735 | _GEN_5772; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6077 = _GEN_32736 | _GEN_5773; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6078 = _T_26 ? _GEN_6070 : _GEN_5766; // @[sequencer-master.scala 154:24]
  wire  _GEN_6079 = _T_26 ? _GEN_6071 : _GEN_5767; // @[sequencer-master.scala 154:24]
  wire  _GEN_6080 = _T_26 ? _GEN_6072 : _GEN_5768; // @[sequencer-master.scala 154:24]
  wire  _GEN_6081 = _T_26 ? _GEN_6073 : _GEN_5769; // @[sequencer-master.scala 154:24]
  wire  _GEN_6082 = _T_26 ? _GEN_6074 : _GEN_5770; // @[sequencer-master.scala 154:24]
  wire  _GEN_6083 = _T_26 ? _GEN_6075 : _GEN_5771; // @[sequencer-master.scala 154:24]
  wire  _GEN_6084 = _T_26 ? _GEN_6076 : _GEN_5772; // @[sequencer-master.scala 154:24]
  wire  _GEN_6085 = _T_26 ? _GEN_6077 : _GEN_5773; // @[sequencer-master.scala 154:24]
  wire  _GEN_6086 = _GEN_32729 | _GEN_5790; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6087 = _GEN_32730 | _GEN_5791; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6088 = _GEN_32731 | _GEN_5792; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6089 = _GEN_32732 | _GEN_5793; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6090 = _GEN_32733 | _GEN_5794; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6091 = _GEN_32734 | _GEN_5795; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6092 = _GEN_32735 | _GEN_5796; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6093 = _GEN_32736 | _GEN_5797; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6094 = _T_48 ? _GEN_6086 : _GEN_5790; // @[sequencer-master.scala 154:24]
  wire  _GEN_6095 = _T_48 ? _GEN_6087 : _GEN_5791; // @[sequencer-master.scala 154:24]
  wire  _GEN_6096 = _T_48 ? _GEN_6088 : _GEN_5792; // @[sequencer-master.scala 154:24]
  wire  _GEN_6097 = _T_48 ? _GEN_6089 : _GEN_5793; // @[sequencer-master.scala 154:24]
  wire  _GEN_6098 = _T_48 ? _GEN_6090 : _GEN_5794; // @[sequencer-master.scala 154:24]
  wire  _GEN_6099 = _T_48 ? _GEN_6091 : _GEN_5795; // @[sequencer-master.scala 154:24]
  wire  _GEN_6100 = _T_48 ? _GEN_6092 : _GEN_5796; // @[sequencer-master.scala 154:24]
  wire  _GEN_6101 = _T_48 ? _GEN_6093 : _GEN_5797; // @[sequencer-master.scala 154:24]
  wire  _GEN_6102 = _GEN_32729 | _GEN_5814; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6103 = _GEN_32730 | _GEN_5815; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6104 = _GEN_32731 | _GEN_5816; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6105 = _GEN_32732 | _GEN_5817; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6106 = _GEN_32733 | _GEN_5818; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6107 = _GEN_32734 | _GEN_5819; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6108 = _GEN_32735 | _GEN_5820; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6109 = _GEN_32736 | _GEN_5821; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6110 = _T_70 ? _GEN_6102 : _GEN_5814; // @[sequencer-master.scala 154:24]
  wire  _GEN_6111 = _T_70 ? _GEN_6103 : _GEN_5815; // @[sequencer-master.scala 154:24]
  wire  _GEN_6112 = _T_70 ? _GEN_6104 : _GEN_5816; // @[sequencer-master.scala 154:24]
  wire  _GEN_6113 = _T_70 ? _GEN_6105 : _GEN_5817; // @[sequencer-master.scala 154:24]
  wire  _GEN_6114 = _T_70 ? _GEN_6106 : _GEN_5818; // @[sequencer-master.scala 154:24]
  wire  _GEN_6115 = _T_70 ? _GEN_6107 : _GEN_5819; // @[sequencer-master.scala 154:24]
  wire  _GEN_6116 = _T_70 ? _GEN_6108 : _GEN_5820; // @[sequencer-master.scala 154:24]
  wire  _GEN_6117 = _T_70 ? _GEN_6109 : _GEN_5821; // @[sequencer-master.scala 154:24]
  wire  _GEN_6118 = _GEN_32729 | _GEN_5838; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6119 = _GEN_32730 | _GEN_5839; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6120 = _GEN_32731 | _GEN_5840; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6121 = _GEN_32732 | _GEN_5841; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6122 = _GEN_32733 | _GEN_5842; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6123 = _GEN_32734 | _GEN_5843; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6124 = _GEN_32735 | _GEN_5844; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6125 = _GEN_32736 | _GEN_5845; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6126 = _T_92 ? _GEN_6118 : _GEN_5838; // @[sequencer-master.scala 154:24]
  wire  _GEN_6127 = _T_92 ? _GEN_6119 : _GEN_5839; // @[sequencer-master.scala 154:24]
  wire  _GEN_6128 = _T_92 ? _GEN_6120 : _GEN_5840; // @[sequencer-master.scala 154:24]
  wire  _GEN_6129 = _T_92 ? _GEN_6121 : _GEN_5841; // @[sequencer-master.scala 154:24]
  wire  _GEN_6130 = _T_92 ? _GEN_6122 : _GEN_5842; // @[sequencer-master.scala 154:24]
  wire  _GEN_6131 = _T_92 ? _GEN_6123 : _GEN_5843; // @[sequencer-master.scala 154:24]
  wire  _GEN_6132 = _T_92 ? _GEN_6124 : _GEN_5844; // @[sequencer-master.scala 154:24]
  wire  _GEN_6133 = _T_92 ? _GEN_6125 : _GEN_5845; // @[sequencer-master.scala 154:24]
  wire  _GEN_6134 = _GEN_32729 | _GEN_5862; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6135 = _GEN_32730 | _GEN_5863; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6136 = _GEN_32731 | _GEN_5864; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6137 = _GEN_32732 | _GEN_5865; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6138 = _GEN_32733 | _GEN_5866; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6139 = _GEN_32734 | _GEN_5867; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6140 = _GEN_32735 | _GEN_5868; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6141 = _GEN_32736 | _GEN_5869; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6142 = _T_114 ? _GEN_6134 : _GEN_5862; // @[sequencer-master.scala 154:24]
  wire  _GEN_6143 = _T_114 ? _GEN_6135 : _GEN_5863; // @[sequencer-master.scala 154:24]
  wire  _GEN_6144 = _T_114 ? _GEN_6136 : _GEN_5864; // @[sequencer-master.scala 154:24]
  wire  _GEN_6145 = _T_114 ? _GEN_6137 : _GEN_5865; // @[sequencer-master.scala 154:24]
  wire  _GEN_6146 = _T_114 ? _GEN_6138 : _GEN_5866; // @[sequencer-master.scala 154:24]
  wire  _GEN_6147 = _T_114 ? _GEN_6139 : _GEN_5867; // @[sequencer-master.scala 154:24]
  wire  _GEN_6148 = _T_114 ? _GEN_6140 : _GEN_5868; // @[sequencer-master.scala 154:24]
  wire  _GEN_6149 = _T_114 ? _GEN_6141 : _GEN_5869; // @[sequencer-master.scala 154:24]
  wire  _GEN_6150 = _GEN_32729 | _GEN_5886; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6151 = _GEN_32730 | _GEN_5887; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6152 = _GEN_32731 | _GEN_5888; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6153 = _GEN_32732 | _GEN_5889; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6154 = _GEN_32733 | _GEN_5890; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6155 = _GEN_32734 | _GEN_5891; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6156 = _GEN_32735 | _GEN_5892; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6157 = _GEN_32736 | _GEN_5893; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6158 = _T_136 ? _GEN_6150 : _GEN_5886; // @[sequencer-master.scala 154:24]
  wire  _GEN_6159 = _T_136 ? _GEN_6151 : _GEN_5887; // @[sequencer-master.scala 154:24]
  wire  _GEN_6160 = _T_136 ? _GEN_6152 : _GEN_5888; // @[sequencer-master.scala 154:24]
  wire  _GEN_6161 = _T_136 ? _GEN_6153 : _GEN_5889; // @[sequencer-master.scala 154:24]
  wire  _GEN_6162 = _T_136 ? _GEN_6154 : _GEN_5890; // @[sequencer-master.scala 154:24]
  wire  _GEN_6163 = _T_136 ? _GEN_6155 : _GEN_5891; // @[sequencer-master.scala 154:24]
  wire  _GEN_6164 = _T_136 ? _GEN_6156 : _GEN_5892; // @[sequencer-master.scala 154:24]
  wire  _GEN_6165 = _T_136 ? _GEN_6157 : _GEN_5893; // @[sequencer-master.scala 154:24]
  wire  _GEN_6166 = _GEN_32729 | _GEN_5910; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6167 = _GEN_32730 | _GEN_5911; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6168 = _GEN_32731 | _GEN_5912; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6169 = _GEN_32732 | _GEN_5913; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6170 = _GEN_32733 | _GEN_5914; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6171 = _GEN_32734 | _GEN_5915; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6172 = _GEN_32735 | _GEN_5916; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6173 = _GEN_32736 | _GEN_5917; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6174 = _T_158 ? _GEN_6166 : _GEN_5910; // @[sequencer-master.scala 154:24]
  wire  _GEN_6175 = _T_158 ? _GEN_6167 : _GEN_5911; // @[sequencer-master.scala 154:24]
  wire  _GEN_6176 = _T_158 ? _GEN_6168 : _GEN_5912; // @[sequencer-master.scala 154:24]
  wire  _GEN_6177 = _T_158 ? _GEN_6169 : _GEN_5913; // @[sequencer-master.scala 154:24]
  wire  _GEN_6178 = _T_158 ? _GEN_6170 : _GEN_5914; // @[sequencer-master.scala 154:24]
  wire  _GEN_6179 = _T_158 ? _GEN_6171 : _GEN_5915; // @[sequencer-master.scala 154:24]
  wire  _GEN_6180 = _T_158 ? _GEN_6172 : _GEN_5916; // @[sequencer-master.scala 154:24]
  wire  _GEN_6181 = _T_158 ? _GEN_6173 : _GEN_5917; // @[sequencer-master.scala 154:24]
  wire  _GEN_6182 = _GEN_32729 | _GEN_5934; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6183 = _GEN_32730 | _GEN_5935; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6184 = _GEN_32731 | _GEN_5936; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6185 = _GEN_32732 | _GEN_5937; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6186 = _GEN_32733 | _GEN_5938; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6187 = _GEN_32734 | _GEN_5939; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6188 = _GEN_32735 | _GEN_5940; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6189 = _GEN_32736 | _GEN_5941; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6190 = _T_180 ? _GEN_6182 : _GEN_5934; // @[sequencer-master.scala 154:24]
  wire  _GEN_6191 = _T_180 ? _GEN_6183 : _GEN_5935; // @[sequencer-master.scala 154:24]
  wire  _GEN_6192 = _T_180 ? _GEN_6184 : _GEN_5936; // @[sequencer-master.scala 154:24]
  wire  _GEN_6193 = _T_180 ? _GEN_6185 : _GEN_5937; // @[sequencer-master.scala 154:24]
  wire  _GEN_6194 = _T_180 ? _GEN_6186 : _GEN_5938; // @[sequencer-master.scala 154:24]
  wire  _GEN_6195 = _T_180 ? _GEN_6187 : _GEN_5939; // @[sequencer-master.scala 154:24]
  wire  _GEN_6196 = _T_180 ? _GEN_6188 : _GEN_5940; // @[sequencer-master.scala 154:24]
  wire  _GEN_6197 = _T_180 ? _GEN_6189 : _GEN_5941; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_6198 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_5540; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6199 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_5541; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6200 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_5542; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6201 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_5543; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6202 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_5544; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6203 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_5545; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6204 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_5546; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6205 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_5547; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6206 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_5726; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6207 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_5727; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6208 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_5728; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6209 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_5729; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6210 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_5730; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6211 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_5731; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6212 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_5732; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6213 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_5733; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6214 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_5548; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6215 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_5549; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6216 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_5550; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6217 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_5551; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6218 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_5552; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6219 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_5553; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6220 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_5554; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6221 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_5555; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6222 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_5556; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6223 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_5557; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6224 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_5558; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6225 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_5559; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6226 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_5560; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6227 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_5561; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6228 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_5562; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6229 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_5563; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6230 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_5564; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6231 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_5565; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6232 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_5566; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6233 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_5567; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6234 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_5568; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6235 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_5569; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6236 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_5570; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6237 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_5571; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6238 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_5572; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6239 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_5573; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6240 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_5574; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6241 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_5575; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6242 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_5576; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6243 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_5577; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6244 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_5578; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6245 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_5579; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_6246 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_5580; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6247 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_5581; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6248 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_5582; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6249 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_5583; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6250 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_5584; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6251 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_5585; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6252 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_5586; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6253 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_5587; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6254 = _T_189 ? _GEN_6246 : _GEN_5580; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6255 = _T_189 ? _GEN_6247 : _GEN_5581; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6256 = _T_189 ? _GEN_6248 : _GEN_5582; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6257 = _T_189 ? _GEN_6249 : _GEN_5583; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6258 = _T_189 ? _GEN_6250 : _GEN_5584; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6259 = _T_189 ? _GEN_6251 : _GEN_5585; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6260 = _T_189 ? _GEN_6252 : _GEN_5586; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6261 = _T_189 ? _GEN_6253 : _GEN_5587; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_6262 = io_op_bits_base_vs1_valid ? _GEN_6198 : _GEN_5540; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6263 = io_op_bits_base_vs1_valid ? _GEN_6199 : _GEN_5541; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6264 = io_op_bits_base_vs1_valid ? _GEN_6200 : _GEN_5542; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6265 = io_op_bits_base_vs1_valid ? _GEN_6201 : _GEN_5543; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6266 = io_op_bits_base_vs1_valid ? _GEN_6202 : _GEN_5544; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6267 = io_op_bits_base_vs1_valid ? _GEN_6203 : _GEN_5545; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6268 = io_op_bits_base_vs1_valid ? _GEN_6204 : _GEN_5546; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6269 = io_op_bits_base_vs1_valid ? _GEN_6205 : _GEN_5547; // @[sequencer-master.scala 328:47]
  wire  _GEN_6270 = io_op_bits_base_vs1_valid ? _GEN_6206 : _GEN_5726; // @[sequencer-master.scala 328:47]
  wire  _GEN_6271 = io_op_bits_base_vs1_valid ? _GEN_6207 : _GEN_5727; // @[sequencer-master.scala 328:47]
  wire  _GEN_6272 = io_op_bits_base_vs1_valid ? _GEN_6208 : _GEN_5728; // @[sequencer-master.scala 328:47]
  wire  _GEN_6273 = io_op_bits_base_vs1_valid ? _GEN_6209 : _GEN_5729; // @[sequencer-master.scala 328:47]
  wire  _GEN_6274 = io_op_bits_base_vs1_valid ? _GEN_6210 : _GEN_5730; // @[sequencer-master.scala 328:47]
  wire  _GEN_6275 = io_op_bits_base_vs1_valid ? _GEN_6211 : _GEN_5731; // @[sequencer-master.scala 328:47]
  wire  _GEN_6276 = io_op_bits_base_vs1_valid ? _GEN_6212 : _GEN_5732; // @[sequencer-master.scala 328:47]
  wire  _GEN_6277 = io_op_bits_base_vs1_valid ? _GEN_6213 : _GEN_5733; // @[sequencer-master.scala 328:47]
  wire  _GEN_6278 = io_op_bits_base_vs1_valid ? _GEN_6214 : _GEN_5548; // @[sequencer-master.scala 328:47]
  wire  _GEN_6279 = io_op_bits_base_vs1_valid ? _GEN_6215 : _GEN_5549; // @[sequencer-master.scala 328:47]
  wire  _GEN_6280 = io_op_bits_base_vs1_valid ? _GEN_6216 : _GEN_5550; // @[sequencer-master.scala 328:47]
  wire  _GEN_6281 = io_op_bits_base_vs1_valid ? _GEN_6217 : _GEN_5551; // @[sequencer-master.scala 328:47]
  wire  _GEN_6282 = io_op_bits_base_vs1_valid ? _GEN_6218 : _GEN_5552; // @[sequencer-master.scala 328:47]
  wire  _GEN_6283 = io_op_bits_base_vs1_valid ? _GEN_6219 : _GEN_5553; // @[sequencer-master.scala 328:47]
  wire  _GEN_6284 = io_op_bits_base_vs1_valid ? _GEN_6220 : _GEN_5554; // @[sequencer-master.scala 328:47]
  wire  _GEN_6285 = io_op_bits_base_vs1_valid ? _GEN_6221 : _GEN_5555; // @[sequencer-master.scala 328:47]
  wire  _GEN_6286 = io_op_bits_base_vs1_valid ? _GEN_6222 : _GEN_5556; // @[sequencer-master.scala 328:47]
  wire  _GEN_6287 = io_op_bits_base_vs1_valid ? _GEN_6223 : _GEN_5557; // @[sequencer-master.scala 328:47]
  wire  _GEN_6288 = io_op_bits_base_vs1_valid ? _GEN_6224 : _GEN_5558; // @[sequencer-master.scala 328:47]
  wire  _GEN_6289 = io_op_bits_base_vs1_valid ? _GEN_6225 : _GEN_5559; // @[sequencer-master.scala 328:47]
  wire  _GEN_6290 = io_op_bits_base_vs1_valid ? _GEN_6226 : _GEN_5560; // @[sequencer-master.scala 328:47]
  wire  _GEN_6291 = io_op_bits_base_vs1_valid ? _GEN_6227 : _GEN_5561; // @[sequencer-master.scala 328:47]
  wire  _GEN_6292 = io_op_bits_base_vs1_valid ? _GEN_6228 : _GEN_5562; // @[sequencer-master.scala 328:47]
  wire  _GEN_6293 = io_op_bits_base_vs1_valid ? _GEN_6229 : _GEN_5563; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6294 = io_op_bits_base_vs1_valid ? _GEN_6230 : _GEN_5564; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6295 = io_op_bits_base_vs1_valid ? _GEN_6231 : _GEN_5565; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6296 = io_op_bits_base_vs1_valid ? _GEN_6232 : _GEN_5566; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6297 = io_op_bits_base_vs1_valid ? _GEN_6233 : _GEN_5567; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6298 = io_op_bits_base_vs1_valid ? _GEN_6234 : _GEN_5568; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6299 = io_op_bits_base_vs1_valid ? _GEN_6235 : _GEN_5569; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6300 = io_op_bits_base_vs1_valid ? _GEN_6236 : _GEN_5570; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6301 = io_op_bits_base_vs1_valid ? _GEN_6237 : _GEN_5571; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6302 = io_op_bits_base_vs1_valid ? _GEN_6238 : _GEN_5572; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6303 = io_op_bits_base_vs1_valid ? _GEN_6239 : _GEN_5573; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6304 = io_op_bits_base_vs1_valid ? _GEN_6240 : _GEN_5574; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6305 = io_op_bits_base_vs1_valid ? _GEN_6241 : _GEN_5575; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6306 = io_op_bits_base_vs1_valid ? _GEN_6242 : _GEN_5576; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6307 = io_op_bits_base_vs1_valid ? _GEN_6243 : _GEN_5577; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6308 = io_op_bits_base_vs1_valid ? _GEN_6244 : _GEN_5578; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6309 = io_op_bits_base_vs1_valid ? _GEN_6245 : _GEN_5579; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6310 = io_op_bits_base_vs1_valid ? _GEN_6254 : _GEN_5580; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6311 = io_op_bits_base_vs1_valid ? _GEN_6255 : _GEN_5581; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6312 = io_op_bits_base_vs1_valid ? _GEN_6256 : _GEN_5582; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6313 = io_op_bits_base_vs1_valid ? _GEN_6257 : _GEN_5583; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6314 = io_op_bits_base_vs1_valid ? _GEN_6258 : _GEN_5584; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6315 = io_op_bits_base_vs1_valid ? _GEN_6259 : _GEN_5585; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6316 = io_op_bits_base_vs1_valid ? _GEN_6260 : _GEN_5586; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6317 = io_op_bits_base_vs1_valid ? _GEN_6261 : _GEN_5587; // @[sequencer-master.scala 328:47]
  wire  _GEN_6318 = _GEN_32729 | _GEN_6078; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6319 = _GEN_32730 | _GEN_6079; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6320 = _GEN_32731 | _GEN_6080; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6321 = _GEN_32732 | _GEN_6081; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6322 = _GEN_32733 | _GEN_6082; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6323 = _GEN_32734 | _GEN_6083; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6324 = _GEN_32735 | _GEN_6084; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6325 = _GEN_32736 | _GEN_6085; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6326 = _T_203 ? _GEN_6318 : _GEN_6078; // @[sequencer-master.scala 154:24]
  wire  _GEN_6327 = _T_203 ? _GEN_6319 : _GEN_6079; // @[sequencer-master.scala 154:24]
  wire  _GEN_6328 = _T_203 ? _GEN_6320 : _GEN_6080; // @[sequencer-master.scala 154:24]
  wire  _GEN_6329 = _T_203 ? _GEN_6321 : _GEN_6081; // @[sequencer-master.scala 154:24]
  wire  _GEN_6330 = _T_203 ? _GEN_6322 : _GEN_6082; // @[sequencer-master.scala 154:24]
  wire  _GEN_6331 = _T_203 ? _GEN_6323 : _GEN_6083; // @[sequencer-master.scala 154:24]
  wire  _GEN_6332 = _T_203 ? _GEN_6324 : _GEN_6084; // @[sequencer-master.scala 154:24]
  wire  _GEN_6333 = _T_203 ? _GEN_6325 : _GEN_6085; // @[sequencer-master.scala 154:24]
  wire  _GEN_6334 = _GEN_32729 | _GEN_6094; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6335 = _GEN_32730 | _GEN_6095; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6336 = _GEN_32731 | _GEN_6096; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6337 = _GEN_32732 | _GEN_6097; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6338 = _GEN_32733 | _GEN_6098; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6339 = _GEN_32734 | _GEN_6099; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6340 = _GEN_32735 | _GEN_6100; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6341 = _GEN_32736 | _GEN_6101; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6342 = _T_225 ? _GEN_6334 : _GEN_6094; // @[sequencer-master.scala 154:24]
  wire  _GEN_6343 = _T_225 ? _GEN_6335 : _GEN_6095; // @[sequencer-master.scala 154:24]
  wire  _GEN_6344 = _T_225 ? _GEN_6336 : _GEN_6096; // @[sequencer-master.scala 154:24]
  wire  _GEN_6345 = _T_225 ? _GEN_6337 : _GEN_6097; // @[sequencer-master.scala 154:24]
  wire  _GEN_6346 = _T_225 ? _GEN_6338 : _GEN_6098; // @[sequencer-master.scala 154:24]
  wire  _GEN_6347 = _T_225 ? _GEN_6339 : _GEN_6099; // @[sequencer-master.scala 154:24]
  wire  _GEN_6348 = _T_225 ? _GEN_6340 : _GEN_6100; // @[sequencer-master.scala 154:24]
  wire  _GEN_6349 = _T_225 ? _GEN_6341 : _GEN_6101; // @[sequencer-master.scala 154:24]
  wire  _GEN_6350 = _GEN_32729 | _GEN_6110; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6351 = _GEN_32730 | _GEN_6111; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6352 = _GEN_32731 | _GEN_6112; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6353 = _GEN_32732 | _GEN_6113; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6354 = _GEN_32733 | _GEN_6114; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6355 = _GEN_32734 | _GEN_6115; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6356 = _GEN_32735 | _GEN_6116; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6357 = _GEN_32736 | _GEN_6117; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6358 = _T_247 ? _GEN_6350 : _GEN_6110; // @[sequencer-master.scala 154:24]
  wire  _GEN_6359 = _T_247 ? _GEN_6351 : _GEN_6111; // @[sequencer-master.scala 154:24]
  wire  _GEN_6360 = _T_247 ? _GEN_6352 : _GEN_6112; // @[sequencer-master.scala 154:24]
  wire  _GEN_6361 = _T_247 ? _GEN_6353 : _GEN_6113; // @[sequencer-master.scala 154:24]
  wire  _GEN_6362 = _T_247 ? _GEN_6354 : _GEN_6114; // @[sequencer-master.scala 154:24]
  wire  _GEN_6363 = _T_247 ? _GEN_6355 : _GEN_6115; // @[sequencer-master.scala 154:24]
  wire  _GEN_6364 = _T_247 ? _GEN_6356 : _GEN_6116; // @[sequencer-master.scala 154:24]
  wire  _GEN_6365 = _T_247 ? _GEN_6357 : _GEN_6117; // @[sequencer-master.scala 154:24]
  wire  _GEN_6366 = _GEN_32729 | _GEN_6126; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6367 = _GEN_32730 | _GEN_6127; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6368 = _GEN_32731 | _GEN_6128; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6369 = _GEN_32732 | _GEN_6129; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6370 = _GEN_32733 | _GEN_6130; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6371 = _GEN_32734 | _GEN_6131; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6372 = _GEN_32735 | _GEN_6132; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6373 = _GEN_32736 | _GEN_6133; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6374 = _T_269 ? _GEN_6366 : _GEN_6126; // @[sequencer-master.scala 154:24]
  wire  _GEN_6375 = _T_269 ? _GEN_6367 : _GEN_6127; // @[sequencer-master.scala 154:24]
  wire  _GEN_6376 = _T_269 ? _GEN_6368 : _GEN_6128; // @[sequencer-master.scala 154:24]
  wire  _GEN_6377 = _T_269 ? _GEN_6369 : _GEN_6129; // @[sequencer-master.scala 154:24]
  wire  _GEN_6378 = _T_269 ? _GEN_6370 : _GEN_6130; // @[sequencer-master.scala 154:24]
  wire  _GEN_6379 = _T_269 ? _GEN_6371 : _GEN_6131; // @[sequencer-master.scala 154:24]
  wire  _GEN_6380 = _T_269 ? _GEN_6372 : _GEN_6132; // @[sequencer-master.scala 154:24]
  wire  _GEN_6381 = _T_269 ? _GEN_6373 : _GEN_6133; // @[sequencer-master.scala 154:24]
  wire  _GEN_6382 = _GEN_32729 | _GEN_6142; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6383 = _GEN_32730 | _GEN_6143; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6384 = _GEN_32731 | _GEN_6144; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6385 = _GEN_32732 | _GEN_6145; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6386 = _GEN_32733 | _GEN_6146; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6387 = _GEN_32734 | _GEN_6147; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6388 = _GEN_32735 | _GEN_6148; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6389 = _GEN_32736 | _GEN_6149; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6390 = _T_291 ? _GEN_6382 : _GEN_6142; // @[sequencer-master.scala 154:24]
  wire  _GEN_6391 = _T_291 ? _GEN_6383 : _GEN_6143; // @[sequencer-master.scala 154:24]
  wire  _GEN_6392 = _T_291 ? _GEN_6384 : _GEN_6144; // @[sequencer-master.scala 154:24]
  wire  _GEN_6393 = _T_291 ? _GEN_6385 : _GEN_6145; // @[sequencer-master.scala 154:24]
  wire  _GEN_6394 = _T_291 ? _GEN_6386 : _GEN_6146; // @[sequencer-master.scala 154:24]
  wire  _GEN_6395 = _T_291 ? _GEN_6387 : _GEN_6147; // @[sequencer-master.scala 154:24]
  wire  _GEN_6396 = _T_291 ? _GEN_6388 : _GEN_6148; // @[sequencer-master.scala 154:24]
  wire  _GEN_6397 = _T_291 ? _GEN_6389 : _GEN_6149; // @[sequencer-master.scala 154:24]
  wire  _GEN_6398 = _GEN_32729 | _GEN_6158; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6399 = _GEN_32730 | _GEN_6159; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6400 = _GEN_32731 | _GEN_6160; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6401 = _GEN_32732 | _GEN_6161; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6402 = _GEN_32733 | _GEN_6162; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6403 = _GEN_32734 | _GEN_6163; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6404 = _GEN_32735 | _GEN_6164; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6405 = _GEN_32736 | _GEN_6165; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6406 = _T_313 ? _GEN_6398 : _GEN_6158; // @[sequencer-master.scala 154:24]
  wire  _GEN_6407 = _T_313 ? _GEN_6399 : _GEN_6159; // @[sequencer-master.scala 154:24]
  wire  _GEN_6408 = _T_313 ? _GEN_6400 : _GEN_6160; // @[sequencer-master.scala 154:24]
  wire  _GEN_6409 = _T_313 ? _GEN_6401 : _GEN_6161; // @[sequencer-master.scala 154:24]
  wire  _GEN_6410 = _T_313 ? _GEN_6402 : _GEN_6162; // @[sequencer-master.scala 154:24]
  wire  _GEN_6411 = _T_313 ? _GEN_6403 : _GEN_6163; // @[sequencer-master.scala 154:24]
  wire  _GEN_6412 = _T_313 ? _GEN_6404 : _GEN_6164; // @[sequencer-master.scala 154:24]
  wire  _GEN_6413 = _T_313 ? _GEN_6405 : _GEN_6165; // @[sequencer-master.scala 154:24]
  wire  _GEN_6414 = _GEN_32729 | _GEN_6174; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6415 = _GEN_32730 | _GEN_6175; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6416 = _GEN_32731 | _GEN_6176; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6417 = _GEN_32732 | _GEN_6177; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6418 = _GEN_32733 | _GEN_6178; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6419 = _GEN_32734 | _GEN_6179; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6420 = _GEN_32735 | _GEN_6180; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6421 = _GEN_32736 | _GEN_6181; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6422 = _T_335 ? _GEN_6414 : _GEN_6174; // @[sequencer-master.scala 154:24]
  wire  _GEN_6423 = _T_335 ? _GEN_6415 : _GEN_6175; // @[sequencer-master.scala 154:24]
  wire  _GEN_6424 = _T_335 ? _GEN_6416 : _GEN_6176; // @[sequencer-master.scala 154:24]
  wire  _GEN_6425 = _T_335 ? _GEN_6417 : _GEN_6177; // @[sequencer-master.scala 154:24]
  wire  _GEN_6426 = _T_335 ? _GEN_6418 : _GEN_6178; // @[sequencer-master.scala 154:24]
  wire  _GEN_6427 = _T_335 ? _GEN_6419 : _GEN_6179; // @[sequencer-master.scala 154:24]
  wire  _GEN_6428 = _T_335 ? _GEN_6420 : _GEN_6180; // @[sequencer-master.scala 154:24]
  wire  _GEN_6429 = _T_335 ? _GEN_6421 : _GEN_6181; // @[sequencer-master.scala 154:24]
  wire  _GEN_6430 = _GEN_32729 | _GEN_6190; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6431 = _GEN_32730 | _GEN_6191; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6432 = _GEN_32731 | _GEN_6192; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6433 = _GEN_32732 | _GEN_6193; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6434 = _GEN_32733 | _GEN_6194; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6435 = _GEN_32734 | _GEN_6195; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6436 = _GEN_32735 | _GEN_6196; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6437 = _GEN_32736 | _GEN_6197; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6438 = _T_357 ? _GEN_6430 : _GEN_6190; // @[sequencer-master.scala 154:24]
  wire  _GEN_6439 = _T_357 ? _GEN_6431 : _GEN_6191; // @[sequencer-master.scala 154:24]
  wire  _GEN_6440 = _T_357 ? _GEN_6432 : _GEN_6192; // @[sequencer-master.scala 154:24]
  wire  _GEN_6441 = _T_357 ? _GEN_6433 : _GEN_6193; // @[sequencer-master.scala 154:24]
  wire  _GEN_6442 = _T_357 ? _GEN_6434 : _GEN_6194; // @[sequencer-master.scala 154:24]
  wire  _GEN_6443 = _T_357 ? _GEN_6435 : _GEN_6195; // @[sequencer-master.scala 154:24]
  wire  _GEN_6444 = _T_357 ? _GEN_6436 : _GEN_6196; // @[sequencer-master.scala 154:24]
  wire  _GEN_6445 = _T_357 ? _GEN_6437 : _GEN_6197; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_6446 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_5588; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6447 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_5589; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6448 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_5590; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6449 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_5591; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6450 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_5592; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6451 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_5593; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6452 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_5594; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6453 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_5595; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6454 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_5734; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6455 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_5735; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6456 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_5736; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6457 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_5737; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6458 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_5738; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6459 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_5739; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6460 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_5740; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6461 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_5741; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6462 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_5596; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6463 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_5597; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6464 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_5598; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6465 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_5599; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6466 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_5600; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6467 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_5601; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6468 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_5602; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6469 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_5603; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6470 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_5604; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6471 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_5605; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6472 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_5606; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6473 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_5607; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6474 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_5608; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6475 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_5609; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6476 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_5610; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_6477 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_5611; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6478 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_5612; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6479 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_5613; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6480 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_5614; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6481 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_5615; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6482 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_5616; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6483 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_5617; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6484 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_5618; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_6485 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_5619; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_6486 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_5620; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6487 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_5621; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6488 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_5622; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6489 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_5623; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6490 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_5624; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6491 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_5625; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6492 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_5626; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_6493 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_5627; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_6494 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_5628; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6495 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_5629; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6496 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_5630; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6497 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_5631; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6498 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_5632; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6499 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_5633; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6500 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_5634; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6501 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_5635; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_6502 = _T_366 ? _GEN_6494 : _GEN_5628; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6503 = _T_366 ? _GEN_6495 : _GEN_5629; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6504 = _T_366 ? _GEN_6496 : _GEN_5630; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6505 = _T_366 ? _GEN_6497 : _GEN_5631; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6506 = _T_366 ? _GEN_6498 : _GEN_5632; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6507 = _T_366 ? _GEN_6499 : _GEN_5633; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6508 = _T_366 ? _GEN_6500 : _GEN_5634; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_6509 = _T_366 ? _GEN_6501 : _GEN_5635; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_6510 = io_op_bits_base_vs2_valid ? _GEN_6446 : _GEN_5588; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6511 = io_op_bits_base_vs2_valid ? _GEN_6447 : _GEN_5589; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6512 = io_op_bits_base_vs2_valid ? _GEN_6448 : _GEN_5590; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6513 = io_op_bits_base_vs2_valid ? _GEN_6449 : _GEN_5591; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6514 = io_op_bits_base_vs2_valid ? _GEN_6450 : _GEN_5592; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6515 = io_op_bits_base_vs2_valid ? _GEN_6451 : _GEN_5593; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6516 = io_op_bits_base_vs2_valid ? _GEN_6452 : _GEN_5594; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6517 = io_op_bits_base_vs2_valid ? _GEN_6453 : _GEN_5595; // @[sequencer-master.scala 328:47]
  wire  _GEN_6518 = io_op_bits_base_vs2_valid ? _GEN_6454 : _GEN_5734; // @[sequencer-master.scala 328:47]
  wire  _GEN_6519 = io_op_bits_base_vs2_valid ? _GEN_6455 : _GEN_5735; // @[sequencer-master.scala 328:47]
  wire  _GEN_6520 = io_op_bits_base_vs2_valid ? _GEN_6456 : _GEN_5736; // @[sequencer-master.scala 328:47]
  wire  _GEN_6521 = io_op_bits_base_vs2_valid ? _GEN_6457 : _GEN_5737; // @[sequencer-master.scala 328:47]
  wire  _GEN_6522 = io_op_bits_base_vs2_valid ? _GEN_6458 : _GEN_5738; // @[sequencer-master.scala 328:47]
  wire  _GEN_6523 = io_op_bits_base_vs2_valid ? _GEN_6459 : _GEN_5739; // @[sequencer-master.scala 328:47]
  wire  _GEN_6524 = io_op_bits_base_vs2_valid ? _GEN_6460 : _GEN_5740; // @[sequencer-master.scala 328:47]
  wire  _GEN_6525 = io_op_bits_base_vs2_valid ? _GEN_6461 : _GEN_5741; // @[sequencer-master.scala 328:47]
  wire  _GEN_6526 = io_op_bits_base_vs2_valid ? _GEN_6462 : _GEN_5596; // @[sequencer-master.scala 328:47]
  wire  _GEN_6527 = io_op_bits_base_vs2_valid ? _GEN_6463 : _GEN_5597; // @[sequencer-master.scala 328:47]
  wire  _GEN_6528 = io_op_bits_base_vs2_valid ? _GEN_6464 : _GEN_5598; // @[sequencer-master.scala 328:47]
  wire  _GEN_6529 = io_op_bits_base_vs2_valid ? _GEN_6465 : _GEN_5599; // @[sequencer-master.scala 328:47]
  wire  _GEN_6530 = io_op_bits_base_vs2_valid ? _GEN_6466 : _GEN_5600; // @[sequencer-master.scala 328:47]
  wire  _GEN_6531 = io_op_bits_base_vs2_valid ? _GEN_6467 : _GEN_5601; // @[sequencer-master.scala 328:47]
  wire  _GEN_6532 = io_op_bits_base_vs2_valid ? _GEN_6468 : _GEN_5602; // @[sequencer-master.scala 328:47]
  wire  _GEN_6533 = io_op_bits_base_vs2_valid ? _GEN_6469 : _GEN_5603; // @[sequencer-master.scala 328:47]
  wire  _GEN_6534 = io_op_bits_base_vs2_valid ? _GEN_6470 : _GEN_5604; // @[sequencer-master.scala 328:47]
  wire  _GEN_6535 = io_op_bits_base_vs2_valid ? _GEN_6471 : _GEN_5605; // @[sequencer-master.scala 328:47]
  wire  _GEN_6536 = io_op_bits_base_vs2_valid ? _GEN_6472 : _GEN_5606; // @[sequencer-master.scala 328:47]
  wire  _GEN_6537 = io_op_bits_base_vs2_valid ? _GEN_6473 : _GEN_5607; // @[sequencer-master.scala 328:47]
  wire  _GEN_6538 = io_op_bits_base_vs2_valid ? _GEN_6474 : _GEN_5608; // @[sequencer-master.scala 328:47]
  wire  _GEN_6539 = io_op_bits_base_vs2_valid ? _GEN_6475 : _GEN_5609; // @[sequencer-master.scala 328:47]
  wire  _GEN_6540 = io_op_bits_base_vs2_valid ? _GEN_6476 : _GEN_5610; // @[sequencer-master.scala 328:47]
  wire  _GEN_6541 = io_op_bits_base_vs2_valid ? _GEN_6477 : _GEN_5611; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6542 = io_op_bits_base_vs2_valid ? _GEN_6478 : _GEN_5612; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6543 = io_op_bits_base_vs2_valid ? _GEN_6479 : _GEN_5613; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6544 = io_op_bits_base_vs2_valid ? _GEN_6480 : _GEN_5614; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6545 = io_op_bits_base_vs2_valid ? _GEN_6481 : _GEN_5615; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6546 = io_op_bits_base_vs2_valid ? _GEN_6482 : _GEN_5616; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6547 = io_op_bits_base_vs2_valid ? _GEN_6483 : _GEN_5617; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6548 = io_op_bits_base_vs2_valid ? _GEN_6484 : _GEN_5618; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_6549 = io_op_bits_base_vs2_valid ? _GEN_6485 : _GEN_5619; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6550 = io_op_bits_base_vs2_valid ? _GEN_6486 : _GEN_5620; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6551 = io_op_bits_base_vs2_valid ? _GEN_6487 : _GEN_5621; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6552 = io_op_bits_base_vs2_valid ? _GEN_6488 : _GEN_5622; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6553 = io_op_bits_base_vs2_valid ? _GEN_6489 : _GEN_5623; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6554 = io_op_bits_base_vs2_valid ? _GEN_6490 : _GEN_5624; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6555 = io_op_bits_base_vs2_valid ? _GEN_6491 : _GEN_5625; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6556 = io_op_bits_base_vs2_valid ? _GEN_6492 : _GEN_5626; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_6557 = io_op_bits_base_vs2_valid ? _GEN_6493 : _GEN_5627; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6558 = io_op_bits_base_vs2_valid ? _GEN_6502 : _GEN_5628; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6559 = io_op_bits_base_vs2_valid ? _GEN_6503 : _GEN_5629; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6560 = io_op_bits_base_vs2_valid ? _GEN_6504 : _GEN_5630; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6561 = io_op_bits_base_vs2_valid ? _GEN_6505 : _GEN_5631; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6562 = io_op_bits_base_vs2_valid ? _GEN_6506 : _GEN_5632; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6563 = io_op_bits_base_vs2_valid ? _GEN_6507 : _GEN_5633; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6564 = io_op_bits_base_vs2_valid ? _GEN_6508 : _GEN_5634; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_6565 = io_op_bits_base_vs2_valid ? _GEN_6509 : _GEN_5635; // @[sequencer-master.scala 328:47]
  wire  _GEN_6566 = _GEN_32729 | _GEN_6326; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6567 = _GEN_32730 | _GEN_6327; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6568 = _GEN_32731 | _GEN_6328; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6569 = _GEN_32732 | _GEN_6329; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6570 = _GEN_32733 | _GEN_6330; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6571 = _GEN_32734 | _GEN_6331; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6572 = _GEN_32735 | _GEN_6332; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6573 = _GEN_32736 | _GEN_6333; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6574 = _T_380 ? _GEN_6566 : _GEN_6326; // @[sequencer-master.scala 154:24]
  wire  _GEN_6575 = _T_380 ? _GEN_6567 : _GEN_6327; // @[sequencer-master.scala 154:24]
  wire  _GEN_6576 = _T_380 ? _GEN_6568 : _GEN_6328; // @[sequencer-master.scala 154:24]
  wire  _GEN_6577 = _T_380 ? _GEN_6569 : _GEN_6329; // @[sequencer-master.scala 154:24]
  wire  _GEN_6578 = _T_380 ? _GEN_6570 : _GEN_6330; // @[sequencer-master.scala 154:24]
  wire  _GEN_6579 = _T_380 ? _GEN_6571 : _GEN_6331; // @[sequencer-master.scala 154:24]
  wire  _GEN_6580 = _T_380 ? _GEN_6572 : _GEN_6332; // @[sequencer-master.scala 154:24]
  wire  _GEN_6581 = _T_380 ? _GEN_6573 : _GEN_6333; // @[sequencer-master.scala 154:24]
  wire  _GEN_6582 = _GEN_32729 | _GEN_6342; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6583 = _GEN_32730 | _GEN_6343; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6584 = _GEN_32731 | _GEN_6344; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6585 = _GEN_32732 | _GEN_6345; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6586 = _GEN_32733 | _GEN_6346; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6587 = _GEN_32734 | _GEN_6347; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6588 = _GEN_32735 | _GEN_6348; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6589 = _GEN_32736 | _GEN_6349; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6590 = _T_402 ? _GEN_6582 : _GEN_6342; // @[sequencer-master.scala 154:24]
  wire  _GEN_6591 = _T_402 ? _GEN_6583 : _GEN_6343; // @[sequencer-master.scala 154:24]
  wire  _GEN_6592 = _T_402 ? _GEN_6584 : _GEN_6344; // @[sequencer-master.scala 154:24]
  wire  _GEN_6593 = _T_402 ? _GEN_6585 : _GEN_6345; // @[sequencer-master.scala 154:24]
  wire  _GEN_6594 = _T_402 ? _GEN_6586 : _GEN_6346; // @[sequencer-master.scala 154:24]
  wire  _GEN_6595 = _T_402 ? _GEN_6587 : _GEN_6347; // @[sequencer-master.scala 154:24]
  wire  _GEN_6596 = _T_402 ? _GEN_6588 : _GEN_6348; // @[sequencer-master.scala 154:24]
  wire  _GEN_6597 = _T_402 ? _GEN_6589 : _GEN_6349; // @[sequencer-master.scala 154:24]
  wire  _GEN_6598 = _GEN_32729 | _GEN_6358; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6599 = _GEN_32730 | _GEN_6359; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6600 = _GEN_32731 | _GEN_6360; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6601 = _GEN_32732 | _GEN_6361; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6602 = _GEN_32733 | _GEN_6362; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6603 = _GEN_32734 | _GEN_6363; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6604 = _GEN_32735 | _GEN_6364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6605 = _GEN_32736 | _GEN_6365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6606 = _T_424 ? _GEN_6598 : _GEN_6358; // @[sequencer-master.scala 154:24]
  wire  _GEN_6607 = _T_424 ? _GEN_6599 : _GEN_6359; // @[sequencer-master.scala 154:24]
  wire  _GEN_6608 = _T_424 ? _GEN_6600 : _GEN_6360; // @[sequencer-master.scala 154:24]
  wire  _GEN_6609 = _T_424 ? _GEN_6601 : _GEN_6361; // @[sequencer-master.scala 154:24]
  wire  _GEN_6610 = _T_424 ? _GEN_6602 : _GEN_6362; // @[sequencer-master.scala 154:24]
  wire  _GEN_6611 = _T_424 ? _GEN_6603 : _GEN_6363; // @[sequencer-master.scala 154:24]
  wire  _GEN_6612 = _T_424 ? _GEN_6604 : _GEN_6364; // @[sequencer-master.scala 154:24]
  wire  _GEN_6613 = _T_424 ? _GEN_6605 : _GEN_6365; // @[sequencer-master.scala 154:24]
  wire  _GEN_6614 = _GEN_32729 | _GEN_6374; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6615 = _GEN_32730 | _GEN_6375; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6616 = _GEN_32731 | _GEN_6376; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6617 = _GEN_32732 | _GEN_6377; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6618 = _GEN_32733 | _GEN_6378; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6619 = _GEN_32734 | _GEN_6379; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6620 = _GEN_32735 | _GEN_6380; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6621 = _GEN_32736 | _GEN_6381; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6622 = _T_446 ? _GEN_6614 : _GEN_6374; // @[sequencer-master.scala 154:24]
  wire  _GEN_6623 = _T_446 ? _GEN_6615 : _GEN_6375; // @[sequencer-master.scala 154:24]
  wire  _GEN_6624 = _T_446 ? _GEN_6616 : _GEN_6376; // @[sequencer-master.scala 154:24]
  wire  _GEN_6625 = _T_446 ? _GEN_6617 : _GEN_6377; // @[sequencer-master.scala 154:24]
  wire  _GEN_6626 = _T_446 ? _GEN_6618 : _GEN_6378; // @[sequencer-master.scala 154:24]
  wire  _GEN_6627 = _T_446 ? _GEN_6619 : _GEN_6379; // @[sequencer-master.scala 154:24]
  wire  _GEN_6628 = _T_446 ? _GEN_6620 : _GEN_6380; // @[sequencer-master.scala 154:24]
  wire  _GEN_6629 = _T_446 ? _GEN_6621 : _GEN_6381; // @[sequencer-master.scala 154:24]
  wire  _GEN_6630 = _GEN_32729 | _GEN_6390; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6631 = _GEN_32730 | _GEN_6391; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6632 = _GEN_32731 | _GEN_6392; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6633 = _GEN_32732 | _GEN_6393; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6634 = _GEN_32733 | _GEN_6394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6635 = _GEN_32734 | _GEN_6395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6636 = _GEN_32735 | _GEN_6396; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6637 = _GEN_32736 | _GEN_6397; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6638 = _T_468 ? _GEN_6630 : _GEN_6390; // @[sequencer-master.scala 154:24]
  wire  _GEN_6639 = _T_468 ? _GEN_6631 : _GEN_6391; // @[sequencer-master.scala 154:24]
  wire  _GEN_6640 = _T_468 ? _GEN_6632 : _GEN_6392; // @[sequencer-master.scala 154:24]
  wire  _GEN_6641 = _T_468 ? _GEN_6633 : _GEN_6393; // @[sequencer-master.scala 154:24]
  wire  _GEN_6642 = _T_468 ? _GEN_6634 : _GEN_6394; // @[sequencer-master.scala 154:24]
  wire  _GEN_6643 = _T_468 ? _GEN_6635 : _GEN_6395; // @[sequencer-master.scala 154:24]
  wire  _GEN_6644 = _T_468 ? _GEN_6636 : _GEN_6396; // @[sequencer-master.scala 154:24]
  wire  _GEN_6645 = _T_468 ? _GEN_6637 : _GEN_6397; // @[sequencer-master.scala 154:24]
  wire  _GEN_6646 = _GEN_32729 | _GEN_6406; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6647 = _GEN_32730 | _GEN_6407; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6648 = _GEN_32731 | _GEN_6408; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6649 = _GEN_32732 | _GEN_6409; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6650 = _GEN_32733 | _GEN_6410; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6651 = _GEN_32734 | _GEN_6411; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6652 = _GEN_32735 | _GEN_6412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6653 = _GEN_32736 | _GEN_6413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6654 = _T_490 ? _GEN_6646 : _GEN_6406; // @[sequencer-master.scala 154:24]
  wire  _GEN_6655 = _T_490 ? _GEN_6647 : _GEN_6407; // @[sequencer-master.scala 154:24]
  wire  _GEN_6656 = _T_490 ? _GEN_6648 : _GEN_6408; // @[sequencer-master.scala 154:24]
  wire  _GEN_6657 = _T_490 ? _GEN_6649 : _GEN_6409; // @[sequencer-master.scala 154:24]
  wire  _GEN_6658 = _T_490 ? _GEN_6650 : _GEN_6410; // @[sequencer-master.scala 154:24]
  wire  _GEN_6659 = _T_490 ? _GEN_6651 : _GEN_6411; // @[sequencer-master.scala 154:24]
  wire  _GEN_6660 = _T_490 ? _GEN_6652 : _GEN_6412; // @[sequencer-master.scala 154:24]
  wire  _GEN_6661 = _T_490 ? _GEN_6653 : _GEN_6413; // @[sequencer-master.scala 154:24]
  wire  _GEN_6662 = _GEN_32729 | _GEN_6422; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6663 = _GEN_32730 | _GEN_6423; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6664 = _GEN_32731 | _GEN_6424; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6665 = _GEN_32732 | _GEN_6425; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6666 = _GEN_32733 | _GEN_6426; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6667 = _GEN_32734 | _GEN_6427; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6668 = _GEN_32735 | _GEN_6428; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6669 = _GEN_32736 | _GEN_6429; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6670 = _T_512 ? _GEN_6662 : _GEN_6422; // @[sequencer-master.scala 154:24]
  wire  _GEN_6671 = _T_512 ? _GEN_6663 : _GEN_6423; // @[sequencer-master.scala 154:24]
  wire  _GEN_6672 = _T_512 ? _GEN_6664 : _GEN_6424; // @[sequencer-master.scala 154:24]
  wire  _GEN_6673 = _T_512 ? _GEN_6665 : _GEN_6425; // @[sequencer-master.scala 154:24]
  wire  _GEN_6674 = _T_512 ? _GEN_6666 : _GEN_6426; // @[sequencer-master.scala 154:24]
  wire  _GEN_6675 = _T_512 ? _GEN_6667 : _GEN_6427; // @[sequencer-master.scala 154:24]
  wire  _GEN_6676 = _T_512 ? _GEN_6668 : _GEN_6428; // @[sequencer-master.scala 154:24]
  wire  _GEN_6677 = _T_512 ? _GEN_6669 : _GEN_6429; // @[sequencer-master.scala 154:24]
  wire  _GEN_6678 = _GEN_32729 | _GEN_6438; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6679 = _GEN_32730 | _GEN_6439; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6680 = _GEN_32731 | _GEN_6440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6681 = _GEN_32732 | _GEN_6441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6682 = _GEN_32733 | _GEN_6442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6683 = _GEN_32734 | _GEN_6443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6684 = _GEN_32735 | _GEN_6444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6685 = _GEN_32736 | _GEN_6445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_6686 = _T_534 ? _GEN_6678 : _GEN_6438; // @[sequencer-master.scala 154:24]
  wire  _GEN_6687 = _T_534 ? _GEN_6679 : _GEN_6439; // @[sequencer-master.scala 154:24]
  wire  _GEN_6688 = _T_534 ? _GEN_6680 : _GEN_6440; // @[sequencer-master.scala 154:24]
  wire  _GEN_6689 = _T_534 ? _GEN_6681 : _GEN_6441; // @[sequencer-master.scala 154:24]
  wire  _GEN_6690 = _T_534 ? _GEN_6682 : _GEN_6442; // @[sequencer-master.scala 154:24]
  wire  _GEN_6691 = _T_534 ? _GEN_6683 : _GEN_6443; // @[sequencer-master.scala 154:24]
  wire  _GEN_6692 = _T_534 ? _GEN_6684 : _GEN_6444; // @[sequencer-master.scala 154:24]
  wire  _GEN_6693 = _T_534 ? _GEN_6685 : _GEN_6445; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_6694 = 3'h0 == tail ? _T_1615[1:0] : _GEN_5676; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6695 = 3'h1 == tail ? _T_1615[1:0] : _GEN_5677; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6696 = 3'h2 == tail ? _T_1615[1:0] : _GEN_5678; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6697 = 3'h3 == tail ? _T_1615[1:0] : _GEN_5679; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6698 = 3'h4 == tail ? _T_1615[1:0] : _GEN_5680; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6699 = 3'h5 == tail ? _T_1615[1:0] : _GEN_5681; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6700 = 3'h6 == tail ? _T_1615[1:0] : _GEN_5682; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_6701 = 3'h7 == tail ? _T_1615[1:0] : _GEN_5683; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_6702 = 3'h0 == tail ? 4'h0 : _GEN_5684; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6703 = 3'h1 == tail ? 4'h0 : _GEN_5685; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6704 = 3'h2 == tail ? 4'h0 : _GEN_5686; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6705 = 3'h3 == tail ? 4'h0 : _GEN_5687; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6706 = 3'h4 == tail ? 4'h0 : _GEN_5688; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6707 = 3'h5 == tail ? 4'h0 : _GEN_5689; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6708 = 3'h6 == tail ? 4'h0 : _GEN_5690; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_6709 = 3'h7 == tail ? 4'h0 : _GEN_5691; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_6710 = 3'h0 == tail ? 3'h0 : _GEN_5692; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6711 = 3'h1 == tail ? 3'h0 : _GEN_5693; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6712 = 3'h2 == tail ? 3'h0 : _GEN_5694; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6713 = 3'h3 == tail ? 3'h0 : _GEN_5695; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6714 = 3'h4 == tail ? 3'h0 : _GEN_5696; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6715 = 3'h5 == tail ? 3'h0 : _GEN_5697; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6716 = 3'h6 == tail ? 3'h0 : _GEN_5698; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_6717 = 3'h7 == tail ? 3'h0 : _GEN_5699; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_6718 = _GEN_32729 | _GEN_5774; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6719 = _GEN_32730 | _GEN_5775; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6720 = _GEN_32731 | _GEN_5776; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6721 = _GEN_32732 | _GEN_5777; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6722 = _GEN_32733 | _GEN_5778; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6723 = _GEN_32734 | _GEN_5779; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6724 = _GEN_32735 | _GEN_5780; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6725 = _GEN_32736 | _GEN_5781; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6726 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6718 : _GEN_5774; // @[sequencer-master.scala 161:86]
  wire  _GEN_6727 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6719 : _GEN_5775; // @[sequencer-master.scala 161:86]
  wire  _GEN_6728 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6720 : _GEN_5776; // @[sequencer-master.scala 161:86]
  wire  _GEN_6729 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6721 : _GEN_5777; // @[sequencer-master.scala 161:86]
  wire  _GEN_6730 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6722 : _GEN_5778; // @[sequencer-master.scala 161:86]
  wire  _GEN_6731 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6723 : _GEN_5779; // @[sequencer-master.scala 161:86]
  wire  _GEN_6732 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6724 : _GEN_5780; // @[sequencer-master.scala 161:86]
  wire  _GEN_6733 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_6725 : _GEN_5781; // @[sequencer-master.scala 161:86]
  wire  _GEN_6734 = _GEN_32729 | _GEN_5798; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6735 = _GEN_32730 | _GEN_5799; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6736 = _GEN_32731 | _GEN_5800; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6737 = _GEN_32732 | _GEN_5801; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6738 = _GEN_32733 | _GEN_5802; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6739 = _GEN_32734 | _GEN_5803; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6740 = _GEN_32735 | _GEN_5804; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6741 = _GEN_32736 | _GEN_5805; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6742 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6734 : _GEN_5798; // @[sequencer-master.scala 161:86]
  wire  _GEN_6743 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6735 : _GEN_5799; // @[sequencer-master.scala 161:86]
  wire  _GEN_6744 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6736 : _GEN_5800; // @[sequencer-master.scala 161:86]
  wire  _GEN_6745 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6737 : _GEN_5801; // @[sequencer-master.scala 161:86]
  wire  _GEN_6746 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6738 : _GEN_5802; // @[sequencer-master.scala 161:86]
  wire  _GEN_6747 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6739 : _GEN_5803; // @[sequencer-master.scala 161:86]
  wire  _GEN_6748 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6740 : _GEN_5804; // @[sequencer-master.scala 161:86]
  wire  _GEN_6749 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_6741 : _GEN_5805; // @[sequencer-master.scala 161:86]
  wire  _GEN_6750 = _GEN_32729 | _GEN_5822; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6751 = _GEN_32730 | _GEN_5823; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6752 = _GEN_32731 | _GEN_5824; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6753 = _GEN_32732 | _GEN_5825; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6754 = _GEN_32733 | _GEN_5826; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6755 = _GEN_32734 | _GEN_5827; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6756 = _GEN_32735 | _GEN_5828; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6757 = _GEN_32736 | _GEN_5829; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6758 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6750 : _GEN_5822; // @[sequencer-master.scala 161:86]
  wire  _GEN_6759 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6751 : _GEN_5823; // @[sequencer-master.scala 161:86]
  wire  _GEN_6760 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6752 : _GEN_5824; // @[sequencer-master.scala 161:86]
  wire  _GEN_6761 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6753 : _GEN_5825; // @[sequencer-master.scala 161:86]
  wire  _GEN_6762 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6754 : _GEN_5826; // @[sequencer-master.scala 161:86]
  wire  _GEN_6763 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6755 : _GEN_5827; // @[sequencer-master.scala 161:86]
  wire  _GEN_6764 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6756 : _GEN_5828; // @[sequencer-master.scala 161:86]
  wire  _GEN_6765 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_6757 : _GEN_5829; // @[sequencer-master.scala 161:86]
  wire  _GEN_6766 = _GEN_32729 | _GEN_5846; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6767 = _GEN_32730 | _GEN_5847; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6768 = _GEN_32731 | _GEN_5848; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6769 = _GEN_32732 | _GEN_5849; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6770 = _GEN_32733 | _GEN_5850; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6771 = _GEN_32734 | _GEN_5851; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6772 = _GEN_32735 | _GEN_5852; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6773 = _GEN_32736 | _GEN_5853; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6774 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6766 : _GEN_5846; // @[sequencer-master.scala 161:86]
  wire  _GEN_6775 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6767 : _GEN_5847; // @[sequencer-master.scala 161:86]
  wire  _GEN_6776 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6768 : _GEN_5848; // @[sequencer-master.scala 161:86]
  wire  _GEN_6777 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6769 : _GEN_5849; // @[sequencer-master.scala 161:86]
  wire  _GEN_6778 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6770 : _GEN_5850; // @[sequencer-master.scala 161:86]
  wire  _GEN_6779 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6771 : _GEN_5851; // @[sequencer-master.scala 161:86]
  wire  _GEN_6780 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6772 : _GEN_5852; // @[sequencer-master.scala 161:86]
  wire  _GEN_6781 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_6773 : _GEN_5853; // @[sequencer-master.scala 161:86]
  wire  _GEN_6782 = _GEN_32729 | _GEN_5870; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6783 = _GEN_32730 | _GEN_5871; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6784 = _GEN_32731 | _GEN_5872; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6785 = _GEN_32732 | _GEN_5873; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6786 = _GEN_32733 | _GEN_5874; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6787 = _GEN_32734 | _GEN_5875; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6788 = _GEN_32735 | _GEN_5876; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6789 = _GEN_32736 | _GEN_5877; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6790 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6782 : _GEN_5870; // @[sequencer-master.scala 161:86]
  wire  _GEN_6791 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6783 : _GEN_5871; // @[sequencer-master.scala 161:86]
  wire  _GEN_6792 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6784 : _GEN_5872; // @[sequencer-master.scala 161:86]
  wire  _GEN_6793 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6785 : _GEN_5873; // @[sequencer-master.scala 161:86]
  wire  _GEN_6794 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6786 : _GEN_5874; // @[sequencer-master.scala 161:86]
  wire  _GEN_6795 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6787 : _GEN_5875; // @[sequencer-master.scala 161:86]
  wire  _GEN_6796 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6788 : _GEN_5876; // @[sequencer-master.scala 161:86]
  wire  _GEN_6797 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_6789 : _GEN_5877; // @[sequencer-master.scala 161:86]
  wire  _GEN_6798 = _GEN_32729 | _GEN_5894; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6799 = _GEN_32730 | _GEN_5895; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6800 = _GEN_32731 | _GEN_5896; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6801 = _GEN_32732 | _GEN_5897; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6802 = _GEN_32733 | _GEN_5898; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6803 = _GEN_32734 | _GEN_5899; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6804 = _GEN_32735 | _GEN_5900; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6805 = _GEN_32736 | _GEN_5901; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6806 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6798 : _GEN_5894; // @[sequencer-master.scala 161:86]
  wire  _GEN_6807 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6799 : _GEN_5895; // @[sequencer-master.scala 161:86]
  wire  _GEN_6808 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6800 : _GEN_5896; // @[sequencer-master.scala 161:86]
  wire  _GEN_6809 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6801 : _GEN_5897; // @[sequencer-master.scala 161:86]
  wire  _GEN_6810 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6802 : _GEN_5898; // @[sequencer-master.scala 161:86]
  wire  _GEN_6811 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6803 : _GEN_5899; // @[sequencer-master.scala 161:86]
  wire  _GEN_6812 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6804 : _GEN_5900; // @[sequencer-master.scala 161:86]
  wire  _GEN_6813 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_6805 : _GEN_5901; // @[sequencer-master.scala 161:86]
  wire  _GEN_6814 = _GEN_32729 | _GEN_5918; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6815 = _GEN_32730 | _GEN_5919; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6816 = _GEN_32731 | _GEN_5920; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6817 = _GEN_32732 | _GEN_5921; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6818 = _GEN_32733 | _GEN_5922; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6819 = _GEN_32734 | _GEN_5923; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6820 = _GEN_32735 | _GEN_5924; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6821 = _GEN_32736 | _GEN_5925; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6822 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6814 : _GEN_5918; // @[sequencer-master.scala 161:86]
  wire  _GEN_6823 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6815 : _GEN_5919; // @[sequencer-master.scala 161:86]
  wire  _GEN_6824 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6816 : _GEN_5920; // @[sequencer-master.scala 161:86]
  wire  _GEN_6825 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6817 : _GEN_5921; // @[sequencer-master.scala 161:86]
  wire  _GEN_6826 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6818 : _GEN_5922; // @[sequencer-master.scala 161:86]
  wire  _GEN_6827 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6819 : _GEN_5923; // @[sequencer-master.scala 161:86]
  wire  _GEN_6828 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6820 : _GEN_5924; // @[sequencer-master.scala 161:86]
  wire  _GEN_6829 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_6821 : _GEN_5925; // @[sequencer-master.scala 161:86]
  wire  _GEN_6830 = _GEN_32729 | _GEN_5942; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6831 = _GEN_32730 | _GEN_5943; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6832 = _GEN_32731 | _GEN_5944; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6833 = _GEN_32732 | _GEN_5945; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6834 = _GEN_32733 | _GEN_5946; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6835 = _GEN_32734 | _GEN_5947; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6836 = _GEN_32735 | _GEN_5948; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6837 = _GEN_32736 | _GEN_5949; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_6838 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6830 : _GEN_5942; // @[sequencer-master.scala 161:86]
  wire  _GEN_6839 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6831 : _GEN_5943; // @[sequencer-master.scala 161:86]
  wire  _GEN_6840 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6832 : _GEN_5944; // @[sequencer-master.scala 161:86]
  wire  _GEN_6841 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6833 : _GEN_5945; // @[sequencer-master.scala 161:86]
  wire  _GEN_6842 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6834 : _GEN_5946; // @[sequencer-master.scala 161:86]
  wire  _GEN_6843 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6835 : _GEN_5947; // @[sequencer-master.scala 161:86]
  wire  _GEN_6844 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6836 : _GEN_5948; // @[sequencer-master.scala 161:86]
  wire  _GEN_6845 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_6837 : _GEN_5949; // @[sequencer-master.scala 161:86]
  wire  _GEN_6846 = _GEN_32729 | _GEN_5782; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6847 = _GEN_32730 | _GEN_5783; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6848 = _GEN_32731 | _GEN_5784; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6849 = _GEN_32732 | _GEN_5785; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6850 = _GEN_32733 | _GEN_5786; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6851 = _GEN_32734 | _GEN_5787; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6852 = _GEN_32735 | _GEN_5788; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6853 = _GEN_32736 | _GEN_5789; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6854 = _T_1442 ? _GEN_6846 : _GEN_5782; // @[sequencer-master.scala 168:32]
  wire  _GEN_6855 = _T_1442 ? _GEN_6847 : _GEN_5783; // @[sequencer-master.scala 168:32]
  wire  _GEN_6856 = _T_1442 ? _GEN_6848 : _GEN_5784; // @[sequencer-master.scala 168:32]
  wire  _GEN_6857 = _T_1442 ? _GEN_6849 : _GEN_5785; // @[sequencer-master.scala 168:32]
  wire  _GEN_6858 = _T_1442 ? _GEN_6850 : _GEN_5786; // @[sequencer-master.scala 168:32]
  wire  _GEN_6859 = _T_1442 ? _GEN_6851 : _GEN_5787; // @[sequencer-master.scala 168:32]
  wire  _GEN_6860 = _T_1442 ? _GEN_6852 : _GEN_5788; // @[sequencer-master.scala 168:32]
  wire  _GEN_6861 = _T_1442 ? _GEN_6853 : _GEN_5789; // @[sequencer-master.scala 168:32]
  wire  _GEN_6862 = _GEN_32729 | _GEN_5806; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6863 = _GEN_32730 | _GEN_5807; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6864 = _GEN_32731 | _GEN_5808; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6865 = _GEN_32732 | _GEN_5809; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6866 = _GEN_32733 | _GEN_5810; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6867 = _GEN_32734 | _GEN_5811; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6868 = _GEN_32735 | _GEN_5812; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6869 = _GEN_32736 | _GEN_5813; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6870 = _T_1464 ? _GEN_6862 : _GEN_5806; // @[sequencer-master.scala 168:32]
  wire  _GEN_6871 = _T_1464 ? _GEN_6863 : _GEN_5807; // @[sequencer-master.scala 168:32]
  wire  _GEN_6872 = _T_1464 ? _GEN_6864 : _GEN_5808; // @[sequencer-master.scala 168:32]
  wire  _GEN_6873 = _T_1464 ? _GEN_6865 : _GEN_5809; // @[sequencer-master.scala 168:32]
  wire  _GEN_6874 = _T_1464 ? _GEN_6866 : _GEN_5810; // @[sequencer-master.scala 168:32]
  wire  _GEN_6875 = _T_1464 ? _GEN_6867 : _GEN_5811; // @[sequencer-master.scala 168:32]
  wire  _GEN_6876 = _T_1464 ? _GEN_6868 : _GEN_5812; // @[sequencer-master.scala 168:32]
  wire  _GEN_6877 = _T_1464 ? _GEN_6869 : _GEN_5813; // @[sequencer-master.scala 168:32]
  wire  _GEN_6878 = _GEN_32729 | _GEN_5830; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6879 = _GEN_32730 | _GEN_5831; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6880 = _GEN_32731 | _GEN_5832; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6881 = _GEN_32732 | _GEN_5833; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6882 = _GEN_32733 | _GEN_5834; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6883 = _GEN_32734 | _GEN_5835; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6884 = _GEN_32735 | _GEN_5836; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6885 = _GEN_32736 | _GEN_5837; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6886 = _T_1486 ? _GEN_6878 : _GEN_5830; // @[sequencer-master.scala 168:32]
  wire  _GEN_6887 = _T_1486 ? _GEN_6879 : _GEN_5831; // @[sequencer-master.scala 168:32]
  wire  _GEN_6888 = _T_1486 ? _GEN_6880 : _GEN_5832; // @[sequencer-master.scala 168:32]
  wire  _GEN_6889 = _T_1486 ? _GEN_6881 : _GEN_5833; // @[sequencer-master.scala 168:32]
  wire  _GEN_6890 = _T_1486 ? _GEN_6882 : _GEN_5834; // @[sequencer-master.scala 168:32]
  wire  _GEN_6891 = _T_1486 ? _GEN_6883 : _GEN_5835; // @[sequencer-master.scala 168:32]
  wire  _GEN_6892 = _T_1486 ? _GEN_6884 : _GEN_5836; // @[sequencer-master.scala 168:32]
  wire  _GEN_6893 = _T_1486 ? _GEN_6885 : _GEN_5837; // @[sequencer-master.scala 168:32]
  wire  _GEN_6894 = _GEN_32729 | _GEN_5854; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6895 = _GEN_32730 | _GEN_5855; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6896 = _GEN_32731 | _GEN_5856; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6897 = _GEN_32732 | _GEN_5857; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6898 = _GEN_32733 | _GEN_5858; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6899 = _GEN_32734 | _GEN_5859; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6900 = _GEN_32735 | _GEN_5860; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6901 = _GEN_32736 | _GEN_5861; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6902 = _T_1508 ? _GEN_6894 : _GEN_5854; // @[sequencer-master.scala 168:32]
  wire  _GEN_6903 = _T_1508 ? _GEN_6895 : _GEN_5855; // @[sequencer-master.scala 168:32]
  wire  _GEN_6904 = _T_1508 ? _GEN_6896 : _GEN_5856; // @[sequencer-master.scala 168:32]
  wire  _GEN_6905 = _T_1508 ? _GEN_6897 : _GEN_5857; // @[sequencer-master.scala 168:32]
  wire  _GEN_6906 = _T_1508 ? _GEN_6898 : _GEN_5858; // @[sequencer-master.scala 168:32]
  wire  _GEN_6907 = _T_1508 ? _GEN_6899 : _GEN_5859; // @[sequencer-master.scala 168:32]
  wire  _GEN_6908 = _T_1508 ? _GEN_6900 : _GEN_5860; // @[sequencer-master.scala 168:32]
  wire  _GEN_6909 = _T_1508 ? _GEN_6901 : _GEN_5861; // @[sequencer-master.scala 168:32]
  wire  _GEN_6910 = _GEN_32729 | _GEN_5878; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6911 = _GEN_32730 | _GEN_5879; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6912 = _GEN_32731 | _GEN_5880; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6913 = _GEN_32732 | _GEN_5881; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6914 = _GEN_32733 | _GEN_5882; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6915 = _GEN_32734 | _GEN_5883; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6916 = _GEN_32735 | _GEN_5884; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6917 = _GEN_32736 | _GEN_5885; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6918 = _T_1530 ? _GEN_6910 : _GEN_5878; // @[sequencer-master.scala 168:32]
  wire  _GEN_6919 = _T_1530 ? _GEN_6911 : _GEN_5879; // @[sequencer-master.scala 168:32]
  wire  _GEN_6920 = _T_1530 ? _GEN_6912 : _GEN_5880; // @[sequencer-master.scala 168:32]
  wire  _GEN_6921 = _T_1530 ? _GEN_6913 : _GEN_5881; // @[sequencer-master.scala 168:32]
  wire  _GEN_6922 = _T_1530 ? _GEN_6914 : _GEN_5882; // @[sequencer-master.scala 168:32]
  wire  _GEN_6923 = _T_1530 ? _GEN_6915 : _GEN_5883; // @[sequencer-master.scala 168:32]
  wire  _GEN_6924 = _T_1530 ? _GEN_6916 : _GEN_5884; // @[sequencer-master.scala 168:32]
  wire  _GEN_6925 = _T_1530 ? _GEN_6917 : _GEN_5885; // @[sequencer-master.scala 168:32]
  wire  _GEN_6926 = _GEN_32729 | _GEN_5902; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6927 = _GEN_32730 | _GEN_5903; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6928 = _GEN_32731 | _GEN_5904; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6929 = _GEN_32732 | _GEN_5905; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6930 = _GEN_32733 | _GEN_5906; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6931 = _GEN_32734 | _GEN_5907; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6932 = _GEN_32735 | _GEN_5908; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6933 = _GEN_32736 | _GEN_5909; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6934 = _T_1552 ? _GEN_6926 : _GEN_5902; // @[sequencer-master.scala 168:32]
  wire  _GEN_6935 = _T_1552 ? _GEN_6927 : _GEN_5903; // @[sequencer-master.scala 168:32]
  wire  _GEN_6936 = _T_1552 ? _GEN_6928 : _GEN_5904; // @[sequencer-master.scala 168:32]
  wire  _GEN_6937 = _T_1552 ? _GEN_6929 : _GEN_5905; // @[sequencer-master.scala 168:32]
  wire  _GEN_6938 = _T_1552 ? _GEN_6930 : _GEN_5906; // @[sequencer-master.scala 168:32]
  wire  _GEN_6939 = _T_1552 ? _GEN_6931 : _GEN_5907; // @[sequencer-master.scala 168:32]
  wire  _GEN_6940 = _T_1552 ? _GEN_6932 : _GEN_5908; // @[sequencer-master.scala 168:32]
  wire  _GEN_6941 = _T_1552 ? _GEN_6933 : _GEN_5909; // @[sequencer-master.scala 168:32]
  wire  _GEN_6942 = _GEN_32729 | _GEN_5926; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6943 = _GEN_32730 | _GEN_5927; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6944 = _GEN_32731 | _GEN_5928; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6945 = _GEN_32732 | _GEN_5929; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6946 = _GEN_32733 | _GEN_5930; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6947 = _GEN_32734 | _GEN_5931; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6948 = _GEN_32735 | _GEN_5932; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6949 = _GEN_32736 | _GEN_5933; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6950 = _T_1574 ? _GEN_6942 : _GEN_5926; // @[sequencer-master.scala 168:32]
  wire  _GEN_6951 = _T_1574 ? _GEN_6943 : _GEN_5927; // @[sequencer-master.scala 168:32]
  wire  _GEN_6952 = _T_1574 ? _GEN_6944 : _GEN_5928; // @[sequencer-master.scala 168:32]
  wire  _GEN_6953 = _T_1574 ? _GEN_6945 : _GEN_5929; // @[sequencer-master.scala 168:32]
  wire  _GEN_6954 = _T_1574 ? _GEN_6946 : _GEN_5930; // @[sequencer-master.scala 168:32]
  wire  _GEN_6955 = _T_1574 ? _GEN_6947 : _GEN_5931; // @[sequencer-master.scala 168:32]
  wire  _GEN_6956 = _T_1574 ? _GEN_6948 : _GEN_5932; // @[sequencer-master.scala 168:32]
  wire  _GEN_6957 = _T_1574 ? _GEN_6949 : _GEN_5933; // @[sequencer-master.scala 168:32]
  wire  _GEN_6958 = _GEN_32729 | _GEN_5950; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6959 = _GEN_32730 | _GEN_5951; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6960 = _GEN_32731 | _GEN_5952; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6961 = _GEN_32732 | _GEN_5953; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6962 = _GEN_32733 | _GEN_5954; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6963 = _GEN_32734 | _GEN_5955; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6964 = _GEN_32735 | _GEN_5956; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6965 = _GEN_32736 | _GEN_5957; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_6966 = _T_1596 ? _GEN_6958 : _GEN_5950; // @[sequencer-master.scala 168:32]
  wire  _GEN_6967 = _T_1596 ? _GEN_6959 : _GEN_5951; // @[sequencer-master.scala 168:32]
  wire  _GEN_6968 = _T_1596 ? _GEN_6960 : _GEN_5952; // @[sequencer-master.scala 168:32]
  wire  _GEN_6969 = _T_1596 ? _GEN_6961 : _GEN_5953; // @[sequencer-master.scala 168:32]
  wire  _GEN_6970 = _T_1596 ? _GEN_6962 : _GEN_5954; // @[sequencer-master.scala 168:32]
  wire  _GEN_6971 = _T_1596 ? _GEN_6963 : _GEN_5955; // @[sequencer-master.scala 168:32]
  wire  _GEN_6972 = _T_1596 ? _GEN_6964 : _GEN_5956; // @[sequencer-master.scala 168:32]
  wire  _GEN_6973 = _T_1596 ? _GEN_6965 : _GEN_5957; // @[sequencer-master.scala 168:32]
  wire  _GEN_34121 = 3'h0 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6974 = 3'h0 == _T_1645 | (_GEN_32729 | _GEN_5220); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34122 = 3'h1 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6975 = 3'h1 == _T_1645 | (_GEN_32730 | _GEN_5221); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34123 = 3'h2 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6976 = 3'h2 == _T_1645 | (_GEN_32731 | _GEN_5222); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34124 = 3'h3 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6977 = 3'h3 == _T_1645 | (_GEN_32732 | _GEN_5223); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34125 = 3'h4 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6978 = 3'h4 == _T_1645 | (_GEN_32733 | _GEN_5224); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34126 = 3'h5 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6979 = 3'h5 == _T_1645 | (_GEN_32734 | _GEN_5225); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34127 = 3'h6 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6980 = 3'h6 == _T_1645 | (_GEN_32735 | _GEN_5226); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_34128 = 3'h7 == _T_1645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6981 = 3'h7 == _T_1645 | (_GEN_32736 | _GEN_5227); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_6990 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6038; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6991 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6039; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6992 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6040; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6993 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6041; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6994 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6042; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6995 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6043; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6996 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6044; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6997 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6045; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_6998 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6270; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_6999 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6271; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7000 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6272; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7001 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6273; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7002 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6274; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7003 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6275; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7004 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6276; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7005 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6277; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_7006 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6518; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7007 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6519; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7008 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6520; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7009 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6521; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7010 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6522; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7011 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6523; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7012 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6524; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7013 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6525; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_7014 = 3'h0 == _T_1645 ? 1'h0 : _GEN_5742; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7015 = 3'h1 == _T_1645 ? 1'h0 : _GEN_5743; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7016 = 3'h2 == _T_1645 ? 1'h0 : _GEN_5744; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7017 = 3'h3 == _T_1645 ? 1'h0 : _GEN_5745; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7018 = 3'h4 == _T_1645 ? 1'h0 : _GEN_5746; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7019 = 3'h5 == _T_1645 ? 1'h0 : _GEN_5747; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7020 = 3'h6 == _T_1645 ? 1'h0 : _GEN_5748; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7021 = 3'h7 == _T_1645 ? 1'h0 : _GEN_5749; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_7022 = 3'h0 == _T_1645 ? 1'h0 : _GEN_5750; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7023 = 3'h1 == _T_1645 ? 1'h0 : _GEN_5751; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7024 = 3'h2 == _T_1645 ? 1'h0 : _GEN_5752; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7025 = 3'h3 == _T_1645 ? 1'h0 : _GEN_5753; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7026 = 3'h4 == _T_1645 ? 1'h0 : _GEN_5754; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7027 = 3'h5 == _T_1645 ? 1'h0 : _GEN_5755; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7028 = 3'h6 == _T_1645 ? 1'h0 : _GEN_5756; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7029 = 3'h7 == _T_1645 ? 1'h0 : _GEN_5757; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_7030 = _GEN_34121 | (_GEN_32729 | _GEN_5276); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7031 = _GEN_34122 | (_GEN_32730 | _GEN_5277); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7032 = _GEN_34123 | (_GEN_32731 | _GEN_5278); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7033 = _GEN_34124 | (_GEN_32732 | _GEN_5279); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7034 = _GEN_34125 | (_GEN_32733 | _GEN_5280); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7035 = _GEN_34126 | (_GEN_32734 | _GEN_5281); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7036 = _GEN_34127 | (_GEN_32735 | _GEN_5282); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7037 = _GEN_34128 | (_GEN_32736 | _GEN_5283); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_7038 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6574; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7039 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6575; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7040 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6576; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7041 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6577; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7042 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6578; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7043 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6579; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7044 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6580; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7045 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6581; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7046 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6726; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7047 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6727; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7048 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6728; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7049 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6729; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7050 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6730; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7051 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6731; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7052 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6732; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7053 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6733; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7054 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6854; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7055 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6855; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7056 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6856; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7057 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6857; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7058 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6858; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7059 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6859; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7060 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6860; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7061 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6861; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7062 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6590; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7063 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6591; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7064 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6592; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7065 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6593; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7066 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6594; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7067 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6595; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7068 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6596; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7069 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6597; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7070 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6742; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7071 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6743; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7072 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6744; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7073 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6745; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7074 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6746; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7075 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6747; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7076 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6748; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7077 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6749; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7078 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6870; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7079 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6871; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7080 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6872; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7081 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6873; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7082 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6874; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7083 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6875; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7084 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6876; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7085 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6877; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7086 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6606; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7087 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6607; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7088 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6608; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7089 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6609; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7090 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6610; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7091 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6611; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7092 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6612; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7093 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6613; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7094 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6758; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7095 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6759; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7096 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6760; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7097 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6761; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7098 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6762; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7099 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6763; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7100 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6764; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7101 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6765; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7102 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6886; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7103 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6887; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7104 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6888; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7105 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6889; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7106 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6890; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7107 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6891; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7108 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6892; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7109 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6893; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7110 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6622; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7111 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6623; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7112 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6624; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7113 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6625; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7114 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6626; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7115 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6627; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7116 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6628; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7117 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6629; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7118 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6774; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7119 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6775; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7120 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6776; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7121 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6777; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7122 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6778; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7123 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6779; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7124 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6780; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7125 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6781; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7126 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6902; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7127 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6903; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7128 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6904; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7129 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6905; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7130 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6906; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7131 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6907; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7132 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6908; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7133 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6909; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7134 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6638; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7135 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6639; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7136 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6640; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7137 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6641; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7138 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6642; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7139 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6643; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7140 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6644; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7141 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6645; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7142 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6790; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7143 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6791; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7144 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6792; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7145 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6793; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7146 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6794; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7147 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6795; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7148 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6796; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7149 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6797; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7150 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6918; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7151 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6919; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7152 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6920; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7153 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6921; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7154 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6922; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7155 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6923; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7156 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6924; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7157 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6925; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7158 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6654; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7159 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6655; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7160 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6656; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7161 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6657; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7162 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6658; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7163 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6659; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7164 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6660; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7165 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6661; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7166 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6806; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7167 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6807; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7168 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6808; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7169 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6809; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7170 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6810; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7171 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6811; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7172 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6812; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7173 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6813; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7174 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6934; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7175 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6935; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7176 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6936; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7177 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6937; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7178 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6938; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7179 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6939; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7180 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6940; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7181 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6941; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7182 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6670; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7183 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6671; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7184 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6672; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7185 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6673; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7186 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6674; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7187 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6675; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7188 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6676; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7189 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6677; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7190 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6822; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7191 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6823; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7192 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6824; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7193 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6825; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7194 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6826; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7195 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6827; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7196 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6828; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7197 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6829; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7198 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6950; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7199 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6951; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7200 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6952; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7201 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6953; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7202 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6954; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7203 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6955; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7204 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6956; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7205 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6957; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7206 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6686; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7207 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6687; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7208 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6688; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7209 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6689; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7210 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6690; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7211 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6691; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7212 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6692; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7213 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6693; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_7214 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6838; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7215 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6839; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7216 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6840; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7217 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6841; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7218 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6842; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7219 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6843; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7220 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6844; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7221 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6845; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_7222 = 3'h0 == _T_1645 ? 1'h0 : _GEN_6966; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7223 = 3'h1 == _T_1645 ? 1'h0 : _GEN_6967; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7224 = 3'h2 == _T_1645 ? 1'h0 : _GEN_6968; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7225 = 3'h3 == _T_1645 ? 1'h0 : _GEN_6969; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7226 = 3'h4 == _T_1645 ? 1'h0 : _GEN_6970; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7227 = 3'h5 == _T_1645 ? 1'h0 : _GEN_6971; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7228 = 3'h6 == _T_1645 ? 1'h0 : _GEN_6972; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7229 = 3'h7 == _T_1645 ? 1'h0 : _GEN_6973; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_7230 = 3'h0 == _T_1645 ? 1'h0 : _GEN_5958; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7231 = 3'h1 == _T_1645 ? 1'h0 : _GEN_5959; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7232 = 3'h2 == _T_1645 ? 1'h0 : _GEN_5960; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7233 = 3'h3 == _T_1645 ? 1'h0 : _GEN_5961; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7234 = 3'h4 == _T_1645 ? 1'h0 : _GEN_5962; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7235 = 3'h5 == _T_1645 ? 1'h0 : _GEN_5963; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7236 = 3'h6 == _T_1645 ? 1'h0 : _GEN_5964; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7237 = 3'h7 == _T_1645 ? 1'h0 : _GEN_5965; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_7246 = _GEN_34121 | e_0_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7247 = _GEN_34122 | e_1_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7248 = _GEN_34123 | e_2_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7249 = _GEN_34124 | e_3_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7250 = _GEN_34125 | e_4_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7251 = _GEN_34126 | e_5_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7252 = _GEN_34127 | e_6_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_7253 = _GEN_34128 | e_7_active_vidu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_7254 = 3'h0 == _T_1645 ? io_op_bits_fn_union : _GEN_5982; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7255 = 3'h1 == _T_1645 ? io_op_bits_fn_union : _GEN_5983; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7256 = 3'h2 == _T_1645 ? io_op_bits_fn_union : _GEN_5984; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7257 = 3'h3 == _T_1645 ? io_op_bits_fn_union : _GEN_5985; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7258 = 3'h4 == _T_1645 ? io_op_bits_fn_union : _GEN_5986; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7259 = 3'h5 == _T_1645 ? io_op_bits_fn_union : _GEN_5987; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7260 = 3'h6 == _T_1645 ? io_op_bits_fn_union : _GEN_5988; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_7261 = 3'h7 == _T_1645 ? io_op_bits_fn_union : _GEN_5989; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [7:0] _GEN_7262 = 3'h0 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5636; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7263 = 3'h1 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5637; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7264 = 3'h2 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5638; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7265 = 3'h3 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5639; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7266 = 3'h4 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5640; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7267 = 3'h5 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5641; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7268 = 3'h6 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5642; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7269 = 3'h7 == _T_1645 ? io_op_bits_base_vd_id : _GEN_5643; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7270 = 3'h0 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7022; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7271 = 3'h1 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7023; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7272 = 3'h2 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7024; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7273 = 3'h3 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7025; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7274 = 3'h4 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7026; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7275 = 3'h5 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7027; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7276 = 3'h6 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7028; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7277 = 3'h7 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_7029; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7278 = 3'h0 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5644; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7279 = 3'h1 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5645; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7280 = 3'h2 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5646; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7281 = 3'h3 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5647; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7282 = 3'h4 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5648; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7283 = 3'h5 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5649; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7284 = 3'h6 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5650; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7285 = 3'h7 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_5651; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7286 = 3'h0 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5652; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7287 = 3'h1 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5653; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7288 = 3'h2 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5654; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7289 = 3'h3 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5655; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7290 = 3'h4 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5656; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7291 = 3'h5 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5657; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7292 = 3'h6 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5658; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_7293 = 3'h7 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_5659; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7294 = 3'h0 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5660; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7295 = 3'h1 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5661; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7296 = 3'h2 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5662; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7297 = 3'h3 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5663; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7298 = 3'h4 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5664; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7299 = 3'h5 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5665; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7300 = 3'h6 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5666; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_7301 = 3'h7 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_5667; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_7302 = 3'h0 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5668; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7303 = 3'h1 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5669; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7304 = 3'h2 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5670; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7305 = 3'h3 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5671; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7306 = 3'h4 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5672; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7307 = 3'h5 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5673; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7308 = 3'h6 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5674; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7309 = 3'h7 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_5675; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_7310 = io_op_bits_base_vd_valid ? _GEN_7262 : _GEN_5636; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7311 = io_op_bits_base_vd_valid ? _GEN_7263 : _GEN_5637; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7312 = io_op_bits_base_vd_valid ? _GEN_7264 : _GEN_5638; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7313 = io_op_bits_base_vd_valid ? _GEN_7265 : _GEN_5639; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7314 = io_op_bits_base_vd_valid ? _GEN_7266 : _GEN_5640; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7315 = io_op_bits_base_vd_valid ? _GEN_7267 : _GEN_5641; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7316 = io_op_bits_base_vd_valid ? _GEN_7268 : _GEN_5642; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7317 = io_op_bits_base_vd_valid ? _GEN_7269 : _GEN_5643; // @[sequencer-master.scala 362:41]
  wire  _GEN_7318 = io_op_bits_base_vd_valid ? _GEN_7270 : _GEN_7022; // @[sequencer-master.scala 362:41]
  wire  _GEN_7319 = io_op_bits_base_vd_valid ? _GEN_7271 : _GEN_7023; // @[sequencer-master.scala 362:41]
  wire  _GEN_7320 = io_op_bits_base_vd_valid ? _GEN_7272 : _GEN_7024; // @[sequencer-master.scala 362:41]
  wire  _GEN_7321 = io_op_bits_base_vd_valid ? _GEN_7273 : _GEN_7025; // @[sequencer-master.scala 362:41]
  wire  _GEN_7322 = io_op_bits_base_vd_valid ? _GEN_7274 : _GEN_7026; // @[sequencer-master.scala 362:41]
  wire  _GEN_7323 = io_op_bits_base_vd_valid ? _GEN_7275 : _GEN_7027; // @[sequencer-master.scala 362:41]
  wire  _GEN_7324 = io_op_bits_base_vd_valid ? _GEN_7276 : _GEN_7028; // @[sequencer-master.scala 362:41]
  wire  _GEN_7325 = io_op_bits_base_vd_valid ? _GEN_7277 : _GEN_7029; // @[sequencer-master.scala 362:41]
  wire  _GEN_7326 = io_op_bits_base_vd_valid ? _GEN_7278 : _GEN_5644; // @[sequencer-master.scala 362:41]
  wire  _GEN_7327 = io_op_bits_base_vd_valid ? _GEN_7279 : _GEN_5645; // @[sequencer-master.scala 362:41]
  wire  _GEN_7328 = io_op_bits_base_vd_valid ? _GEN_7280 : _GEN_5646; // @[sequencer-master.scala 362:41]
  wire  _GEN_7329 = io_op_bits_base_vd_valid ? _GEN_7281 : _GEN_5647; // @[sequencer-master.scala 362:41]
  wire  _GEN_7330 = io_op_bits_base_vd_valid ? _GEN_7282 : _GEN_5648; // @[sequencer-master.scala 362:41]
  wire  _GEN_7331 = io_op_bits_base_vd_valid ? _GEN_7283 : _GEN_5649; // @[sequencer-master.scala 362:41]
  wire  _GEN_7332 = io_op_bits_base_vd_valid ? _GEN_7284 : _GEN_5650; // @[sequencer-master.scala 362:41]
  wire  _GEN_7333 = io_op_bits_base_vd_valid ? _GEN_7285 : _GEN_5651; // @[sequencer-master.scala 362:41]
  wire  _GEN_7334 = io_op_bits_base_vd_valid ? _GEN_7286 : _GEN_5652; // @[sequencer-master.scala 362:41]
  wire  _GEN_7335 = io_op_bits_base_vd_valid ? _GEN_7287 : _GEN_5653; // @[sequencer-master.scala 362:41]
  wire  _GEN_7336 = io_op_bits_base_vd_valid ? _GEN_7288 : _GEN_5654; // @[sequencer-master.scala 362:41]
  wire  _GEN_7337 = io_op_bits_base_vd_valid ? _GEN_7289 : _GEN_5655; // @[sequencer-master.scala 362:41]
  wire  _GEN_7338 = io_op_bits_base_vd_valid ? _GEN_7290 : _GEN_5656; // @[sequencer-master.scala 362:41]
  wire  _GEN_7339 = io_op_bits_base_vd_valid ? _GEN_7291 : _GEN_5657; // @[sequencer-master.scala 362:41]
  wire  _GEN_7340 = io_op_bits_base_vd_valid ? _GEN_7292 : _GEN_5658; // @[sequencer-master.scala 362:41]
  wire  _GEN_7341 = io_op_bits_base_vd_valid ? _GEN_7293 : _GEN_5659; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7342 = io_op_bits_base_vd_valid ? _GEN_7294 : _GEN_5660; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7343 = io_op_bits_base_vd_valid ? _GEN_7295 : _GEN_5661; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7344 = io_op_bits_base_vd_valid ? _GEN_7296 : _GEN_5662; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7345 = io_op_bits_base_vd_valid ? _GEN_7297 : _GEN_5663; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7346 = io_op_bits_base_vd_valid ? _GEN_7298 : _GEN_5664; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7347 = io_op_bits_base_vd_valid ? _GEN_7299 : _GEN_5665; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7348 = io_op_bits_base_vd_valid ? _GEN_7300 : _GEN_5666; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_7349 = io_op_bits_base_vd_valid ? _GEN_7301 : _GEN_5667; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7350 = io_op_bits_base_vd_valid ? _GEN_7302 : _GEN_5668; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7351 = io_op_bits_base_vd_valid ? _GEN_7303 : _GEN_5669; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7352 = io_op_bits_base_vd_valid ? _GEN_7304 : _GEN_5670; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7353 = io_op_bits_base_vd_valid ? _GEN_7305 : _GEN_5671; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7354 = io_op_bits_base_vd_valid ? _GEN_7306 : _GEN_5672; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7355 = io_op_bits_base_vd_valid ? _GEN_7307 : _GEN_5673; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7356 = io_op_bits_base_vd_valid ? _GEN_7308 : _GEN_5674; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_7357 = io_op_bits_base_vd_valid ? _GEN_7309 : _GEN_5675; // @[sequencer-master.scala 362:41]
  wire  _GEN_7358 = _GEN_34121 | _GEN_7046; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7359 = _GEN_34122 | _GEN_7047; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7360 = _GEN_34123 | _GEN_7048; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7361 = _GEN_34124 | _GEN_7049; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7362 = _GEN_34125 | _GEN_7050; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7363 = _GEN_34126 | _GEN_7051; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7364 = _GEN_34127 | _GEN_7052; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7365 = _GEN_34128 | _GEN_7053; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7366 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7358 : _GEN_7046; // @[sequencer-master.scala 161:86]
  wire  _GEN_7367 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7359 : _GEN_7047; // @[sequencer-master.scala 161:86]
  wire  _GEN_7368 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7360 : _GEN_7048; // @[sequencer-master.scala 161:86]
  wire  _GEN_7369 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7361 : _GEN_7049; // @[sequencer-master.scala 161:86]
  wire  _GEN_7370 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7362 : _GEN_7050; // @[sequencer-master.scala 161:86]
  wire  _GEN_7371 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7363 : _GEN_7051; // @[sequencer-master.scala 161:86]
  wire  _GEN_7372 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7364 : _GEN_7052; // @[sequencer-master.scala 161:86]
  wire  _GEN_7373 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_7365 : _GEN_7053; // @[sequencer-master.scala 161:86]
  wire  _GEN_7374 = _GEN_34121 | _GEN_7070; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7375 = _GEN_34122 | _GEN_7071; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7376 = _GEN_34123 | _GEN_7072; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7377 = _GEN_34124 | _GEN_7073; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7378 = _GEN_34125 | _GEN_7074; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7379 = _GEN_34126 | _GEN_7075; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7380 = _GEN_34127 | _GEN_7076; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7381 = _GEN_34128 | _GEN_7077; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7382 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7374 : _GEN_7070; // @[sequencer-master.scala 161:86]
  wire  _GEN_7383 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7375 : _GEN_7071; // @[sequencer-master.scala 161:86]
  wire  _GEN_7384 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7376 : _GEN_7072; // @[sequencer-master.scala 161:86]
  wire  _GEN_7385 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7377 : _GEN_7073; // @[sequencer-master.scala 161:86]
  wire  _GEN_7386 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7378 : _GEN_7074; // @[sequencer-master.scala 161:86]
  wire  _GEN_7387 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7379 : _GEN_7075; // @[sequencer-master.scala 161:86]
  wire  _GEN_7388 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7380 : _GEN_7076; // @[sequencer-master.scala 161:86]
  wire  _GEN_7389 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_7381 : _GEN_7077; // @[sequencer-master.scala 161:86]
  wire  _GEN_7390 = _GEN_34121 | _GEN_7094; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7391 = _GEN_34122 | _GEN_7095; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7392 = _GEN_34123 | _GEN_7096; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7393 = _GEN_34124 | _GEN_7097; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7394 = _GEN_34125 | _GEN_7098; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7395 = _GEN_34126 | _GEN_7099; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7396 = _GEN_34127 | _GEN_7100; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7397 = _GEN_34128 | _GEN_7101; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7398 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7390 : _GEN_7094; // @[sequencer-master.scala 161:86]
  wire  _GEN_7399 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7391 : _GEN_7095; // @[sequencer-master.scala 161:86]
  wire  _GEN_7400 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7392 : _GEN_7096; // @[sequencer-master.scala 161:86]
  wire  _GEN_7401 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7393 : _GEN_7097; // @[sequencer-master.scala 161:86]
  wire  _GEN_7402 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7394 : _GEN_7098; // @[sequencer-master.scala 161:86]
  wire  _GEN_7403 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7395 : _GEN_7099; // @[sequencer-master.scala 161:86]
  wire  _GEN_7404 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7396 : _GEN_7100; // @[sequencer-master.scala 161:86]
  wire  _GEN_7405 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_7397 : _GEN_7101; // @[sequencer-master.scala 161:86]
  wire  _GEN_7406 = _GEN_34121 | _GEN_7118; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7407 = _GEN_34122 | _GEN_7119; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7408 = _GEN_34123 | _GEN_7120; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7409 = _GEN_34124 | _GEN_7121; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7410 = _GEN_34125 | _GEN_7122; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7411 = _GEN_34126 | _GEN_7123; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7412 = _GEN_34127 | _GEN_7124; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7413 = _GEN_34128 | _GEN_7125; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7414 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7406 : _GEN_7118; // @[sequencer-master.scala 161:86]
  wire  _GEN_7415 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7407 : _GEN_7119; // @[sequencer-master.scala 161:86]
  wire  _GEN_7416 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7408 : _GEN_7120; // @[sequencer-master.scala 161:86]
  wire  _GEN_7417 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7409 : _GEN_7121; // @[sequencer-master.scala 161:86]
  wire  _GEN_7418 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7410 : _GEN_7122; // @[sequencer-master.scala 161:86]
  wire  _GEN_7419 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7411 : _GEN_7123; // @[sequencer-master.scala 161:86]
  wire  _GEN_7420 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7412 : _GEN_7124; // @[sequencer-master.scala 161:86]
  wire  _GEN_7421 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_7413 : _GEN_7125; // @[sequencer-master.scala 161:86]
  wire  _GEN_7422 = _GEN_34121 | _GEN_7142; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7423 = _GEN_34122 | _GEN_7143; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7424 = _GEN_34123 | _GEN_7144; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7425 = _GEN_34124 | _GEN_7145; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7426 = _GEN_34125 | _GEN_7146; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7427 = _GEN_34126 | _GEN_7147; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7428 = _GEN_34127 | _GEN_7148; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7429 = _GEN_34128 | _GEN_7149; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7430 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7422 : _GEN_7142; // @[sequencer-master.scala 161:86]
  wire  _GEN_7431 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7423 : _GEN_7143; // @[sequencer-master.scala 161:86]
  wire  _GEN_7432 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7424 : _GEN_7144; // @[sequencer-master.scala 161:86]
  wire  _GEN_7433 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7425 : _GEN_7145; // @[sequencer-master.scala 161:86]
  wire  _GEN_7434 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7426 : _GEN_7146; // @[sequencer-master.scala 161:86]
  wire  _GEN_7435 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7427 : _GEN_7147; // @[sequencer-master.scala 161:86]
  wire  _GEN_7436 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7428 : _GEN_7148; // @[sequencer-master.scala 161:86]
  wire  _GEN_7437 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_7429 : _GEN_7149; // @[sequencer-master.scala 161:86]
  wire  _GEN_7438 = _GEN_34121 | _GEN_7166; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7439 = _GEN_34122 | _GEN_7167; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7440 = _GEN_34123 | _GEN_7168; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7441 = _GEN_34124 | _GEN_7169; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7442 = _GEN_34125 | _GEN_7170; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7443 = _GEN_34126 | _GEN_7171; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7444 = _GEN_34127 | _GEN_7172; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7445 = _GEN_34128 | _GEN_7173; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7446 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7438 : _GEN_7166; // @[sequencer-master.scala 161:86]
  wire  _GEN_7447 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7439 : _GEN_7167; // @[sequencer-master.scala 161:86]
  wire  _GEN_7448 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7440 : _GEN_7168; // @[sequencer-master.scala 161:86]
  wire  _GEN_7449 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7441 : _GEN_7169; // @[sequencer-master.scala 161:86]
  wire  _GEN_7450 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7442 : _GEN_7170; // @[sequencer-master.scala 161:86]
  wire  _GEN_7451 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7443 : _GEN_7171; // @[sequencer-master.scala 161:86]
  wire  _GEN_7452 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7444 : _GEN_7172; // @[sequencer-master.scala 161:86]
  wire  _GEN_7453 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_7445 : _GEN_7173; // @[sequencer-master.scala 161:86]
  wire  _GEN_7454 = _GEN_34121 | _GEN_7190; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7455 = _GEN_34122 | _GEN_7191; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7456 = _GEN_34123 | _GEN_7192; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7457 = _GEN_34124 | _GEN_7193; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7458 = _GEN_34125 | _GEN_7194; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7459 = _GEN_34126 | _GEN_7195; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7460 = _GEN_34127 | _GEN_7196; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7461 = _GEN_34128 | _GEN_7197; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7462 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7454 : _GEN_7190; // @[sequencer-master.scala 161:86]
  wire  _GEN_7463 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7455 : _GEN_7191; // @[sequencer-master.scala 161:86]
  wire  _GEN_7464 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7456 : _GEN_7192; // @[sequencer-master.scala 161:86]
  wire  _GEN_7465 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7457 : _GEN_7193; // @[sequencer-master.scala 161:86]
  wire  _GEN_7466 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7458 : _GEN_7194; // @[sequencer-master.scala 161:86]
  wire  _GEN_7467 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7459 : _GEN_7195; // @[sequencer-master.scala 161:86]
  wire  _GEN_7468 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7460 : _GEN_7196; // @[sequencer-master.scala 161:86]
  wire  _GEN_7469 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_7461 : _GEN_7197; // @[sequencer-master.scala 161:86]
  wire  _GEN_7470 = _GEN_34121 | _GEN_7214; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7471 = _GEN_34122 | _GEN_7215; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7472 = _GEN_34123 | _GEN_7216; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7473 = _GEN_34124 | _GEN_7217; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7474 = _GEN_34125 | _GEN_7218; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7475 = _GEN_34126 | _GEN_7219; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7476 = _GEN_34127 | _GEN_7220; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7477 = _GEN_34128 | _GEN_7221; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_7478 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7470 : _GEN_7214; // @[sequencer-master.scala 161:86]
  wire  _GEN_7479 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7471 : _GEN_7215; // @[sequencer-master.scala 161:86]
  wire  _GEN_7480 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7472 : _GEN_7216; // @[sequencer-master.scala 161:86]
  wire  _GEN_7481 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7473 : _GEN_7217; // @[sequencer-master.scala 161:86]
  wire  _GEN_7482 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7474 : _GEN_7218; // @[sequencer-master.scala 161:86]
  wire  _GEN_7483 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7475 : _GEN_7219; // @[sequencer-master.scala 161:86]
  wire  _GEN_7484 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7476 : _GEN_7220; // @[sequencer-master.scala 161:86]
  wire  _GEN_7485 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_7477 : _GEN_7221; // @[sequencer-master.scala 161:86]
  wire  _GEN_7486 = _GEN_34121 | _GEN_7054; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7487 = _GEN_34122 | _GEN_7055; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7488 = _GEN_34123 | _GEN_7056; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7489 = _GEN_34124 | _GEN_7057; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7490 = _GEN_34125 | _GEN_7058; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7491 = _GEN_34126 | _GEN_7059; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7492 = _GEN_34127 | _GEN_7060; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7493 = _GEN_34128 | _GEN_7061; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7494 = _T_1442 ? _GEN_7486 : _GEN_7054; // @[sequencer-master.scala 168:32]
  wire  _GEN_7495 = _T_1442 ? _GEN_7487 : _GEN_7055; // @[sequencer-master.scala 168:32]
  wire  _GEN_7496 = _T_1442 ? _GEN_7488 : _GEN_7056; // @[sequencer-master.scala 168:32]
  wire  _GEN_7497 = _T_1442 ? _GEN_7489 : _GEN_7057; // @[sequencer-master.scala 168:32]
  wire  _GEN_7498 = _T_1442 ? _GEN_7490 : _GEN_7058; // @[sequencer-master.scala 168:32]
  wire  _GEN_7499 = _T_1442 ? _GEN_7491 : _GEN_7059; // @[sequencer-master.scala 168:32]
  wire  _GEN_7500 = _T_1442 ? _GEN_7492 : _GEN_7060; // @[sequencer-master.scala 168:32]
  wire  _GEN_7501 = _T_1442 ? _GEN_7493 : _GEN_7061; // @[sequencer-master.scala 168:32]
  wire  _GEN_7502 = _GEN_34121 | _GEN_7078; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7503 = _GEN_34122 | _GEN_7079; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7504 = _GEN_34123 | _GEN_7080; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7505 = _GEN_34124 | _GEN_7081; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7506 = _GEN_34125 | _GEN_7082; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7507 = _GEN_34126 | _GEN_7083; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7508 = _GEN_34127 | _GEN_7084; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7509 = _GEN_34128 | _GEN_7085; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7510 = _T_1464 ? _GEN_7502 : _GEN_7078; // @[sequencer-master.scala 168:32]
  wire  _GEN_7511 = _T_1464 ? _GEN_7503 : _GEN_7079; // @[sequencer-master.scala 168:32]
  wire  _GEN_7512 = _T_1464 ? _GEN_7504 : _GEN_7080; // @[sequencer-master.scala 168:32]
  wire  _GEN_7513 = _T_1464 ? _GEN_7505 : _GEN_7081; // @[sequencer-master.scala 168:32]
  wire  _GEN_7514 = _T_1464 ? _GEN_7506 : _GEN_7082; // @[sequencer-master.scala 168:32]
  wire  _GEN_7515 = _T_1464 ? _GEN_7507 : _GEN_7083; // @[sequencer-master.scala 168:32]
  wire  _GEN_7516 = _T_1464 ? _GEN_7508 : _GEN_7084; // @[sequencer-master.scala 168:32]
  wire  _GEN_7517 = _T_1464 ? _GEN_7509 : _GEN_7085; // @[sequencer-master.scala 168:32]
  wire  _GEN_7518 = _GEN_34121 | _GEN_7102; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7519 = _GEN_34122 | _GEN_7103; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7520 = _GEN_34123 | _GEN_7104; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7521 = _GEN_34124 | _GEN_7105; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7522 = _GEN_34125 | _GEN_7106; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7523 = _GEN_34126 | _GEN_7107; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7524 = _GEN_34127 | _GEN_7108; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7525 = _GEN_34128 | _GEN_7109; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7526 = _T_1486 ? _GEN_7518 : _GEN_7102; // @[sequencer-master.scala 168:32]
  wire  _GEN_7527 = _T_1486 ? _GEN_7519 : _GEN_7103; // @[sequencer-master.scala 168:32]
  wire  _GEN_7528 = _T_1486 ? _GEN_7520 : _GEN_7104; // @[sequencer-master.scala 168:32]
  wire  _GEN_7529 = _T_1486 ? _GEN_7521 : _GEN_7105; // @[sequencer-master.scala 168:32]
  wire  _GEN_7530 = _T_1486 ? _GEN_7522 : _GEN_7106; // @[sequencer-master.scala 168:32]
  wire  _GEN_7531 = _T_1486 ? _GEN_7523 : _GEN_7107; // @[sequencer-master.scala 168:32]
  wire  _GEN_7532 = _T_1486 ? _GEN_7524 : _GEN_7108; // @[sequencer-master.scala 168:32]
  wire  _GEN_7533 = _T_1486 ? _GEN_7525 : _GEN_7109; // @[sequencer-master.scala 168:32]
  wire  _GEN_7534 = _GEN_34121 | _GEN_7126; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7535 = _GEN_34122 | _GEN_7127; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7536 = _GEN_34123 | _GEN_7128; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7537 = _GEN_34124 | _GEN_7129; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7538 = _GEN_34125 | _GEN_7130; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7539 = _GEN_34126 | _GEN_7131; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7540 = _GEN_34127 | _GEN_7132; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7541 = _GEN_34128 | _GEN_7133; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7542 = _T_1508 ? _GEN_7534 : _GEN_7126; // @[sequencer-master.scala 168:32]
  wire  _GEN_7543 = _T_1508 ? _GEN_7535 : _GEN_7127; // @[sequencer-master.scala 168:32]
  wire  _GEN_7544 = _T_1508 ? _GEN_7536 : _GEN_7128; // @[sequencer-master.scala 168:32]
  wire  _GEN_7545 = _T_1508 ? _GEN_7537 : _GEN_7129; // @[sequencer-master.scala 168:32]
  wire  _GEN_7546 = _T_1508 ? _GEN_7538 : _GEN_7130; // @[sequencer-master.scala 168:32]
  wire  _GEN_7547 = _T_1508 ? _GEN_7539 : _GEN_7131; // @[sequencer-master.scala 168:32]
  wire  _GEN_7548 = _T_1508 ? _GEN_7540 : _GEN_7132; // @[sequencer-master.scala 168:32]
  wire  _GEN_7549 = _T_1508 ? _GEN_7541 : _GEN_7133; // @[sequencer-master.scala 168:32]
  wire  _GEN_7550 = _GEN_34121 | _GEN_7150; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7551 = _GEN_34122 | _GEN_7151; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7552 = _GEN_34123 | _GEN_7152; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7553 = _GEN_34124 | _GEN_7153; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7554 = _GEN_34125 | _GEN_7154; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7555 = _GEN_34126 | _GEN_7155; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7556 = _GEN_34127 | _GEN_7156; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7557 = _GEN_34128 | _GEN_7157; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7558 = _T_1530 ? _GEN_7550 : _GEN_7150; // @[sequencer-master.scala 168:32]
  wire  _GEN_7559 = _T_1530 ? _GEN_7551 : _GEN_7151; // @[sequencer-master.scala 168:32]
  wire  _GEN_7560 = _T_1530 ? _GEN_7552 : _GEN_7152; // @[sequencer-master.scala 168:32]
  wire  _GEN_7561 = _T_1530 ? _GEN_7553 : _GEN_7153; // @[sequencer-master.scala 168:32]
  wire  _GEN_7562 = _T_1530 ? _GEN_7554 : _GEN_7154; // @[sequencer-master.scala 168:32]
  wire  _GEN_7563 = _T_1530 ? _GEN_7555 : _GEN_7155; // @[sequencer-master.scala 168:32]
  wire  _GEN_7564 = _T_1530 ? _GEN_7556 : _GEN_7156; // @[sequencer-master.scala 168:32]
  wire  _GEN_7565 = _T_1530 ? _GEN_7557 : _GEN_7157; // @[sequencer-master.scala 168:32]
  wire  _GEN_7566 = _GEN_34121 | _GEN_7174; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7567 = _GEN_34122 | _GEN_7175; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7568 = _GEN_34123 | _GEN_7176; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7569 = _GEN_34124 | _GEN_7177; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7570 = _GEN_34125 | _GEN_7178; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7571 = _GEN_34126 | _GEN_7179; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7572 = _GEN_34127 | _GEN_7180; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7573 = _GEN_34128 | _GEN_7181; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7574 = _T_1552 ? _GEN_7566 : _GEN_7174; // @[sequencer-master.scala 168:32]
  wire  _GEN_7575 = _T_1552 ? _GEN_7567 : _GEN_7175; // @[sequencer-master.scala 168:32]
  wire  _GEN_7576 = _T_1552 ? _GEN_7568 : _GEN_7176; // @[sequencer-master.scala 168:32]
  wire  _GEN_7577 = _T_1552 ? _GEN_7569 : _GEN_7177; // @[sequencer-master.scala 168:32]
  wire  _GEN_7578 = _T_1552 ? _GEN_7570 : _GEN_7178; // @[sequencer-master.scala 168:32]
  wire  _GEN_7579 = _T_1552 ? _GEN_7571 : _GEN_7179; // @[sequencer-master.scala 168:32]
  wire  _GEN_7580 = _T_1552 ? _GEN_7572 : _GEN_7180; // @[sequencer-master.scala 168:32]
  wire  _GEN_7581 = _T_1552 ? _GEN_7573 : _GEN_7181; // @[sequencer-master.scala 168:32]
  wire  _GEN_7582 = _GEN_34121 | _GEN_7198; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7583 = _GEN_34122 | _GEN_7199; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7584 = _GEN_34123 | _GEN_7200; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7585 = _GEN_34124 | _GEN_7201; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7586 = _GEN_34125 | _GEN_7202; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7587 = _GEN_34126 | _GEN_7203; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7588 = _GEN_34127 | _GEN_7204; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7589 = _GEN_34128 | _GEN_7205; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7590 = _T_1574 ? _GEN_7582 : _GEN_7198; // @[sequencer-master.scala 168:32]
  wire  _GEN_7591 = _T_1574 ? _GEN_7583 : _GEN_7199; // @[sequencer-master.scala 168:32]
  wire  _GEN_7592 = _T_1574 ? _GEN_7584 : _GEN_7200; // @[sequencer-master.scala 168:32]
  wire  _GEN_7593 = _T_1574 ? _GEN_7585 : _GEN_7201; // @[sequencer-master.scala 168:32]
  wire  _GEN_7594 = _T_1574 ? _GEN_7586 : _GEN_7202; // @[sequencer-master.scala 168:32]
  wire  _GEN_7595 = _T_1574 ? _GEN_7587 : _GEN_7203; // @[sequencer-master.scala 168:32]
  wire  _GEN_7596 = _T_1574 ? _GEN_7588 : _GEN_7204; // @[sequencer-master.scala 168:32]
  wire  _GEN_7597 = _T_1574 ? _GEN_7589 : _GEN_7205; // @[sequencer-master.scala 168:32]
  wire  _GEN_7598 = _GEN_34121 | _GEN_7222; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7599 = _GEN_34122 | _GEN_7223; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7600 = _GEN_34123 | _GEN_7224; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7601 = _GEN_34124 | _GEN_7225; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7602 = _GEN_34125 | _GEN_7226; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7603 = _GEN_34126 | _GEN_7227; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7604 = _GEN_34127 | _GEN_7228; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7605 = _GEN_34128 | _GEN_7229; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_7606 = _T_1596 ? _GEN_7598 : _GEN_7222; // @[sequencer-master.scala 168:32]
  wire  _GEN_7607 = _T_1596 ? _GEN_7599 : _GEN_7223; // @[sequencer-master.scala 168:32]
  wire  _GEN_7608 = _T_1596 ? _GEN_7600 : _GEN_7224; // @[sequencer-master.scala 168:32]
  wire  _GEN_7609 = _T_1596 ? _GEN_7601 : _GEN_7225; // @[sequencer-master.scala 168:32]
  wire  _GEN_7610 = _T_1596 ? _GEN_7602 : _GEN_7226; // @[sequencer-master.scala 168:32]
  wire  _GEN_7611 = _T_1596 ? _GEN_7603 : _GEN_7227; // @[sequencer-master.scala 168:32]
  wire  _GEN_7612 = _T_1596 ? _GEN_7604 : _GEN_7228; // @[sequencer-master.scala 168:32]
  wire  _GEN_7613 = _T_1596 ? _GEN_7605 : _GEN_7229; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_7614 = 3'h0 == _T_1645 ? 2'h0 : _GEN_6694; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7615 = 3'h1 == _T_1645 ? 2'h0 : _GEN_6695; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7616 = 3'h2 == _T_1645 ? 2'h0 : _GEN_6696; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7617 = 3'h3 == _T_1645 ? 2'h0 : _GEN_6697; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7618 = 3'h4 == _T_1645 ? 2'h0 : _GEN_6698; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7619 = 3'h5 == _T_1645 ? 2'h0 : _GEN_6699; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7620 = 3'h6 == _T_1645 ? 2'h0 : _GEN_6700; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_7621 = 3'h7 == _T_1645 ? 2'h0 : _GEN_6701; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_7622 = 3'h0 == _T_1645 ? 4'h0 : _GEN_6702; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7623 = 3'h1 == _T_1645 ? 4'h0 : _GEN_6703; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7624 = 3'h2 == _T_1645 ? 4'h0 : _GEN_6704; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7625 = 3'h3 == _T_1645 ? 4'h0 : _GEN_6705; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7626 = 3'h4 == _T_1645 ? 4'h0 : _GEN_6706; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7627 = 3'h5 == _T_1645 ? 4'h0 : _GEN_6707; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7628 = 3'h6 == _T_1645 ? 4'h0 : _GEN_6708; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_7629 = 3'h7 == _T_1645 ? 4'h0 : _GEN_6709; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_7630 = 3'h0 == _T_1645 ? 3'h0 : _GEN_6710; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7631 = 3'h1 == _T_1645 ? 3'h0 : _GEN_6711; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7632 = 3'h2 == _T_1645 ? 3'h0 : _GEN_6712; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7633 = 3'h3 == _T_1645 ? 3'h0 : _GEN_6713; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7634 = 3'h4 == _T_1645 ? 3'h0 : _GEN_6714; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7635 = 3'h5 == _T_1645 ? 3'h0 : _GEN_6715; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7636 = 3'h6 == _T_1645 ? 3'h0 : _GEN_6716; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_7637 = 3'h7 == _T_1645 ? 3'h0 : _GEN_6717; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_7638 = io_op_bits_active_vidiv ? _GEN_6974 : _GEN_5220; // @[sequencer-master.scala 643:40]
  wire  _GEN_7639 = io_op_bits_active_vidiv ? _GEN_6975 : _GEN_5221; // @[sequencer-master.scala 643:40]
  wire  _GEN_7640 = io_op_bits_active_vidiv ? _GEN_6976 : _GEN_5222; // @[sequencer-master.scala 643:40]
  wire  _GEN_7641 = io_op_bits_active_vidiv ? _GEN_6977 : _GEN_5223; // @[sequencer-master.scala 643:40]
  wire  _GEN_7642 = io_op_bits_active_vidiv ? _GEN_6978 : _GEN_5224; // @[sequencer-master.scala 643:40]
  wire  _GEN_7643 = io_op_bits_active_vidiv ? _GEN_6979 : _GEN_5225; // @[sequencer-master.scala 643:40]
  wire  _GEN_7644 = io_op_bits_active_vidiv ? _GEN_6980 : _GEN_5226; // @[sequencer-master.scala 643:40]
  wire  _GEN_7645 = io_op_bits_active_vidiv ? _GEN_6981 : _GEN_5227; // @[sequencer-master.scala 643:40]
  wire  _GEN_7654 = io_op_bits_active_vidiv ? _GEN_6990 : _GEN_5236; // @[sequencer-master.scala 643:40]
  wire  _GEN_7655 = io_op_bits_active_vidiv ? _GEN_6991 : _GEN_5237; // @[sequencer-master.scala 643:40]
  wire  _GEN_7656 = io_op_bits_active_vidiv ? _GEN_6992 : _GEN_5238; // @[sequencer-master.scala 643:40]
  wire  _GEN_7657 = io_op_bits_active_vidiv ? _GEN_6993 : _GEN_5239; // @[sequencer-master.scala 643:40]
  wire  _GEN_7658 = io_op_bits_active_vidiv ? _GEN_6994 : _GEN_5240; // @[sequencer-master.scala 643:40]
  wire  _GEN_7659 = io_op_bits_active_vidiv ? _GEN_6995 : _GEN_5241; // @[sequencer-master.scala 643:40]
  wire  _GEN_7660 = io_op_bits_active_vidiv ? _GEN_6996 : _GEN_5242; // @[sequencer-master.scala 643:40]
  wire  _GEN_7661 = io_op_bits_active_vidiv ? _GEN_6997 : _GEN_5243; // @[sequencer-master.scala 643:40]
  wire  _GEN_7662 = io_op_bits_active_vidiv ? _GEN_6998 : _GEN_5244; // @[sequencer-master.scala 643:40]
  wire  _GEN_7663 = io_op_bits_active_vidiv ? _GEN_6999 : _GEN_5245; // @[sequencer-master.scala 643:40]
  wire  _GEN_7664 = io_op_bits_active_vidiv ? _GEN_7000 : _GEN_5246; // @[sequencer-master.scala 643:40]
  wire  _GEN_7665 = io_op_bits_active_vidiv ? _GEN_7001 : _GEN_5247; // @[sequencer-master.scala 643:40]
  wire  _GEN_7666 = io_op_bits_active_vidiv ? _GEN_7002 : _GEN_5248; // @[sequencer-master.scala 643:40]
  wire  _GEN_7667 = io_op_bits_active_vidiv ? _GEN_7003 : _GEN_5249; // @[sequencer-master.scala 643:40]
  wire  _GEN_7668 = io_op_bits_active_vidiv ? _GEN_7004 : _GEN_5250; // @[sequencer-master.scala 643:40]
  wire  _GEN_7669 = io_op_bits_active_vidiv ? _GEN_7005 : _GEN_5251; // @[sequencer-master.scala 643:40]
  wire  _GEN_7670 = io_op_bits_active_vidiv ? _GEN_7006 : _GEN_5252; // @[sequencer-master.scala 643:40]
  wire  _GEN_7671 = io_op_bits_active_vidiv ? _GEN_7007 : _GEN_5253; // @[sequencer-master.scala 643:40]
  wire  _GEN_7672 = io_op_bits_active_vidiv ? _GEN_7008 : _GEN_5254; // @[sequencer-master.scala 643:40]
  wire  _GEN_7673 = io_op_bits_active_vidiv ? _GEN_7009 : _GEN_5255; // @[sequencer-master.scala 643:40]
  wire  _GEN_7674 = io_op_bits_active_vidiv ? _GEN_7010 : _GEN_5256; // @[sequencer-master.scala 643:40]
  wire  _GEN_7675 = io_op_bits_active_vidiv ? _GEN_7011 : _GEN_5257; // @[sequencer-master.scala 643:40]
  wire  _GEN_7676 = io_op_bits_active_vidiv ? _GEN_7012 : _GEN_5258; // @[sequencer-master.scala 643:40]
  wire  _GEN_7677 = io_op_bits_active_vidiv ? _GEN_7013 : _GEN_5259; // @[sequencer-master.scala 643:40]
  wire  _GEN_7678 = io_op_bits_active_vidiv ? _GEN_7014 : _GEN_5260; // @[sequencer-master.scala 643:40]
  wire  _GEN_7679 = io_op_bits_active_vidiv ? _GEN_7015 : _GEN_5261; // @[sequencer-master.scala 643:40]
  wire  _GEN_7680 = io_op_bits_active_vidiv ? _GEN_7016 : _GEN_5262; // @[sequencer-master.scala 643:40]
  wire  _GEN_7681 = io_op_bits_active_vidiv ? _GEN_7017 : _GEN_5263; // @[sequencer-master.scala 643:40]
  wire  _GEN_7682 = io_op_bits_active_vidiv ? _GEN_7018 : _GEN_5264; // @[sequencer-master.scala 643:40]
  wire  _GEN_7683 = io_op_bits_active_vidiv ? _GEN_7019 : _GEN_5265; // @[sequencer-master.scala 643:40]
  wire  _GEN_7684 = io_op_bits_active_vidiv ? _GEN_7020 : _GEN_5266; // @[sequencer-master.scala 643:40]
  wire  _GEN_7685 = io_op_bits_active_vidiv ? _GEN_7021 : _GEN_5267; // @[sequencer-master.scala 643:40]
  wire  _GEN_7686 = io_op_bits_active_vidiv ? _GEN_7318 : _GEN_5268; // @[sequencer-master.scala 643:40]
  wire  _GEN_7687 = io_op_bits_active_vidiv ? _GEN_7319 : _GEN_5269; // @[sequencer-master.scala 643:40]
  wire  _GEN_7688 = io_op_bits_active_vidiv ? _GEN_7320 : _GEN_5270; // @[sequencer-master.scala 643:40]
  wire  _GEN_7689 = io_op_bits_active_vidiv ? _GEN_7321 : _GEN_5271; // @[sequencer-master.scala 643:40]
  wire  _GEN_7690 = io_op_bits_active_vidiv ? _GEN_7322 : _GEN_5272; // @[sequencer-master.scala 643:40]
  wire  _GEN_7691 = io_op_bits_active_vidiv ? _GEN_7323 : _GEN_5273; // @[sequencer-master.scala 643:40]
  wire  _GEN_7692 = io_op_bits_active_vidiv ? _GEN_7324 : _GEN_5274; // @[sequencer-master.scala 643:40]
  wire  _GEN_7693 = io_op_bits_active_vidiv ? _GEN_7325 : _GEN_5275; // @[sequencer-master.scala 643:40]
  wire  _GEN_7694 = io_op_bits_active_vidiv ? _GEN_7030 : _GEN_5276; // @[sequencer-master.scala 643:40]
  wire  _GEN_7695 = io_op_bits_active_vidiv ? _GEN_7031 : _GEN_5277; // @[sequencer-master.scala 643:40]
  wire  _GEN_7696 = io_op_bits_active_vidiv ? _GEN_7032 : _GEN_5278; // @[sequencer-master.scala 643:40]
  wire  _GEN_7697 = io_op_bits_active_vidiv ? _GEN_7033 : _GEN_5279; // @[sequencer-master.scala 643:40]
  wire  _GEN_7698 = io_op_bits_active_vidiv ? _GEN_7034 : _GEN_5280; // @[sequencer-master.scala 643:40]
  wire  _GEN_7699 = io_op_bits_active_vidiv ? _GEN_7035 : _GEN_5281; // @[sequencer-master.scala 643:40]
  wire  _GEN_7700 = io_op_bits_active_vidiv ? _GEN_7036 : _GEN_5282; // @[sequencer-master.scala 643:40]
  wire  _GEN_7701 = io_op_bits_active_vidiv ? _GEN_7037 : _GEN_5283; // @[sequencer-master.scala 643:40]
  wire  _GEN_7702 = io_op_bits_active_vidiv ? _GEN_7038 : _GEN_5284; // @[sequencer-master.scala 643:40]
  wire  _GEN_7703 = io_op_bits_active_vidiv ? _GEN_7039 : _GEN_5285; // @[sequencer-master.scala 643:40]
  wire  _GEN_7704 = io_op_bits_active_vidiv ? _GEN_7040 : _GEN_5286; // @[sequencer-master.scala 643:40]
  wire  _GEN_7705 = io_op_bits_active_vidiv ? _GEN_7041 : _GEN_5287; // @[sequencer-master.scala 643:40]
  wire  _GEN_7706 = io_op_bits_active_vidiv ? _GEN_7042 : _GEN_5288; // @[sequencer-master.scala 643:40]
  wire  _GEN_7707 = io_op_bits_active_vidiv ? _GEN_7043 : _GEN_5289; // @[sequencer-master.scala 643:40]
  wire  _GEN_7708 = io_op_bits_active_vidiv ? _GEN_7044 : _GEN_5290; // @[sequencer-master.scala 643:40]
  wire  _GEN_7709 = io_op_bits_active_vidiv ? _GEN_7045 : _GEN_5291; // @[sequencer-master.scala 643:40]
  wire  _GEN_7710 = io_op_bits_active_vidiv ? _GEN_7366 : _GEN_5292; // @[sequencer-master.scala 643:40]
  wire  _GEN_7711 = io_op_bits_active_vidiv ? _GEN_7367 : _GEN_5293; // @[sequencer-master.scala 643:40]
  wire  _GEN_7712 = io_op_bits_active_vidiv ? _GEN_7368 : _GEN_5294; // @[sequencer-master.scala 643:40]
  wire  _GEN_7713 = io_op_bits_active_vidiv ? _GEN_7369 : _GEN_5295; // @[sequencer-master.scala 643:40]
  wire  _GEN_7714 = io_op_bits_active_vidiv ? _GEN_7370 : _GEN_5296; // @[sequencer-master.scala 643:40]
  wire  _GEN_7715 = io_op_bits_active_vidiv ? _GEN_7371 : _GEN_5297; // @[sequencer-master.scala 643:40]
  wire  _GEN_7716 = io_op_bits_active_vidiv ? _GEN_7372 : _GEN_5298; // @[sequencer-master.scala 643:40]
  wire  _GEN_7717 = io_op_bits_active_vidiv ? _GEN_7373 : _GEN_5299; // @[sequencer-master.scala 643:40]
  wire  _GEN_7718 = io_op_bits_active_vidiv ? _GEN_7494 : _GEN_5300; // @[sequencer-master.scala 643:40]
  wire  _GEN_7719 = io_op_bits_active_vidiv ? _GEN_7495 : _GEN_5301; // @[sequencer-master.scala 643:40]
  wire  _GEN_7720 = io_op_bits_active_vidiv ? _GEN_7496 : _GEN_5302; // @[sequencer-master.scala 643:40]
  wire  _GEN_7721 = io_op_bits_active_vidiv ? _GEN_7497 : _GEN_5303; // @[sequencer-master.scala 643:40]
  wire  _GEN_7722 = io_op_bits_active_vidiv ? _GEN_7498 : _GEN_5304; // @[sequencer-master.scala 643:40]
  wire  _GEN_7723 = io_op_bits_active_vidiv ? _GEN_7499 : _GEN_5305; // @[sequencer-master.scala 643:40]
  wire  _GEN_7724 = io_op_bits_active_vidiv ? _GEN_7500 : _GEN_5306; // @[sequencer-master.scala 643:40]
  wire  _GEN_7725 = io_op_bits_active_vidiv ? _GEN_7501 : _GEN_5307; // @[sequencer-master.scala 643:40]
  wire  _GEN_7726 = io_op_bits_active_vidiv ? _GEN_7062 : _GEN_5308; // @[sequencer-master.scala 643:40]
  wire  _GEN_7727 = io_op_bits_active_vidiv ? _GEN_7063 : _GEN_5309; // @[sequencer-master.scala 643:40]
  wire  _GEN_7728 = io_op_bits_active_vidiv ? _GEN_7064 : _GEN_5310; // @[sequencer-master.scala 643:40]
  wire  _GEN_7729 = io_op_bits_active_vidiv ? _GEN_7065 : _GEN_5311; // @[sequencer-master.scala 643:40]
  wire  _GEN_7730 = io_op_bits_active_vidiv ? _GEN_7066 : _GEN_5312; // @[sequencer-master.scala 643:40]
  wire  _GEN_7731 = io_op_bits_active_vidiv ? _GEN_7067 : _GEN_5313; // @[sequencer-master.scala 643:40]
  wire  _GEN_7732 = io_op_bits_active_vidiv ? _GEN_7068 : _GEN_5314; // @[sequencer-master.scala 643:40]
  wire  _GEN_7733 = io_op_bits_active_vidiv ? _GEN_7069 : _GEN_5315; // @[sequencer-master.scala 643:40]
  wire  _GEN_7734 = io_op_bits_active_vidiv ? _GEN_7382 : _GEN_5316; // @[sequencer-master.scala 643:40]
  wire  _GEN_7735 = io_op_bits_active_vidiv ? _GEN_7383 : _GEN_5317; // @[sequencer-master.scala 643:40]
  wire  _GEN_7736 = io_op_bits_active_vidiv ? _GEN_7384 : _GEN_5318; // @[sequencer-master.scala 643:40]
  wire  _GEN_7737 = io_op_bits_active_vidiv ? _GEN_7385 : _GEN_5319; // @[sequencer-master.scala 643:40]
  wire  _GEN_7738 = io_op_bits_active_vidiv ? _GEN_7386 : _GEN_5320; // @[sequencer-master.scala 643:40]
  wire  _GEN_7739 = io_op_bits_active_vidiv ? _GEN_7387 : _GEN_5321; // @[sequencer-master.scala 643:40]
  wire  _GEN_7740 = io_op_bits_active_vidiv ? _GEN_7388 : _GEN_5322; // @[sequencer-master.scala 643:40]
  wire  _GEN_7741 = io_op_bits_active_vidiv ? _GEN_7389 : _GEN_5323; // @[sequencer-master.scala 643:40]
  wire  _GEN_7742 = io_op_bits_active_vidiv ? _GEN_7510 : _GEN_5324; // @[sequencer-master.scala 643:40]
  wire  _GEN_7743 = io_op_bits_active_vidiv ? _GEN_7511 : _GEN_5325; // @[sequencer-master.scala 643:40]
  wire  _GEN_7744 = io_op_bits_active_vidiv ? _GEN_7512 : _GEN_5326; // @[sequencer-master.scala 643:40]
  wire  _GEN_7745 = io_op_bits_active_vidiv ? _GEN_7513 : _GEN_5327; // @[sequencer-master.scala 643:40]
  wire  _GEN_7746 = io_op_bits_active_vidiv ? _GEN_7514 : _GEN_5328; // @[sequencer-master.scala 643:40]
  wire  _GEN_7747 = io_op_bits_active_vidiv ? _GEN_7515 : _GEN_5329; // @[sequencer-master.scala 643:40]
  wire  _GEN_7748 = io_op_bits_active_vidiv ? _GEN_7516 : _GEN_5330; // @[sequencer-master.scala 643:40]
  wire  _GEN_7749 = io_op_bits_active_vidiv ? _GEN_7517 : _GEN_5331; // @[sequencer-master.scala 643:40]
  wire  _GEN_7750 = io_op_bits_active_vidiv ? _GEN_7086 : _GEN_5332; // @[sequencer-master.scala 643:40]
  wire  _GEN_7751 = io_op_bits_active_vidiv ? _GEN_7087 : _GEN_5333; // @[sequencer-master.scala 643:40]
  wire  _GEN_7752 = io_op_bits_active_vidiv ? _GEN_7088 : _GEN_5334; // @[sequencer-master.scala 643:40]
  wire  _GEN_7753 = io_op_bits_active_vidiv ? _GEN_7089 : _GEN_5335; // @[sequencer-master.scala 643:40]
  wire  _GEN_7754 = io_op_bits_active_vidiv ? _GEN_7090 : _GEN_5336; // @[sequencer-master.scala 643:40]
  wire  _GEN_7755 = io_op_bits_active_vidiv ? _GEN_7091 : _GEN_5337; // @[sequencer-master.scala 643:40]
  wire  _GEN_7756 = io_op_bits_active_vidiv ? _GEN_7092 : _GEN_5338; // @[sequencer-master.scala 643:40]
  wire  _GEN_7757 = io_op_bits_active_vidiv ? _GEN_7093 : _GEN_5339; // @[sequencer-master.scala 643:40]
  wire  _GEN_7758 = io_op_bits_active_vidiv ? _GEN_7398 : _GEN_5340; // @[sequencer-master.scala 643:40]
  wire  _GEN_7759 = io_op_bits_active_vidiv ? _GEN_7399 : _GEN_5341; // @[sequencer-master.scala 643:40]
  wire  _GEN_7760 = io_op_bits_active_vidiv ? _GEN_7400 : _GEN_5342; // @[sequencer-master.scala 643:40]
  wire  _GEN_7761 = io_op_bits_active_vidiv ? _GEN_7401 : _GEN_5343; // @[sequencer-master.scala 643:40]
  wire  _GEN_7762 = io_op_bits_active_vidiv ? _GEN_7402 : _GEN_5344; // @[sequencer-master.scala 643:40]
  wire  _GEN_7763 = io_op_bits_active_vidiv ? _GEN_7403 : _GEN_5345; // @[sequencer-master.scala 643:40]
  wire  _GEN_7764 = io_op_bits_active_vidiv ? _GEN_7404 : _GEN_5346; // @[sequencer-master.scala 643:40]
  wire  _GEN_7765 = io_op_bits_active_vidiv ? _GEN_7405 : _GEN_5347; // @[sequencer-master.scala 643:40]
  wire  _GEN_7766 = io_op_bits_active_vidiv ? _GEN_7526 : _GEN_5348; // @[sequencer-master.scala 643:40]
  wire  _GEN_7767 = io_op_bits_active_vidiv ? _GEN_7527 : _GEN_5349; // @[sequencer-master.scala 643:40]
  wire  _GEN_7768 = io_op_bits_active_vidiv ? _GEN_7528 : _GEN_5350; // @[sequencer-master.scala 643:40]
  wire  _GEN_7769 = io_op_bits_active_vidiv ? _GEN_7529 : _GEN_5351; // @[sequencer-master.scala 643:40]
  wire  _GEN_7770 = io_op_bits_active_vidiv ? _GEN_7530 : _GEN_5352; // @[sequencer-master.scala 643:40]
  wire  _GEN_7771 = io_op_bits_active_vidiv ? _GEN_7531 : _GEN_5353; // @[sequencer-master.scala 643:40]
  wire  _GEN_7772 = io_op_bits_active_vidiv ? _GEN_7532 : _GEN_5354; // @[sequencer-master.scala 643:40]
  wire  _GEN_7773 = io_op_bits_active_vidiv ? _GEN_7533 : _GEN_5355; // @[sequencer-master.scala 643:40]
  wire  _GEN_7774 = io_op_bits_active_vidiv ? _GEN_7110 : _GEN_5356; // @[sequencer-master.scala 643:40]
  wire  _GEN_7775 = io_op_bits_active_vidiv ? _GEN_7111 : _GEN_5357; // @[sequencer-master.scala 643:40]
  wire  _GEN_7776 = io_op_bits_active_vidiv ? _GEN_7112 : _GEN_5358; // @[sequencer-master.scala 643:40]
  wire  _GEN_7777 = io_op_bits_active_vidiv ? _GEN_7113 : _GEN_5359; // @[sequencer-master.scala 643:40]
  wire  _GEN_7778 = io_op_bits_active_vidiv ? _GEN_7114 : _GEN_5360; // @[sequencer-master.scala 643:40]
  wire  _GEN_7779 = io_op_bits_active_vidiv ? _GEN_7115 : _GEN_5361; // @[sequencer-master.scala 643:40]
  wire  _GEN_7780 = io_op_bits_active_vidiv ? _GEN_7116 : _GEN_5362; // @[sequencer-master.scala 643:40]
  wire  _GEN_7781 = io_op_bits_active_vidiv ? _GEN_7117 : _GEN_5363; // @[sequencer-master.scala 643:40]
  wire  _GEN_7782 = io_op_bits_active_vidiv ? _GEN_7414 : _GEN_5364; // @[sequencer-master.scala 643:40]
  wire  _GEN_7783 = io_op_bits_active_vidiv ? _GEN_7415 : _GEN_5365; // @[sequencer-master.scala 643:40]
  wire  _GEN_7784 = io_op_bits_active_vidiv ? _GEN_7416 : _GEN_5366; // @[sequencer-master.scala 643:40]
  wire  _GEN_7785 = io_op_bits_active_vidiv ? _GEN_7417 : _GEN_5367; // @[sequencer-master.scala 643:40]
  wire  _GEN_7786 = io_op_bits_active_vidiv ? _GEN_7418 : _GEN_5368; // @[sequencer-master.scala 643:40]
  wire  _GEN_7787 = io_op_bits_active_vidiv ? _GEN_7419 : _GEN_5369; // @[sequencer-master.scala 643:40]
  wire  _GEN_7788 = io_op_bits_active_vidiv ? _GEN_7420 : _GEN_5370; // @[sequencer-master.scala 643:40]
  wire  _GEN_7789 = io_op_bits_active_vidiv ? _GEN_7421 : _GEN_5371; // @[sequencer-master.scala 643:40]
  wire  _GEN_7790 = io_op_bits_active_vidiv ? _GEN_7542 : _GEN_5372; // @[sequencer-master.scala 643:40]
  wire  _GEN_7791 = io_op_bits_active_vidiv ? _GEN_7543 : _GEN_5373; // @[sequencer-master.scala 643:40]
  wire  _GEN_7792 = io_op_bits_active_vidiv ? _GEN_7544 : _GEN_5374; // @[sequencer-master.scala 643:40]
  wire  _GEN_7793 = io_op_bits_active_vidiv ? _GEN_7545 : _GEN_5375; // @[sequencer-master.scala 643:40]
  wire  _GEN_7794 = io_op_bits_active_vidiv ? _GEN_7546 : _GEN_5376; // @[sequencer-master.scala 643:40]
  wire  _GEN_7795 = io_op_bits_active_vidiv ? _GEN_7547 : _GEN_5377; // @[sequencer-master.scala 643:40]
  wire  _GEN_7796 = io_op_bits_active_vidiv ? _GEN_7548 : _GEN_5378; // @[sequencer-master.scala 643:40]
  wire  _GEN_7797 = io_op_bits_active_vidiv ? _GEN_7549 : _GEN_5379; // @[sequencer-master.scala 643:40]
  wire  _GEN_7798 = io_op_bits_active_vidiv ? _GEN_7134 : _GEN_5380; // @[sequencer-master.scala 643:40]
  wire  _GEN_7799 = io_op_bits_active_vidiv ? _GEN_7135 : _GEN_5381; // @[sequencer-master.scala 643:40]
  wire  _GEN_7800 = io_op_bits_active_vidiv ? _GEN_7136 : _GEN_5382; // @[sequencer-master.scala 643:40]
  wire  _GEN_7801 = io_op_bits_active_vidiv ? _GEN_7137 : _GEN_5383; // @[sequencer-master.scala 643:40]
  wire  _GEN_7802 = io_op_bits_active_vidiv ? _GEN_7138 : _GEN_5384; // @[sequencer-master.scala 643:40]
  wire  _GEN_7803 = io_op_bits_active_vidiv ? _GEN_7139 : _GEN_5385; // @[sequencer-master.scala 643:40]
  wire  _GEN_7804 = io_op_bits_active_vidiv ? _GEN_7140 : _GEN_5386; // @[sequencer-master.scala 643:40]
  wire  _GEN_7805 = io_op_bits_active_vidiv ? _GEN_7141 : _GEN_5387; // @[sequencer-master.scala 643:40]
  wire  _GEN_7806 = io_op_bits_active_vidiv ? _GEN_7430 : _GEN_5388; // @[sequencer-master.scala 643:40]
  wire  _GEN_7807 = io_op_bits_active_vidiv ? _GEN_7431 : _GEN_5389; // @[sequencer-master.scala 643:40]
  wire  _GEN_7808 = io_op_bits_active_vidiv ? _GEN_7432 : _GEN_5390; // @[sequencer-master.scala 643:40]
  wire  _GEN_7809 = io_op_bits_active_vidiv ? _GEN_7433 : _GEN_5391; // @[sequencer-master.scala 643:40]
  wire  _GEN_7810 = io_op_bits_active_vidiv ? _GEN_7434 : _GEN_5392; // @[sequencer-master.scala 643:40]
  wire  _GEN_7811 = io_op_bits_active_vidiv ? _GEN_7435 : _GEN_5393; // @[sequencer-master.scala 643:40]
  wire  _GEN_7812 = io_op_bits_active_vidiv ? _GEN_7436 : _GEN_5394; // @[sequencer-master.scala 643:40]
  wire  _GEN_7813 = io_op_bits_active_vidiv ? _GEN_7437 : _GEN_5395; // @[sequencer-master.scala 643:40]
  wire  _GEN_7814 = io_op_bits_active_vidiv ? _GEN_7558 : _GEN_5396; // @[sequencer-master.scala 643:40]
  wire  _GEN_7815 = io_op_bits_active_vidiv ? _GEN_7559 : _GEN_5397; // @[sequencer-master.scala 643:40]
  wire  _GEN_7816 = io_op_bits_active_vidiv ? _GEN_7560 : _GEN_5398; // @[sequencer-master.scala 643:40]
  wire  _GEN_7817 = io_op_bits_active_vidiv ? _GEN_7561 : _GEN_5399; // @[sequencer-master.scala 643:40]
  wire  _GEN_7818 = io_op_bits_active_vidiv ? _GEN_7562 : _GEN_5400; // @[sequencer-master.scala 643:40]
  wire  _GEN_7819 = io_op_bits_active_vidiv ? _GEN_7563 : _GEN_5401; // @[sequencer-master.scala 643:40]
  wire  _GEN_7820 = io_op_bits_active_vidiv ? _GEN_7564 : _GEN_5402; // @[sequencer-master.scala 643:40]
  wire  _GEN_7821 = io_op_bits_active_vidiv ? _GEN_7565 : _GEN_5403; // @[sequencer-master.scala 643:40]
  wire  _GEN_7822 = io_op_bits_active_vidiv ? _GEN_7158 : _GEN_5404; // @[sequencer-master.scala 643:40]
  wire  _GEN_7823 = io_op_bits_active_vidiv ? _GEN_7159 : _GEN_5405; // @[sequencer-master.scala 643:40]
  wire  _GEN_7824 = io_op_bits_active_vidiv ? _GEN_7160 : _GEN_5406; // @[sequencer-master.scala 643:40]
  wire  _GEN_7825 = io_op_bits_active_vidiv ? _GEN_7161 : _GEN_5407; // @[sequencer-master.scala 643:40]
  wire  _GEN_7826 = io_op_bits_active_vidiv ? _GEN_7162 : _GEN_5408; // @[sequencer-master.scala 643:40]
  wire  _GEN_7827 = io_op_bits_active_vidiv ? _GEN_7163 : _GEN_5409; // @[sequencer-master.scala 643:40]
  wire  _GEN_7828 = io_op_bits_active_vidiv ? _GEN_7164 : _GEN_5410; // @[sequencer-master.scala 643:40]
  wire  _GEN_7829 = io_op_bits_active_vidiv ? _GEN_7165 : _GEN_5411; // @[sequencer-master.scala 643:40]
  wire  _GEN_7830 = io_op_bits_active_vidiv ? _GEN_7446 : _GEN_5412; // @[sequencer-master.scala 643:40]
  wire  _GEN_7831 = io_op_bits_active_vidiv ? _GEN_7447 : _GEN_5413; // @[sequencer-master.scala 643:40]
  wire  _GEN_7832 = io_op_bits_active_vidiv ? _GEN_7448 : _GEN_5414; // @[sequencer-master.scala 643:40]
  wire  _GEN_7833 = io_op_bits_active_vidiv ? _GEN_7449 : _GEN_5415; // @[sequencer-master.scala 643:40]
  wire  _GEN_7834 = io_op_bits_active_vidiv ? _GEN_7450 : _GEN_5416; // @[sequencer-master.scala 643:40]
  wire  _GEN_7835 = io_op_bits_active_vidiv ? _GEN_7451 : _GEN_5417; // @[sequencer-master.scala 643:40]
  wire  _GEN_7836 = io_op_bits_active_vidiv ? _GEN_7452 : _GEN_5418; // @[sequencer-master.scala 643:40]
  wire  _GEN_7837 = io_op_bits_active_vidiv ? _GEN_7453 : _GEN_5419; // @[sequencer-master.scala 643:40]
  wire  _GEN_7838 = io_op_bits_active_vidiv ? _GEN_7574 : _GEN_5420; // @[sequencer-master.scala 643:40]
  wire  _GEN_7839 = io_op_bits_active_vidiv ? _GEN_7575 : _GEN_5421; // @[sequencer-master.scala 643:40]
  wire  _GEN_7840 = io_op_bits_active_vidiv ? _GEN_7576 : _GEN_5422; // @[sequencer-master.scala 643:40]
  wire  _GEN_7841 = io_op_bits_active_vidiv ? _GEN_7577 : _GEN_5423; // @[sequencer-master.scala 643:40]
  wire  _GEN_7842 = io_op_bits_active_vidiv ? _GEN_7578 : _GEN_5424; // @[sequencer-master.scala 643:40]
  wire  _GEN_7843 = io_op_bits_active_vidiv ? _GEN_7579 : _GEN_5425; // @[sequencer-master.scala 643:40]
  wire  _GEN_7844 = io_op_bits_active_vidiv ? _GEN_7580 : _GEN_5426; // @[sequencer-master.scala 643:40]
  wire  _GEN_7845 = io_op_bits_active_vidiv ? _GEN_7581 : _GEN_5427; // @[sequencer-master.scala 643:40]
  wire  _GEN_7846 = io_op_bits_active_vidiv ? _GEN_7182 : _GEN_5428; // @[sequencer-master.scala 643:40]
  wire  _GEN_7847 = io_op_bits_active_vidiv ? _GEN_7183 : _GEN_5429; // @[sequencer-master.scala 643:40]
  wire  _GEN_7848 = io_op_bits_active_vidiv ? _GEN_7184 : _GEN_5430; // @[sequencer-master.scala 643:40]
  wire  _GEN_7849 = io_op_bits_active_vidiv ? _GEN_7185 : _GEN_5431; // @[sequencer-master.scala 643:40]
  wire  _GEN_7850 = io_op_bits_active_vidiv ? _GEN_7186 : _GEN_5432; // @[sequencer-master.scala 643:40]
  wire  _GEN_7851 = io_op_bits_active_vidiv ? _GEN_7187 : _GEN_5433; // @[sequencer-master.scala 643:40]
  wire  _GEN_7852 = io_op_bits_active_vidiv ? _GEN_7188 : _GEN_5434; // @[sequencer-master.scala 643:40]
  wire  _GEN_7853 = io_op_bits_active_vidiv ? _GEN_7189 : _GEN_5435; // @[sequencer-master.scala 643:40]
  wire  _GEN_7854 = io_op_bits_active_vidiv ? _GEN_7462 : _GEN_5436; // @[sequencer-master.scala 643:40]
  wire  _GEN_7855 = io_op_bits_active_vidiv ? _GEN_7463 : _GEN_5437; // @[sequencer-master.scala 643:40]
  wire  _GEN_7856 = io_op_bits_active_vidiv ? _GEN_7464 : _GEN_5438; // @[sequencer-master.scala 643:40]
  wire  _GEN_7857 = io_op_bits_active_vidiv ? _GEN_7465 : _GEN_5439; // @[sequencer-master.scala 643:40]
  wire  _GEN_7858 = io_op_bits_active_vidiv ? _GEN_7466 : _GEN_5440; // @[sequencer-master.scala 643:40]
  wire  _GEN_7859 = io_op_bits_active_vidiv ? _GEN_7467 : _GEN_5441; // @[sequencer-master.scala 643:40]
  wire  _GEN_7860 = io_op_bits_active_vidiv ? _GEN_7468 : _GEN_5442; // @[sequencer-master.scala 643:40]
  wire  _GEN_7861 = io_op_bits_active_vidiv ? _GEN_7469 : _GEN_5443; // @[sequencer-master.scala 643:40]
  wire  _GEN_7862 = io_op_bits_active_vidiv ? _GEN_7590 : _GEN_5444; // @[sequencer-master.scala 643:40]
  wire  _GEN_7863 = io_op_bits_active_vidiv ? _GEN_7591 : _GEN_5445; // @[sequencer-master.scala 643:40]
  wire  _GEN_7864 = io_op_bits_active_vidiv ? _GEN_7592 : _GEN_5446; // @[sequencer-master.scala 643:40]
  wire  _GEN_7865 = io_op_bits_active_vidiv ? _GEN_7593 : _GEN_5447; // @[sequencer-master.scala 643:40]
  wire  _GEN_7866 = io_op_bits_active_vidiv ? _GEN_7594 : _GEN_5448; // @[sequencer-master.scala 643:40]
  wire  _GEN_7867 = io_op_bits_active_vidiv ? _GEN_7595 : _GEN_5449; // @[sequencer-master.scala 643:40]
  wire  _GEN_7868 = io_op_bits_active_vidiv ? _GEN_7596 : _GEN_5450; // @[sequencer-master.scala 643:40]
  wire  _GEN_7869 = io_op_bits_active_vidiv ? _GEN_7597 : _GEN_5451; // @[sequencer-master.scala 643:40]
  wire  _GEN_7870 = io_op_bits_active_vidiv ? _GEN_7206 : _GEN_5452; // @[sequencer-master.scala 643:40]
  wire  _GEN_7871 = io_op_bits_active_vidiv ? _GEN_7207 : _GEN_5453; // @[sequencer-master.scala 643:40]
  wire  _GEN_7872 = io_op_bits_active_vidiv ? _GEN_7208 : _GEN_5454; // @[sequencer-master.scala 643:40]
  wire  _GEN_7873 = io_op_bits_active_vidiv ? _GEN_7209 : _GEN_5455; // @[sequencer-master.scala 643:40]
  wire  _GEN_7874 = io_op_bits_active_vidiv ? _GEN_7210 : _GEN_5456; // @[sequencer-master.scala 643:40]
  wire  _GEN_7875 = io_op_bits_active_vidiv ? _GEN_7211 : _GEN_5457; // @[sequencer-master.scala 643:40]
  wire  _GEN_7876 = io_op_bits_active_vidiv ? _GEN_7212 : _GEN_5458; // @[sequencer-master.scala 643:40]
  wire  _GEN_7877 = io_op_bits_active_vidiv ? _GEN_7213 : _GEN_5459; // @[sequencer-master.scala 643:40]
  wire  _GEN_7878 = io_op_bits_active_vidiv ? _GEN_7478 : _GEN_5460; // @[sequencer-master.scala 643:40]
  wire  _GEN_7879 = io_op_bits_active_vidiv ? _GEN_7479 : _GEN_5461; // @[sequencer-master.scala 643:40]
  wire  _GEN_7880 = io_op_bits_active_vidiv ? _GEN_7480 : _GEN_5462; // @[sequencer-master.scala 643:40]
  wire  _GEN_7881 = io_op_bits_active_vidiv ? _GEN_7481 : _GEN_5463; // @[sequencer-master.scala 643:40]
  wire  _GEN_7882 = io_op_bits_active_vidiv ? _GEN_7482 : _GEN_5464; // @[sequencer-master.scala 643:40]
  wire  _GEN_7883 = io_op_bits_active_vidiv ? _GEN_7483 : _GEN_5465; // @[sequencer-master.scala 643:40]
  wire  _GEN_7884 = io_op_bits_active_vidiv ? _GEN_7484 : _GEN_5466; // @[sequencer-master.scala 643:40]
  wire  _GEN_7885 = io_op_bits_active_vidiv ? _GEN_7485 : _GEN_5467; // @[sequencer-master.scala 643:40]
  wire  _GEN_7886 = io_op_bits_active_vidiv ? _GEN_7606 : _GEN_5468; // @[sequencer-master.scala 643:40]
  wire  _GEN_7887 = io_op_bits_active_vidiv ? _GEN_7607 : _GEN_5469; // @[sequencer-master.scala 643:40]
  wire  _GEN_7888 = io_op_bits_active_vidiv ? _GEN_7608 : _GEN_5470; // @[sequencer-master.scala 643:40]
  wire  _GEN_7889 = io_op_bits_active_vidiv ? _GEN_7609 : _GEN_5471; // @[sequencer-master.scala 643:40]
  wire  _GEN_7890 = io_op_bits_active_vidiv ? _GEN_7610 : _GEN_5472; // @[sequencer-master.scala 643:40]
  wire  _GEN_7891 = io_op_bits_active_vidiv ? _GEN_7611 : _GEN_5473; // @[sequencer-master.scala 643:40]
  wire  _GEN_7892 = io_op_bits_active_vidiv ? _GEN_7612 : _GEN_5474; // @[sequencer-master.scala 643:40]
  wire  _GEN_7893 = io_op_bits_active_vidiv ? _GEN_7613 : _GEN_5475; // @[sequencer-master.scala 643:40]
  wire  _GEN_7894 = io_op_bits_active_vidiv ? _GEN_7230 : _GEN_5476; // @[sequencer-master.scala 643:40]
  wire  _GEN_7895 = io_op_bits_active_vidiv ? _GEN_7231 : _GEN_5477; // @[sequencer-master.scala 643:40]
  wire  _GEN_7896 = io_op_bits_active_vidiv ? _GEN_7232 : _GEN_5478; // @[sequencer-master.scala 643:40]
  wire  _GEN_7897 = io_op_bits_active_vidiv ? _GEN_7233 : _GEN_5479; // @[sequencer-master.scala 643:40]
  wire  _GEN_7898 = io_op_bits_active_vidiv ? _GEN_7234 : _GEN_5480; // @[sequencer-master.scala 643:40]
  wire  _GEN_7899 = io_op_bits_active_vidiv ? _GEN_7235 : _GEN_5481; // @[sequencer-master.scala 643:40]
  wire  _GEN_7900 = io_op_bits_active_vidiv ? _GEN_7236 : _GEN_5482; // @[sequencer-master.scala 643:40]
  wire  _GEN_7901 = io_op_bits_active_vidiv ? _GEN_7237 : _GEN_5483; // @[sequencer-master.scala 643:40]
  wire  _GEN_7910 = io_op_bits_active_vidiv ? _GEN_5974 : e_0_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7911 = io_op_bits_active_vidiv ? _GEN_5975 : e_1_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7912 = io_op_bits_active_vidiv ? _GEN_5976 : e_2_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7913 = io_op_bits_active_vidiv ? _GEN_5977 : e_3_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7914 = io_op_bits_active_vidiv ? _GEN_5978 : e_4_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7915 = io_op_bits_active_vidiv ? _GEN_5979 : e_5_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7916 = io_op_bits_active_vidiv ? _GEN_5980 : e_6_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_7917 = io_op_bits_active_vidiv ? _GEN_5981 : e_7_active_vqu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire [9:0] _GEN_7918 = io_op_bits_active_vidiv ? _GEN_7254 : _GEN_5500; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7919 = io_op_bits_active_vidiv ? _GEN_7255 : _GEN_5501; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7920 = io_op_bits_active_vidiv ? _GEN_7256 : _GEN_5502; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7921 = io_op_bits_active_vidiv ? _GEN_7257 : _GEN_5503; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7922 = io_op_bits_active_vidiv ? _GEN_7258 : _GEN_5504; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7923 = io_op_bits_active_vidiv ? _GEN_7259 : _GEN_5505; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7924 = io_op_bits_active_vidiv ? _GEN_7260 : _GEN_5506; // @[sequencer-master.scala 643:40]
  wire [9:0] _GEN_7925 = io_op_bits_active_vidiv ? _GEN_7261 : _GEN_5507; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7926 = io_op_bits_active_vidiv ? _GEN_6030 : _GEN_5508; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7927 = io_op_bits_active_vidiv ? _GEN_6031 : _GEN_5509; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7928 = io_op_bits_active_vidiv ? _GEN_6032 : _GEN_5510; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7929 = io_op_bits_active_vidiv ? _GEN_6033 : _GEN_5511; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7930 = io_op_bits_active_vidiv ? _GEN_6034 : _GEN_5512; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7931 = io_op_bits_active_vidiv ? _GEN_6035 : _GEN_5513; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7932 = io_op_bits_active_vidiv ? _GEN_6036 : _GEN_5514; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_7933 = io_op_bits_active_vidiv ? _GEN_6037 : _GEN_5515; // @[sequencer-master.scala 643:40]
  wire  _GEN_7934 = io_op_bits_active_vidiv ? _GEN_6046 : _GEN_5516; // @[sequencer-master.scala 643:40]
  wire  _GEN_7935 = io_op_bits_active_vidiv ? _GEN_6047 : _GEN_5517; // @[sequencer-master.scala 643:40]
  wire  _GEN_7936 = io_op_bits_active_vidiv ? _GEN_6048 : _GEN_5518; // @[sequencer-master.scala 643:40]
  wire  _GEN_7937 = io_op_bits_active_vidiv ? _GEN_6049 : _GEN_5519; // @[sequencer-master.scala 643:40]
  wire  _GEN_7938 = io_op_bits_active_vidiv ? _GEN_6050 : _GEN_5520; // @[sequencer-master.scala 643:40]
  wire  _GEN_7939 = io_op_bits_active_vidiv ? _GEN_6051 : _GEN_5521; // @[sequencer-master.scala 643:40]
  wire  _GEN_7940 = io_op_bits_active_vidiv ? _GEN_6052 : _GEN_5522; // @[sequencer-master.scala 643:40]
  wire  _GEN_7941 = io_op_bits_active_vidiv ? _GEN_6053 : _GEN_5523; // @[sequencer-master.scala 643:40]
  wire  _GEN_7942 = io_op_bits_active_vidiv ? _GEN_6054 : _GEN_5524; // @[sequencer-master.scala 643:40]
  wire  _GEN_7943 = io_op_bits_active_vidiv ? _GEN_6055 : _GEN_5525; // @[sequencer-master.scala 643:40]
  wire  _GEN_7944 = io_op_bits_active_vidiv ? _GEN_6056 : _GEN_5526; // @[sequencer-master.scala 643:40]
  wire  _GEN_7945 = io_op_bits_active_vidiv ? _GEN_6057 : _GEN_5527; // @[sequencer-master.scala 643:40]
  wire  _GEN_7946 = io_op_bits_active_vidiv ? _GEN_6058 : _GEN_5528; // @[sequencer-master.scala 643:40]
  wire  _GEN_7947 = io_op_bits_active_vidiv ? _GEN_6059 : _GEN_5529; // @[sequencer-master.scala 643:40]
  wire  _GEN_7948 = io_op_bits_active_vidiv ? _GEN_6060 : _GEN_5530; // @[sequencer-master.scala 643:40]
  wire  _GEN_7949 = io_op_bits_active_vidiv ? _GEN_6061 : _GEN_5531; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7950 = io_op_bits_active_vidiv ? _GEN_6062 : _GEN_5532; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7951 = io_op_bits_active_vidiv ? _GEN_6063 : _GEN_5533; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7952 = io_op_bits_active_vidiv ? _GEN_6064 : _GEN_5534; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7953 = io_op_bits_active_vidiv ? _GEN_6065 : _GEN_5535; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7954 = io_op_bits_active_vidiv ? _GEN_6066 : _GEN_5536; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7955 = io_op_bits_active_vidiv ? _GEN_6067 : _GEN_5537; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7956 = io_op_bits_active_vidiv ? _GEN_6068 : _GEN_5538; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7957 = io_op_bits_active_vidiv ? _GEN_6069 : _GEN_5539; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7958 = io_op_bits_active_vidiv ? _GEN_6262 : _GEN_5540; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7959 = io_op_bits_active_vidiv ? _GEN_6263 : _GEN_5541; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7960 = io_op_bits_active_vidiv ? _GEN_6264 : _GEN_5542; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7961 = io_op_bits_active_vidiv ? _GEN_6265 : _GEN_5543; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7962 = io_op_bits_active_vidiv ? _GEN_6266 : _GEN_5544; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7963 = io_op_bits_active_vidiv ? _GEN_6267 : _GEN_5545; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7964 = io_op_bits_active_vidiv ? _GEN_6268 : _GEN_5546; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7965 = io_op_bits_active_vidiv ? _GEN_6269 : _GEN_5547; // @[sequencer-master.scala 643:40]
  wire  _GEN_7966 = io_op_bits_active_vidiv ? _GEN_6278 : _GEN_5548; // @[sequencer-master.scala 643:40]
  wire  _GEN_7967 = io_op_bits_active_vidiv ? _GEN_6279 : _GEN_5549; // @[sequencer-master.scala 643:40]
  wire  _GEN_7968 = io_op_bits_active_vidiv ? _GEN_6280 : _GEN_5550; // @[sequencer-master.scala 643:40]
  wire  _GEN_7969 = io_op_bits_active_vidiv ? _GEN_6281 : _GEN_5551; // @[sequencer-master.scala 643:40]
  wire  _GEN_7970 = io_op_bits_active_vidiv ? _GEN_6282 : _GEN_5552; // @[sequencer-master.scala 643:40]
  wire  _GEN_7971 = io_op_bits_active_vidiv ? _GEN_6283 : _GEN_5553; // @[sequencer-master.scala 643:40]
  wire  _GEN_7972 = io_op_bits_active_vidiv ? _GEN_6284 : _GEN_5554; // @[sequencer-master.scala 643:40]
  wire  _GEN_7973 = io_op_bits_active_vidiv ? _GEN_6285 : _GEN_5555; // @[sequencer-master.scala 643:40]
  wire  _GEN_7974 = io_op_bits_active_vidiv ? _GEN_6286 : _GEN_5556; // @[sequencer-master.scala 643:40]
  wire  _GEN_7975 = io_op_bits_active_vidiv ? _GEN_6287 : _GEN_5557; // @[sequencer-master.scala 643:40]
  wire  _GEN_7976 = io_op_bits_active_vidiv ? _GEN_6288 : _GEN_5558; // @[sequencer-master.scala 643:40]
  wire  _GEN_7977 = io_op_bits_active_vidiv ? _GEN_6289 : _GEN_5559; // @[sequencer-master.scala 643:40]
  wire  _GEN_7978 = io_op_bits_active_vidiv ? _GEN_6290 : _GEN_5560; // @[sequencer-master.scala 643:40]
  wire  _GEN_7979 = io_op_bits_active_vidiv ? _GEN_6291 : _GEN_5561; // @[sequencer-master.scala 643:40]
  wire  _GEN_7980 = io_op_bits_active_vidiv ? _GEN_6292 : _GEN_5562; // @[sequencer-master.scala 643:40]
  wire  _GEN_7981 = io_op_bits_active_vidiv ? _GEN_6293 : _GEN_5563; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7982 = io_op_bits_active_vidiv ? _GEN_6294 : _GEN_5564; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7983 = io_op_bits_active_vidiv ? _GEN_6295 : _GEN_5565; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7984 = io_op_bits_active_vidiv ? _GEN_6296 : _GEN_5566; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7985 = io_op_bits_active_vidiv ? _GEN_6297 : _GEN_5567; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7986 = io_op_bits_active_vidiv ? _GEN_6298 : _GEN_5568; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7987 = io_op_bits_active_vidiv ? _GEN_6299 : _GEN_5569; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7988 = io_op_bits_active_vidiv ? _GEN_6300 : _GEN_5570; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_7989 = io_op_bits_active_vidiv ? _GEN_6301 : _GEN_5571; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7990 = io_op_bits_active_vidiv ? _GEN_6302 : _GEN_5572; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7991 = io_op_bits_active_vidiv ? _GEN_6303 : _GEN_5573; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7992 = io_op_bits_active_vidiv ? _GEN_6304 : _GEN_5574; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7993 = io_op_bits_active_vidiv ? _GEN_6305 : _GEN_5575; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7994 = io_op_bits_active_vidiv ? _GEN_6306 : _GEN_5576; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7995 = io_op_bits_active_vidiv ? _GEN_6307 : _GEN_5577; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7996 = io_op_bits_active_vidiv ? _GEN_6308 : _GEN_5578; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_7997 = io_op_bits_active_vidiv ? _GEN_6309 : _GEN_5579; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_7998 = io_op_bits_active_vidiv ? _GEN_6310 : _GEN_5580; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_7999 = io_op_bits_active_vidiv ? _GEN_6311 : _GEN_5581; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8000 = io_op_bits_active_vidiv ? _GEN_6312 : _GEN_5582; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8001 = io_op_bits_active_vidiv ? _GEN_6313 : _GEN_5583; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8002 = io_op_bits_active_vidiv ? _GEN_6314 : _GEN_5584; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8003 = io_op_bits_active_vidiv ? _GEN_6315 : _GEN_5585; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8004 = io_op_bits_active_vidiv ? _GEN_6316 : _GEN_5586; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8005 = io_op_bits_active_vidiv ? _GEN_6317 : _GEN_5587; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8006 = io_op_bits_active_vidiv ? _GEN_6510 : _GEN_5588; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8007 = io_op_bits_active_vidiv ? _GEN_6511 : _GEN_5589; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8008 = io_op_bits_active_vidiv ? _GEN_6512 : _GEN_5590; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8009 = io_op_bits_active_vidiv ? _GEN_6513 : _GEN_5591; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8010 = io_op_bits_active_vidiv ? _GEN_6514 : _GEN_5592; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8011 = io_op_bits_active_vidiv ? _GEN_6515 : _GEN_5593; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8012 = io_op_bits_active_vidiv ? _GEN_6516 : _GEN_5594; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8013 = io_op_bits_active_vidiv ? _GEN_6517 : _GEN_5595; // @[sequencer-master.scala 643:40]
  wire  _GEN_8014 = io_op_bits_active_vidiv ? _GEN_6526 : _GEN_5596; // @[sequencer-master.scala 643:40]
  wire  _GEN_8015 = io_op_bits_active_vidiv ? _GEN_6527 : _GEN_5597; // @[sequencer-master.scala 643:40]
  wire  _GEN_8016 = io_op_bits_active_vidiv ? _GEN_6528 : _GEN_5598; // @[sequencer-master.scala 643:40]
  wire  _GEN_8017 = io_op_bits_active_vidiv ? _GEN_6529 : _GEN_5599; // @[sequencer-master.scala 643:40]
  wire  _GEN_8018 = io_op_bits_active_vidiv ? _GEN_6530 : _GEN_5600; // @[sequencer-master.scala 643:40]
  wire  _GEN_8019 = io_op_bits_active_vidiv ? _GEN_6531 : _GEN_5601; // @[sequencer-master.scala 643:40]
  wire  _GEN_8020 = io_op_bits_active_vidiv ? _GEN_6532 : _GEN_5602; // @[sequencer-master.scala 643:40]
  wire  _GEN_8021 = io_op_bits_active_vidiv ? _GEN_6533 : _GEN_5603; // @[sequencer-master.scala 643:40]
  wire  _GEN_8022 = io_op_bits_active_vidiv ? _GEN_6534 : _GEN_5604; // @[sequencer-master.scala 643:40]
  wire  _GEN_8023 = io_op_bits_active_vidiv ? _GEN_6535 : _GEN_5605; // @[sequencer-master.scala 643:40]
  wire  _GEN_8024 = io_op_bits_active_vidiv ? _GEN_6536 : _GEN_5606; // @[sequencer-master.scala 643:40]
  wire  _GEN_8025 = io_op_bits_active_vidiv ? _GEN_6537 : _GEN_5607; // @[sequencer-master.scala 643:40]
  wire  _GEN_8026 = io_op_bits_active_vidiv ? _GEN_6538 : _GEN_5608; // @[sequencer-master.scala 643:40]
  wire  _GEN_8027 = io_op_bits_active_vidiv ? _GEN_6539 : _GEN_5609; // @[sequencer-master.scala 643:40]
  wire  _GEN_8028 = io_op_bits_active_vidiv ? _GEN_6540 : _GEN_5610; // @[sequencer-master.scala 643:40]
  wire  _GEN_8029 = io_op_bits_active_vidiv ? _GEN_6541 : _GEN_5611; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8030 = io_op_bits_active_vidiv ? _GEN_6542 : _GEN_5612; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8031 = io_op_bits_active_vidiv ? _GEN_6543 : _GEN_5613; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8032 = io_op_bits_active_vidiv ? _GEN_6544 : _GEN_5614; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8033 = io_op_bits_active_vidiv ? _GEN_6545 : _GEN_5615; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8034 = io_op_bits_active_vidiv ? _GEN_6546 : _GEN_5616; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8035 = io_op_bits_active_vidiv ? _GEN_6547 : _GEN_5617; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8036 = io_op_bits_active_vidiv ? _GEN_6548 : _GEN_5618; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8037 = io_op_bits_active_vidiv ? _GEN_6549 : _GEN_5619; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8038 = io_op_bits_active_vidiv ? _GEN_6550 : _GEN_5620; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8039 = io_op_bits_active_vidiv ? _GEN_6551 : _GEN_5621; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8040 = io_op_bits_active_vidiv ? _GEN_6552 : _GEN_5622; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8041 = io_op_bits_active_vidiv ? _GEN_6553 : _GEN_5623; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8042 = io_op_bits_active_vidiv ? _GEN_6554 : _GEN_5624; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8043 = io_op_bits_active_vidiv ? _GEN_6555 : _GEN_5625; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8044 = io_op_bits_active_vidiv ? _GEN_6556 : _GEN_5626; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8045 = io_op_bits_active_vidiv ? _GEN_6557 : _GEN_5627; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8046 = io_op_bits_active_vidiv ? _GEN_6558 : _GEN_5628; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8047 = io_op_bits_active_vidiv ? _GEN_6559 : _GEN_5629; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8048 = io_op_bits_active_vidiv ? _GEN_6560 : _GEN_5630; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8049 = io_op_bits_active_vidiv ? _GEN_6561 : _GEN_5631; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8050 = io_op_bits_active_vidiv ? _GEN_6562 : _GEN_5632; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8051 = io_op_bits_active_vidiv ? _GEN_6563 : _GEN_5633; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8052 = io_op_bits_active_vidiv ? _GEN_6564 : _GEN_5634; // @[sequencer-master.scala 643:40]
  wire [63:0] _GEN_8053 = io_op_bits_active_vidiv ? _GEN_6565 : _GEN_5635; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8054 = io_op_bits_active_vidiv ? _GEN_7614 : _GEN_5676; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8055 = io_op_bits_active_vidiv ? _GEN_7615 : _GEN_5677; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8056 = io_op_bits_active_vidiv ? _GEN_7616 : _GEN_5678; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8057 = io_op_bits_active_vidiv ? _GEN_7617 : _GEN_5679; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8058 = io_op_bits_active_vidiv ? _GEN_7618 : _GEN_5680; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8059 = io_op_bits_active_vidiv ? _GEN_7619 : _GEN_5681; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8060 = io_op_bits_active_vidiv ? _GEN_7620 : _GEN_5682; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8061 = io_op_bits_active_vidiv ? _GEN_7621 : _GEN_5683; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8062 = io_op_bits_active_vidiv ? _GEN_7622 : _GEN_5684; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8063 = io_op_bits_active_vidiv ? _GEN_7623 : _GEN_5685; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8064 = io_op_bits_active_vidiv ? _GEN_7624 : _GEN_5686; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8065 = io_op_bits_active_vidiv ? _GEN_7625 : _GEN_5687; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8066 = io_op_bits_active_vidiv ? _GEN_7626 : _GEN_5688; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8067 = io_op_bits_active_vidiv ? _GEN_7627 : _GEN_5689; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8068 = io_op_bits_active_vidiv ? _GEN_7628 : _GEN_5690; // @[sequencer-master.scala 643:40]
  wire [3:0] _GEN_8069 = io_op_bits_active_vidiv ? _GEN_7629 : _GEN_5691; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8070 = io_op_bits_active_vidiv ? _GEN_7630 : _GEN_5692; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8071 = io_op_bits_active_vidiv ? _GEN_7631 : _GEN_5693; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8072 = io_op_bits_active_vidiv ? _GEN_7632 : _GEN_5694; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8073 = io_op_bits_active_vidiv ? _GEN_7633 : _GEN_5695; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8074 = io_op_bits_active_vidiv ? _GEN_7634 : _GEN_5696; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8075 = io_op_bits_active_vidiv ? _GEN_7635 : _GEN_5697; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8076 = io_op_bits_active_vidiv ? _GEN_7636 : _GEN_5698; // @[sequencer-master.scala 643:40]
  wire [2:0] _GEN_8077 = io_op_bits_active_vidiv ? _GEN_7637 : _GEN_5699; // @[sequencer-master.scala 643:40]
  wire  _GEN_8078 = io_op_bits_active_vidiv ? _GEN_7246 : e_0_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8079 = io_op_bits_active_vidiv ? _GEN_7247 : e_1_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8080 = io_op_bits_active_vidiv ? _GEN_7248 : e_2_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8081 = io_op_bits_active_vidiv ? _GEN_7249 : e_3_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8082 = io_op_bits_active_vidiv ? _GEN_7250 : e_4_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8083 = io_op_bits_active_vidiv ? _GEN_7251 : e_5_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8084 = io_op_bits_active_vidiv ? _GEN_7252 : e_6_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire  _GEN_8085 = io_op_bits_active_vidiv ? _GEN_7253 : e_7_active_vidu; // @[sequencer-master.scala 643:40 sequencer-master.scala 109:14]
  wire [7:0] _GEN_8086 = io_op_bits_active_vidiv ? _GEN_7310 : _GEN_5636; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8087 = io_op_bits_active_vidiv ? _GEN_7311 : _GEN_5637; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8088 = io_op_bits_active_vidiv ? _GEN_7312 : _GEN_5638; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8089 = io_op_bits_active_vidiv ? _GEN_7313 : _GEN_5639; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8090 = io_op_bits_active_vidiv ? _GEN_7314 : _GEN_5640; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8091 = io_op_bits_active_vidiv ? _GEN_7315 : _GEN_5641; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8092 = io_op_bits_active_vidiv ? _GEN_7316 : _GEN_5642; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8093 = io_op_bits_active_vidiv ? _GEN_7317 : _GEN_5643; // @[sequencer-master.scala 643:40]
  wire  _GEN_8094 = io_op_bits_active_vidiv ? _GEN_7326 : _GEN_5644; // @[sequencer-master.scala 643:40]
  wire  _GEN_8095 = io_op_bits_active_vidiv ? _GEN_7327 : _GEN_5645; // @[sequencer-master.scala 643:40]
  wire  _GEN_8096 = io_op_bits_active_vidiv ? _GEN_7328 : _GEN_5646; // @[sequencer-master.scala 643:40]
  wire  _GEN_8097 = io_op_bits_active_vidiv ? _GEN_7329 : _GEN_5647; // @[sequencer-master.scala 643:40]
  wire  _GEN_8098 = io_op_bits_active_vidiv ? _GEN_7330 : _GEN_5648; // @[sequencer-master.scala 643:40]
  wire  _GEN_8099 = io_op_bits_active_vidiv ? _GEN_7331 : _GEN_5649; // @[sequencer-master.scala 643:40]
  wire  _GEN_8100 = io_op_bits_active_vidiv ? _GEN_7332 : _GEN_5650; // @[sequencer-master.scala 643:40]
  wire  _GEN_8101 = io_op_bits_active_vidiv ? _GEN_7333 : _GEN_5651; // @[sequencer-master.scala 643:40]
  wire  _GEN_8102 = io_op_bits_active_vidiv ? _GEN_7334 : _GEN_5652; // @[sequencer-master.scala 643:40]
  wire  _GEN_8103 = io_op_bits_active_vidiv ? _GEN_7335 : _GEN_5653; // @[sequencer-master.scala 643:40]
  wire  _GEN_8104 = io_op_bits_active_vidiv ? _GEN_7336 : _GEN_5654; // @[sequencer-master.scala 643:40]
  wire  _GEN_8105 = io_op_bits_active_vidiv ? _GEN_7337 : _GEN_5655; // @[sequencer-master.scala 643:40]
  wire  _GEN_8106 = io_op_bits_active_vidiv ? _GEN_7338 : _GEN_5656; // @[sequencer-master.scala 643:40]
  wire  _GEN_8107 = io_op_bits_active_vidiv ? _GEN_7339 : _GEN_5657; // @[sequencer-master.scala 643:40]
  wire  _GEN_8108 = io_op_bits_active_vidiv ? _GEN_7340 : _GEN_5658; // @[sequencer-master.scala 643:40]
  wire  _GEN_8109 = io_op_bits_active_vidiv ? _GEN_7341 : _GEN_5659; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8110 = io_op_bits_active_vidiv ? _GEN_7342 : _GEN_5660; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8111 = io_op_bits_active_vidiv ? _GEN_7343 : _GEN_5661; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8112 = io_op_bits_active_vidiv ? _GEN_7344 : _GEN_5662; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8113 = io_op_bits_active_vidiv ? _GEN_7345 : _GEN_5663; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8114 = io_op_bits_active_vidiv ? _GEN_7346 : _GEN_5664; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8115 = io_op_bits_active_vidiv ? _GEN_7347 : _GEN_5665; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8116 = io_op_bits_active_vidiv ? _GEN_7348 : _GEN_5666; // @[sequencer-master.scala 643:40]
  wire [1:0] _GEN_8117 = io_op_bits_active_vidiv ? _GEN_7349 : _GEN_5667; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8118 = io_op_bits_active_vidiv ? _GEN_7350 : _GEN_5668; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8119 = io_op_bits_active_vidiv ? _GEN_7351 : _GEN_5669; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8120 = io_op_bits_active_vidiv ? _GEN_7352 : _GEN_5670; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8121 = io_op_bits_active_vidiv ? _GEN_7353 : _GEN_5671; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8122 = io_op_bits_active_vidiv ? _GEN_7354 : _GEN_5672; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8123 = io_op_bits_active_vidiv ? _GEN_7355 : _GEN_5673; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8124 = io_op_bits_active_vidiv ? _GEN_7356 : _GEN_5674; // @[sequencer-master.scala 643:40]
  wire [7:0] _GEN_8125 = io_op_bits_active_vidiv ? _GEN_7357 : _GEN_5675; // @[sequencer-master.scala 643:40]
  wire  _GEN_8126 = io_op_bits_active_vidiv | _GEN_5700; // @[sequencer-master.scala 643:40 sequencer-master.scala 265:41]
  wire [2:0] _GEN_8127 = io_op_bits_active_vidiv ? _T_1647 : _GEN_5701; // @[sequencer-master.scala 643:40 sequencer-master.scala 265:66]
  wire  _T_1966 = io_op_bits_fn_union[7:6] == 2'h1; // @[types-vxu.scala 53:51]
  wire  _T_1967 = io_op_bits_fn_union[7:6] == 2'h0; // @[types-vxu.scala 53:51]
  wire  _T_1968 = io_op_bits_fn_union[7:6] == 2'h2; // @[types-vxu.scala 53:51]
  wire  _GEN_8128 = _GEN_32729 | _GEN_7638; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8129 = _GEN_32730 | _GEN_7639; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8130 = _GEN_32731 | _GEN_7640; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8131 = _GEN_32732 | _GEN_7641; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8132 = _GEN_32733 | _GEN_7642; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8133 = _GEN_32734 | _GEN_7643; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8134 = _GEN_32735 | _GEN_7644; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8135 = _GEN_32736 | _GEN_7645; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_8144 = 3'h0 == tail ? 1'h0 : _GEN_7654; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8145 = 3'h1 == tail ? 1'h0 : _GEN_7655; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8146 = 3'h2 == tail ? 1'h0 : _GEN_7656; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8147 = 3'h3 == tail ? 1'h0 : _GEN_7657; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8148 = 3'h4 == tail ? 1'h0 : _GEN_7658; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8149 = 3'h5 == tail ? 1'h0 : _GEN_7659; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8150 = 3'h6 == tail ? 1'h0 : _GEN_7660; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8151 = 3'h7 == tail ? 1'h0 : _GEN_7661; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_8152 = 3'h0 == tail ? 1'h0 : _GEN_7662; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8153 = 3'h1 == tail ? 1'h0 : _GEN_7663; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8154 = 3'h2 == tail ? 1'h0 : _GEN_7664; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8155 = 3'h3 == tail ? 1'h0 : _GEN_7665; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8156 = 3'h4 == tail ? 1'h0 : _GEN_7666; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8157 = 3'h5 == tail ? 1'h0 : _GEN_7667; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8158 = 3'h6 == tail ? 1'h0 : _GEN_7668; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8159 = 3'h7 == tail ? 1'h0 : _GEN_7669; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_8160 = 3'h0 == tail ? 1'h0 : _GEN_7670; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8161 = 3'h1 == tail ? 1'h0 : _GEN_7671; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8162 = 3'h2 == tail ? 1'h0 : _GEN_7672; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8163 = 3'h3 == tail ? 1'h0 : _GEN_7673; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8164 = 3'h4 == tail ? 1'h0 : _GEN_7674; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8165 = 3'h5 == tail ? 1'h0 : _GEN_7675; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8166 = 3'h6 == tail ? 1'h0 : _GEN_7676; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8167 = 3'h7 == tail ? 1'h0 : _GEN_7677; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_8168 = 3'h0 == tail ? 1'h0 : _GEN_7678; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8169 = 3'h1 == tail ? 1'h0 : _GEN_7679; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8170 = 3'h2 == tail ? 1'h0 : _GEN_7680; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8171 = 3'h3 == tail ? 1'h0 : _GEN_7681; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8172 = 3'h4 == tail ? 1'h0 : _GEN_7682; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8173 = 3'h5 == tail ? 1'h0 : _GEN_7683; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8174 = 3'h6 == tail ? 1'h0 : _GEN_7684; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8175 = 3'h7 == tail ? 1'h0 : _GEN_7685; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_8176 = 3'h0 == tail ? 1'h0 : _GEN_7686; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8177 = 3'h1 == tail ? 1'h0 : _GEN_7687; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8178 = 3'h2 == tail ? 1'h0 : _GEN_7688; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8179 = 3'h3 == tail ? 1'h0 : _GEN_7689; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8180 = 3'h4 == tail ? 1'h0 : _GEN_7690; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8181 = 3'h5 == tail ? 1'h0 : _GEN_7691; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8182 = 3'h6 == tail ? 1'h0 : _GEN_7692; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8183 = 3'h7 == tail ? 1'h0 : _GEN_7693; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_8184 = _GEN_32729 | _GEN_7694; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8185 = _GEN_32730 | _GEN_7695; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8186 = _GEN_32731 | _GEN_7696; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8187 = _GEN_32732 | _GEN_7697; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8188 = _GEN_32733 | _GEN_7698; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8189 = _GEN_32734 | _GEN_7699; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8190 = _GEN_32735 | _GEN_7700; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8191 = _GEN_32736 | _GEN_7701; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_8192 = 3'h0 == tail ? 1'h0 : _GEN_7702; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8193 = 3'h1 == tail ? 1'h0 : _GEN_7703; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8194 = 3'h2 == tail ? 1'h0 : _GEN_7704; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8195 = 3'h3 == tail ? 1'h0 : _GEN_7705; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8196 = 3'h4 == tail ? 1'h0 : _GEN_7706; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8197 = 3'h5 == tail ? 1'h0 : _GEN_7707; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8198 = 3'h6 == tail ? 1'h0 : _GEN_7708; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8199 = 3'h7 == tail ? 1'h0 : _GEN_7709; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8200 = 3'h0 == tail ? 1'h0 : _GEN_7710; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8201 = 3'h1 == tail ? 1'h0 : _GEN_7711; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8202 = 3'h2 == tail ? 1'h0 : _GEN_7712; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8203 = 3'h3 == tail ? 1'h0 : _GEN_7713; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8204 = 3'h4 == tail ? 1'h0 : _GEN_7714; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8205 = 3'h5 == tail ? 1'h0 : _GEN_7715; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8206 = 3'h6 == tail ? 1'h0 : _GEN_7716; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8207 = 3'h7 == tail ? 1'h0 : _GEN_7717; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8208 = 3'h0 == tail ? 1'h0 : _GEN_7718; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8209 = 3'h1 == tail ? 1'h0 : _GEN_7719; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8210 = 3'h2 == tail ? 1'h0 : _GEN_7720; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8211 = 3'h3 == tail ? 1'h0 : _GEN_7721; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8212 = 3'h4 == tail ? 1'h0 : _GEN_7722; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8213 = 3'h5 == tail ? 1'h0 : _GEN_7723; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8214 = 3'h6 == tail ? 1'h0 : _GEN_7724; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8215 = 3'h7 == tail ? 1'h0 : _GEN_7725; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8216 = 3'h0 == tail ? 1'h0 : _GEN_7726; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8217 = 3'h1 == tail ? 1'h0 : _GEN_7727; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8218 = 3'h2 == tail ? 1'h0 : _GEN_7728; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8219 = 3'h3 == tail ? 1'h0 : _GEN_7729; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8220 = 3'h4 == tail ? 1'h0 : _GEN_7730; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8221 = 3'h5 == tail ? 1'h0 : _GEN_7731; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8222 = 3'h6 == tail ? 1'h0 : _GEN_7732; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8223 = 3'h7 == tail ? 1'h0 : _GEN_7733; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8224 = 3'h0 == tail ? 1'h0 : _GEN_7734; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8225 = 3'h1 == tail ? 1'h0 : _GEN_7735; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8226 = 3'h2 == tail ? 1'h0 : _GEN_7736; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8227 = 3'h3 == tail ? 1'h0 : _GEN_7737; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8228 = 3'h4 == tail ? 1'h0 : _GEN_7738; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8229 = 3'h5 == tail ? 1'h0 : _GEN_7739; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8230 = 3'h6 == tail ? 1'h0 : _GEN_7740; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8231 = 3'h7 == tail ? 1'h0 : _GEN_7741; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8232 = 3'h0 == tail ? 1'h0 : _GEN_7742; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8233 = 3'h1 == tail ? 1'h0 : _GEN_7743; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8234 = 3'h2 == tail ? 1'h0 : _GEN_7744; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8235 = 3'h3 == tail ? 1'h0 : _GEN_7745; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8236 = 3'h4 == tail ? 1'h0 : _GEN_7746; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8237 = 3'h5 == tail ? 1'h0 : _GEN_7747; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8238 = 3'h6 == tail ? 1'h0 : _GEN_7748; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8239 = 3'h7 == tail ? 1'h0 : _GEN_7749; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8240 = 3'h0 == tail ? 1'h0 : _GEN_7750; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8241 = 3'h1 == tail ? 1'h0 : _GEN_7751; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8242 = 3'h2 == tail ? 1'h0 : _GEN_7752; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8243 = 3'h3 == tail ? 1'h0 : _GEN_7753; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8244 = 3'h4 == tail ? 1'h0 : _GEN_7754; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8245 = 3'h5 == tail ? 1'h0 : _GEN_7755; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8246 = 3'h6 == tail ? 1'h0 : _GEN_7756; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8247 = 3'h7 == tail ? 1'h0 : _GEN_7757; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8248 = 3'h0 == tail ? 1'h0 : _GEN_7758; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8249 = 3'h1 == tail ? 1'h0 : _GEN_7759; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8250 = 3'h2 == tail ? 1'h0 : _GEN_7760; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8251 = 3'h3 == tail ? 1'h0 : _GEN_7761; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8252 = 3'h4 == tail ? 1'h0 : _GEN_7762; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8253 = 3'h5 == tail ? 1'h0 : _GEN_7763; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8254 = 3'h6 == tail ? 1'h0 : _GEN_7764; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8255 = 3'h7 == tail ? 1'h0 : _GEN_7765; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8256 = 3'h0 == tail ? 1'h0 : _GEN_7766; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8257 = 3'h1 == tail ? 1'h0 : _GEN_7767; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8258 = 3'h2 == tail ? 1'h0 : _GEN_7768; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8259 = 3'h3 == tail ? 1'h0 : _GEN_7769; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8260 = 3'h4 == tail ? 1'h0 : _GEN_7770; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8261 = 3'h5 == tail ? 1'h0 : _GEN_7771; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8262 = 3'h6 == tail ? 1'h0 : _GEN_7772; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8263 = 3'h7 == tail ? 1'h0 : _GEN_7773; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8264 = 3'h0 == tail ? 1'h0 : _GEN_7774; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8265 = 3'h1 == tail ? 1'h0 : _GEN_7775; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8266 = 3'h2 == tail ? 1'h0 : _GEN_7776; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8267 = 3'h3 == tail ? 1'h0 : _GEN_7777; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8268 = 3'h4 == tail ? 1'h0 : _GEN_7778; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8269 = 3'h5 == tail ? 1'h0 : _GEN_7779; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8270 = 3'h6 == tail ? 1'h0 : _GEN_7780; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8271 = 3'h7 == tail ? 1'h0 : _GEN_7781; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8272 = 3'h0 == tail ? 1'h0 : _GEN_7782; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8273 = 3'h1 == tail ? 1'h0 : _GEN_7783; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8274 = 3'h2 == tail ? 1'h0 : _GEN_7784; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8275 = 3'h3 == tail ? 1'h0 : _GEN_7785; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8276 = 3'h4 == tail ? 1'h0 : _GEN_7786; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8277 = 3'h5 == tail ? 1'h0 : _GEN_7787; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8278 = 3'h6 == tail ? 1'h0 : _GEN_7788; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8279 = 3'h7 == tail ? 1'h0 : _GEN_7789; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8280 = 3'h0 == tail ? 1'h0 : _GEN_7790; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8281 = 3'h1 == tail ? 1'h0 : _GEN_7791; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8282 = 3'h2 == tail ? 1'h0 : _GEN_7792; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8283 = 3'h3 == tail ? 1'h0 : _GEN_7793; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8284 = 3'h4 == tail ? 1'h0 : _GEN_7794; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8285 = 3'h5 == tail ? 1'h0 : _GEN_7795; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8286 = 3'h6 == tail ? 1'h0 : _GEN_7796; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8287 = 3'h7 == tail ? 1'h0 : _GEN_7797; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8288 = 3'h0 == tail ? 1'h0 : _GEN_7798; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8289 = 3'h1 == tail ? 1'h0 : _GEN_7799; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8290 = 3'h2 == tail ? 1'h0 : _GEN_7800; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8291 = 3'h3 == tail ? 1'h0 : _GEN_7801; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8292 = 3'h4 == tail ? 1'h0 : _GEN_7802; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8293 = 3'h5 == tail ? 1'h0 : _GEN_7803; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8294 = 3'h6 == tail ? 1'h0 : _GEN_7804; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8295 = 3'h7 == tail ? 1'h0 : _GEN_7805; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8296 = 3'h0 == tail ? 1'h0 : _GEN_7806; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8297 = 3'h1 == tail ? 1'h0 : _GEN_7807; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8298 = 3'h2 == tail ? 1'h0 : _GEN_7808; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8299 = 3'h3 == tail ? 1'h0 : _GEN_7809; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8300 = 3'h4 == tail ? 1'h0 : _GEN_7810; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8301 = 3'h5 == tail ? 1'h0 : _GEN_7811; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8302 = 3'h6 == tail ? 1'h0 : _GEN_7812; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8303 = 3'h7 == tail ? 1'h0 : _GEN_7813; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8304 = 3'h0 == tail ? 1'h0 : _GEN_7814; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8305 = 3'h1 == tail ? 1'h0 : _GEN_7815; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8306 = 3'h2 == tail ? 1'h0 : _GEN_7816; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8307 = 3'h3 == tail ? 1'h0 : _GEN_7817; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8308 = 3'h4 == tail ? 1'h0 : _GEN_7818; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8309 = 3'h5 == tail ? 1'h0 : _GEN_7819; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8310 = 3'h6 == tail ? 1'h0 : _GEN_7820; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8311 = 3'h7 == tail ? 1'h0 : _GEN_7821; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8312 = 3'h0 == tail ? 1'h0 : _GEN_7822; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8313 = 3'h1 == tail ? 1'h0 : _GEN_7823; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8314 = 3'h2 == tail ? 1'h0 : _GEN_7824; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8315 = 3'h3 == tail ? 1'h0 : _GEN_7825; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8316 = 3'h4 == tail ? 1'h0 : _GEN_7826; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8317 = 3'h5 == tail ? 1'h0 : _GEN_7827; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8318 = 3'h6 == tail ? 1'h0 : _GEN_7828; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8319 = 3'h7 == tail ? 1'h0 : _GEN_7829; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8320 = 3'h0 == tail ? 1'h0 : _GEN_7830; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8321 = 3'h1 == tail ? 1'h0 : _GEN_7831; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8322 = 3'h2 == tail ? 1'h0 : _GEN_7832; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8323 = 3'h3 == tail ? 1'h0 : _GEN_7833; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8324 = 3'h4 == tail ? 1'h0 : _GEN_7834; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8325 = 3'h5 == tail ? 1'h0 : _GEN_7835; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8326 = 3'h6 == tail ? 1'h0 : _GEN_7836; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8327 = 3'h7 == tail ? 1'h0 : _GEN_7837; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8328 = 3'h0 == tail ? 1'h0 : _GEN_7838; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8329 = 3'h1 == tail ? 1'h0 : _GEN_7839; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8330 = 3'h2 == tail ? 1'h0 : _GEN_7840; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8331 = 3'h3 == tail ? 1'h0 : _GEN_7841; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8332 = 3'h4 == tail ? 1'h0 : _GEN_7842; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8333 = 3'h5 == tail ? 1'h0 : _GEN_7843; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8334 = 3'h6 == tail ? 1'h0 : _GEN_7844; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8335 = 3'h7 == tail ? 1'h0 : _GEN_7845; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8336 = 3'h0 == tail ? 1'h0 : _GEN_7846; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8337 = 3'h1 == tail ? 1'h0 : _GEN_7847; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8338 = 3'h2 == tail ? 1'h0 : _GEN_7848; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8339 = 3'h3 == tail ? 1'h0 : _GEN_7849; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8340 = 3'h4 == tail ? 1'h0 : _GEN_7850; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8341 = 3'h5 == tail ? 1'h0 : _GEN_7851; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8342 = 3'h6 == tail ? 1'h0 : _GEN_7852; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8343 = 3'h7 == tail ? 1'h0 : _GEN_7853; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8344 = 3'h0 == tail ? 1'h0 : _GEN_7854; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8345 = 3'h1 == tail ? 1'h0 : _GEN_7855; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8346 = 3'h2 == tail ? 1'h0 : _GEN_7856; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8347 = 3'h3 == tail ? 1'h0 : _GEN_7857; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8348 = 3'h4 == tail ? 1'h0 : _GEN_7858; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8349 = 3'h5 == tail ? 1'h0 : _GEN_7859; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8350 = 3'h6 == tail ? 1'h0 : _GEN_7860; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8351 = 3'h7 == tail ? 1'h0 : _GEN_7861; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8352 = 3'h0 == tail ? 1'h0 : _GEN_7862; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8353 = 3'h1 == tail ? 1'h0 : _GEN_7863; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8354 = 3'h2 == tail ? 1'h0 : _GEN_7864; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8355 = 3'h3 == tail ? 1'h0 : _GEN_7865; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8356 = 3'h4 == tail ? 1'h0 : _GEN_7866; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8357 = 3'h5 == tail ? 1'h0 : _GEN_7867; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8358 = 3'h6 == tail ? 1'h0 : _GEN_7868; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8359 = 3'h7 == tail ? 1'h0 : _GEN_7869; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8360 = 3'h0 == tail ? 1'h0 : _GEN_7870; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8361 = 3'h1 == tail ? 1'h0 : _GEN_7871; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8362 = 3'h2 == tail ? 1'h0 : _GEN_7872; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8363 = 3'h3 == tail ? 1'h0 : _GEN_7873; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8364 = 3'h4 == tail ? 1'h0 : _GEN_7874; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8365 = 3'h5 == tail ? 1'h0 : _GEN_7875; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8366 = 3'h6 == tail ? 1'h0 : _GEN_7876; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8367 = 3'h7 == tail ? 1'h0 : _GEN_7877; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_8368 = 3'h0 == tail ? 1'h0 : _GEN_7878; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8369 = 3'h1 == tail ? 1'h0 : _GEN_7879; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8370 = 3'h2 == tail ? 1'h0 : _GEN_7880; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8371 = 3'h3 == tail ? 1'h0 : _GEN_7881; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8372 = 3'h4 == tail ? 1'h0 : _GEN_7882; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8373 = 3'h5 == tail ? 1'h0 : _GEN_7883; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8374 = 3'h6 == tail ? 1'h0 : _GEN_7884; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8375 = 3'h7 == tail ? 1'h0 : _GEN_7885; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_8376 = 3'h0 == tail ? 1'h0 : _GEN_7886; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8377 = 3'h1 == tail ? 1'h0 : _GEN_7887; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8378 = 3'h2 == tail ? 1'h0 : _GEN_7888; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8379 = 3'h3 == tail ? 1'h0 : _GEN_7889; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8380 = 3'h4 == tail ? 1'h0 : _GEN_7890; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8381 = 3'h5 == tail ? 1'h0 : _GEN_7891; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8382 = 3'h6 == tail ? 1'h0 : _GEN_7892; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8383 = 3'h7 == tail ? 1'h0 : _GEN_7893; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_8384 = 3'h0 == tail ? 1'h0 : _GEN_7894; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8385 = 3'h1 == tail ? 1'h0 : _GEN_7895; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8386 = 3'h2 == tail ? 1'h0 : _GEN_7896; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8387 = 3'h3 == tail ? 1'h0 : _GEN_7897; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8388 = 3'h4 == tail ? 1'h0 : _GEN_7898; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8389 = 3'h5 == tail ? 1'h0 : _GEN_7899; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8390 = 3'h6 == tail ? 1'h0 : _GEN_7900; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8391 = 3'h7 == tail ? 1'h0 : _GEN_7901; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_8400 = _GEN_32729 | e_0_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8401 = _GEN_32730 | e_1_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8402 = _GEN_32731 | e_2_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8403 = _GEN_32732 | e_3_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8404 = _GEN_32733 | e_4_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8405 = _GEN_32734 | e_5_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8406 = _GEN_32735 | e_6_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_8407 = _GEN_32736 | e_7_active_vfmu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_8408 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_7918; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8409 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_7919; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8410 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_7920; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8411 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_7921; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8412 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_7922; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8413 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_7923; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8414 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_7924; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_8415 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_7925; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_8416 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_7926; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8417 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_7927; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8418 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_7928; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8419 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_7929; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8420 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_7930; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8421 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_7931; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8422 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_7932; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_8423 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_7933; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8424 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_8144; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8425 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_8145; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8426 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_8146; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8427 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_8147; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8428 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_8148; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8429 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_8149; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8430 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_8150; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8431 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_8151; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8432 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_7934; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8433 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_7935; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8434 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_7936; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8435 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_7937; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8436 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_7938; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8437 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_7939; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8438 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_7940; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8439 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_7941; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8440 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_7942; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8441 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_7943; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8442 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_7944; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8443 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_7945; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8444 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_7946; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8445 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_7947; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8446 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_7948; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_8447 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_7949; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_8448 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_7950; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8449 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_7951; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8450 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_7952; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8451 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_7953; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8452 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_7954; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8453 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_7955; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8454 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_7956; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_8455 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_7957; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_8456 = io_op_bits_base_vp_valid ? _GEN_8416 : _GEN_7926; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8457 = io_op_bits_base_vp_valid ? _GEN_8417 : _GEN_7927; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8458 = io_op_bits_base_vp_valid ? _GEN_8418 : _GEN_7928; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8459 = io_op_bits_base_vp_valid ? _GEN_8419 : _GEN_7929; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8460 = io_op_bits_base_vp_valid ? _GEN_8420 : _GEN_7930; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8461 = io_op_bits_base_vp_valid ? _GEN_8421 : _GEN_7931; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8462 = io_op_bits_base_vp_valid ? _GEN_8422 : _GEN_7932; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_8463 = io_op_bits_base_vp_valid ? _GEN_8423 : _GEN_7933; // @[sequencer-master.scala 320:41]
  wire  _GEN_8464 = io_op_bits_base_vp_valid ? _GEN_8424 : _GEN_8144; // @[sequencer-master.scala 320:41]
  wire  _GEN_8465 = io_op_bits_base_vp_valid ? _GEN_8425 : _GEN_8145; // @[sequencer-master.scala 320:41]
  wire  _GEN_8466 = io_op_bits_base_vp_valid ? _GEN_8426 : _GEN_8146; // @[sequencer-master.scala 320:41]
  wire  _GEN_8467 = io_op_bits_base_vp_valid ? _GEN_8427 : _GEN_8147; // @[sequencer-master.scala 320:41]
  wire  _GEN_8468 = io_op_bits_base_vp_valid ? _GEN_8428 : _GEN_8148; // @[sequencer-master.scala 320:41]
  wire  _GEN_8469 = io_op_bits_base_vp_valid ? _GEN_8429 : _GEN_8149; // @[sequencer-master.scala 320:41]
  wire  _GEN_8470 = io_op_bits_base_vp_valid ? _GEN_8430 : _GEN_8150; // @[sequencer-master.scala 320:41]
  wire  _GEN_8471 = io_op_bits_base_vp_valid ? _GEN_8431 : _GEN_8151; // @[sequencer-master.scala 320:41]
  wire  _GEN_8472 = io_op_bits_base_vp_valid ? _GEN_8432 : _GEN_7934; // @[sequencer-master.scala 320:41]
  wire  _GEN_8473 = io_op_bits_base_vp_valid ? _GEN_8433 : _GEN_7935; // @[sequencer-master.scala 320:41]
  wire  _GEN_8474 = io_op_bits_base_vp_valid ? _GEN_8434 : _GEN_7936; // @[sequencer-master.scala 320:41]
  wire  _GEN_8475 = io_op_bits_base_vp_valid ? _GEN_8435 : _GEN_7937; // @[sequencer-master.scala 320:41]
  wire  _GEN_8476 = io_op_bits_base_vp_valid ? _GEN_8436 : _GEN_7938; // @[sequencer-master.scala 320:41]
  wire  _GEN_8477 = io_op_bits_base_vp_valid ? _GEN_8437 : _GEN_7939; // @[sequencer-master.scala 320:41]
  wire  _GEN_8478 = io_op_bits_base_vp_valid ? _GEN_8438 : _GEN_7940; // @[sequencer-master.scala 320:41]
  wire  _GEN_8479 = io_op_bits_base_vp_valid ? _GEN_8439 : _GEN_7941; // @[sequencer-master.scala 320:41]
  wire  _GEN_8480 = io_op_bits_base_vp_valid ? _GEN_8440 : _GEN_7942; // @[sequencer-master.scala 320:41]
  wire  _GEN_8481 = io_op_bits_base_vp_valid ? _GEN_8441 : _GEN_7943; // @[sequencer-master.scala 320:41]
  wire  _GEN_8482 = io_op_bits_base_vp_valid ? _GEN_8442 : _GEN_7944; // @[sequencer-master.scala 320:41]
  wire  _GEN_8483 = io_op_bits_base_vp_valid ? _GEN_8443 : _GEN_7945; // @[sequencer-master.scala 320:41]
  wire  _GEN_8484 = io_op_bits_base_vp_valid ? _GEN_8444 : _GEN_7946; // @[sequencer-master.scala 320:41]
  wire  _GEN_8485 = io_op_bits_base_vp_valid ? _GEN_8445 : _GEN_7947; // @[sequencer-master.scala 320:41]
  wire  _GEN_8486 = io_op_bits_base_vp_valid ? _GEN_8446 : _GEN_7948; // @[sequencer-master.scala 320:41]
  wire  _GEN_8487 = io_op_bits_base_vp_valid ? _GEN_8447 : _GEN_7949; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8488 = io_op_bits_base_vp_valid ? _GEN_8448 : _GEN_7950; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8489 = io_op_bits_base_vp_valid ? _GEN_8449 : _GEN_7951; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8490 = io_op_bits_base_vp_valid ? _GEN_8450 : _GEN_7952; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8491 = io_op_bits_base_vp_valid ? _GEN_8451 : _GEN_7953; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8492 = io_op_bits_base_vp_valid ? _GEN_8452 : _GEN_7954; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8493 = io_op_bits_base_vp_valid ? _GEN_8453 : _GEN_7955; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8494 = io_op_bits_base_vp_valid ? _GEN_8454 : _GEN_7956; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_8495 = io_op_bits_base_vp_valid ? _GEN_8455 : _GEN_7957; // @[sequencer-master.scala 320:41]
  wire  _GEN_8496 = _GEN_32729 | _GEN_8192; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8497 = _GEN_32730 | _GEN_8193; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8498 = _GEN_32731 | _GEN_8194; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8499 = _GEN_32732 | _GEN_8195; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8500 = _GEN_32733 | _GEN_8196; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8501 = _GEN_32734 | _GEN_8197; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8502 = _GEN_32735 | _GEN_8198; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8503 = _GEN_32736 | _GEN_8199; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8504 = _T_26 ? _GEN_8496 : _GEN_8192; // @[sequencer-master.scala 154:24]
  wire  _GEN_8505 = _T_26 ? _GEN_8497 : _GEN_8193; // @[sequencer-master.scala 154:24]
  wire  _GEN_8506 = _T_26 ? _GEN_8498 : _GEN_8194; // @[sequencer-master.scala 154:24]
  wire  _GEN_8507 = _T_26 ? _GEN_8499 : _GEN_8195; // @[sequencer-master.scala 154:24]
  wire  _GEN_8508 = _T_26 ? _GEN_8500 : _GEN_8196; // @[sequencer-master.scala 154:24]
  wire  _GEN_8509 = _T_26 ? _GEN_8501 : _GEN_8197; // @[sequencer-master.scala 154:24]
  wire  _GEN_8510 = _T_26 ? _GEN_8502 : _GEN_8198; // @[sequencer-master.scala 154:24]
  wire  _GEN_8511 = _T_26 ? _GEN_8503 : _GEN_8199; // @[sequencer-master.scala 154:24]
  wire  _GEN_8512 = _GEN_32729 | _GEN_8216; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8513 = _GEN_32730 | _GEN_8217; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8514 = _GEN_32731 | _GEN_8218; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8515 = _GEN_32732 | _GEN_8219; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8516 = _GEN_32733 | _GEN_8220; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8517 = _GEN_32734 | _GEN_8221; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8518 = _GEN_32735 | _GEN_8222; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8519 = _GEN_32736 | _GEN_8223; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8520 = _T_48 ? _GEN_8512 : _GEN_8216; // @[sequencer-master.scala 154:24]
  wire  _GEN_8521 = _T_48 ? _GEN_8513 : _GEN_8217; // @[sequencer-master.scala 154:24]
  wire  _GEN_8522 = _T_48 ? _GEN_8514 : _GEN_8218; // @[sequencer-master.scala 154:24]
  wire  _GEN_8523 = _T_48 ? _GEN_8515 : _GEN_8219; // @[sequencer-master.scala 154:24]
  wire  _GEN_8524 = _T_48 ? _GEN_8516 : _GEN_8220; // @[sequencer-master.scala 154:24]
  wire  _GEN_8525 = _T_48 ? _GEN_8517 : _GEN_8221; // @[sequencer-master.scala 154:24]
  wire  _GEN_8526 = _T_48 ? _GEN_8518 : _GEN_8222; // @[sequencer-master.scala 154:24]
  wire  _GEN_8527 = _T_48 ? _GEN_8519 : _GEN_8223; // @[sequencer-master.scala 154:24]
  wire  _GEN_8528 = _GEN_32729 | _GEN_8240; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8529 = _GEN_32730 | _GEN_8241; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8530 = _GEN_32731 | _GEN_8242; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8531 = _GEN_32732 | _GEN_8243; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8532 = _GEN_32733 | _GEN_8244; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8533 = _GEN_32734 | _GEN_8245; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8534 = _GEN_32735 | _GEN_8246; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8535 = _GEN_32736 | _GEN_8247; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8536 = _T_70 ? _GEN_8528 : _GEN_8240; // @[sequencer-master.scala 154:24]
  wire  _GEN_8537 = _T_70 ? _GEN_8529 : _GEN_8241; // @[sequencer-master.scala 154:24]
  wire  _GEN_8538 = _T_70 ? _GEN_8530 : _GEN_8242; // @[sequencer-master.scala 154:24]
  wire  _GEN_8539 = _T_70 ? _GEN_8531 : _GEN_8243; // @[sequencer-master.scala 154:24]
  wire  _GEN_8540 = _T_70 ? _GEN_8532 : _GEN_8244; // @[sequencer-master.scala 154:24]
  wire  _GEN_8541 = _T_70 ? _GEN_8533 : _GEN_8245; // @[sequencer-master.scala 154:24]
  wire  _GEN_8542 = _T_70 ? _GEN_8534 : _GEN_8246; // @[sequencer-master.scala 154:24]
  wire  _GEN_8543 = _T_70 ? _GEN_8535 : _GEN_8247; // @[sequencer-master.scala 154:24]
  wire  _GEN_8544 = _GEN_32729 | _GEN_8264; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8545 = _GEN_32730 | _GEN_8265; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8546 = _GEN_32731 | _GEN_8266; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8547 = _GEN_32732 | _GEN_8267; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8548 = _GEN_32733 | _GEN_8268; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8549 = _GEN_32734 | _GEN_8269; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8550 = _GEN_32735 | _GEN_8270; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8551 = _GEN_32736 | _GEN_8271; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8552 = _T_92 ? _GEN_8544 : _GEN_8264; // @[sequencer-master.scala 154:24]
  wire  _GEN_8553 = _T_92 ? _GEN_8545 : _GEN_8265; // @[sequencer-master.scala 154:24]
  wire  _GEN_8554 = _T_92 ? _GEN_8546 : _GEN_8266; // @[sequencer-master.scala 154:24]
  wire  _GEN_8555 = _T_92 ? _GEN_8547 : _GEN_8267; // @[sequencer-master.scala 154:24]
  wire  _GEN_8556 = _T_92 ? _GEN_8548 : _GEN_8268; // @[sequencer-master.scala 154:24]
  wire  _GEN_8557 = _T_92 ? _GEN_8549 : _GEN_8269; // @[sequencer-master.scala 154:24]
  wire  _GEN_8558 = _T_92 ? _GEN_8550 : _GEN_8270; // @[sequencer-master.scala 154:24]
  wire  _GEN_8559 = _T_92 ? _GEN_8551 : _GEN_8271; // @[sequencer-master.scala 154:24]
  wire  _GEN_8560 = _GEN_32729 | _GEN_8288; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8561 = _GEN_32730 | _GEN_8289; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8562 = _GEN_32731 | _GEN_8290; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8563 = _GEN_32732 | _GEN_8291; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8564 = _GEN_32733 | _GEN_8292; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8565 = _GEN_32734 | _GEN_8293; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8566 = _GEN_32735 | _GEN_8294; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8567 = _GEN_32736 | _GEN_8295; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8568 = _T_114 ? _GEN_8560 : _GEN_8288; // @[sequencer-master.scala 154:24]
  wire  _GEN_8569 = _T_114 ? _GEN_8561 : _GEN_8289; // @[sequencer-master.scala 154:24]
  wire  _GEN_8570 = _T_114 ? _GEN_8562 : _GEN_8290; // @[sequencer-master.scala 154:24]
  wire  _GEN_8571 = _T_114 ? _GEN_8563 : _GEN_8291; // @[sequencer-master.scala 154:24]
  wire  _GEN_8572 = _T_114 ? _GEN_8564 : _GEN_8292; // @[sequencer-master.scala 154:24]
  wire  _GEN_8573 = _T_114 ? _GEN_8565 : _GEN_8293; // @[sequencer-master.scala 154:24]
  wire  _GEN_8574 = _T_114 ? _GEN_8566 : _GEN_8294; // @[sequencer-master.scala 154:24]
  wire  _GEN_8575 = _T_114 ? _GEN_8567 : _GEN_8295; // @[sequencer-master.scala 154:24]
  wire  _GEN_8576 = _GEN_32729 | _GEN_8312; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8577 = _GEN_32730 | _GEN_8313; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8578 = _GEN_32731 | _GEN_8314; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8579 = _GEN_32732 | _GEN_8315; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8580 = _GEN_32733 | _GEN_8316; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8581 = _GEN_32734 | _GEN_8317; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8582 = _GEN_32735 | _GEN_8318; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8583 = _GEN_32736 | _GEN_8319; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8584 = _T_136 ? _GEN_8576 : _GEN_8312; // @[sequencer-master.scala 154:24]
  wire  _GEN_8585 = _T_136 ? _GEN_8577 : _GEN_8313; // @[sequencer-master.scala 154:24]
  wire  _GEN_8586 = _T_136 ? _GEN_8578 : _GEN_8314; // @[sequencer-master.scala 154:24]
  wire  _GEN_8587 = _T_136 ? _GEN_8579 : _GEN_8315; // @[sequencer-master.scala 154:24]
  wire  _GEN_8588 = _T_136 ? _GEN_8580 : _GEN_8316; // @[sequencer-master.scala 154:24]
  wire  _GEN_8589 = _T_136 ? _GEN_8581 : _GEN_8317; // @[sequencer-master.scala 154:24]
  wire  _GEN_8590 = _T_136 ? _GEN_8582 : _GEN_8318; // @[sequencer-master.scala 154:24]
  wire  _GEN_8591 = _T_136 ? _GEN_8583 : _GEN_8319; // @[sequencer-master.scala 154:24]
  wire  _GEN_8592 = _GEN_32729 | _GEN_8336; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8593 = _GEN_32730 | _GEN_8337; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8594 = _GEN_32731 | _GEN_8338; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8595 = _GEN_32732 | _GEN_8339; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8596 = _GEN_32733 | _GEN_8340; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8597 = _GEN_32734 | _GEN_8341; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8598 = _GEN_32735 | _GEN_8342; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8599 = _GEN_32736 | _GEN_8343; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8600 = _T_158 ? _GEN_8592 : _GEN_8336; // @[sequencer-master.scala 154:24]
  wire  _GEN_8601 = _T_158 ? _GEN_8593 : _GEN_8337; // @[sequencer-master.scala 154:24]
  wire  _GEN_8602 = _T_158 ? _GEN_8594 : _GEN_8338; // @[sequencer-master.scala 154:24]
  wire  _GEN_8603 = _T_158 ? _GEN_8595 : _GEN_8339; // @[sequencer-master.scala 154:24]
  wire  _GEN_8604 = _T_158 ? _GEN_8596 : _GEN_8340; // @[sequencer-master.scala 154:24]
  wire  _GEN_8605 = _T_158 ? _GEN_8597 : _GEN_8341; // @[sequencer-master.scala 154:24]
  wire  _GEN_8606 = _T_158 ? _GEN_8598 : _GEN_8342; // @[sequencer-master.scala 154:24]
  wire  _GEN_8607 = _T_158 ? _GEN_8599 : _GEN_8343; // @[sequencer-master.scala 154:24]
  wire  _GEN_8608 = _GEN_32729 | _GEN_8360; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8609 = _GEN_32730 | _GEN_8361; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8610 = _GEN_32731 | _GEN_8362; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8611 = _GEN_32732 | _GEN_8363; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8612 = _GEN_32733 | _GEN_8364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8613 = _GEN_32734 | _GEN_8365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8614 = _GEN_32735 | _GEN_8366; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8615 = _GEN_32736 | _GEN_8367; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8616 = _T_180 ? _GEN_8608 : _GEN_8360; // @[sequencer-master.scala 154:24]
  wire  _GEN_8617 = _T_180 ? _GEN_8609 : _GEN_8361; // @[sequencer-master.scala 154:24]
  wire  _GEN_8618 = _T_180 ? _GEN_8610 : _GEN_8362; // @[sequencer-master.scala 154:24]
  wire  _GEN_8619 = _T_180 ? _GEN_8611 : _GEN_8363; // @[sequencer-master.scala 154:24]
  wire  _GEN_8620 = _T_180 ? _GEN_8612 : _GEN_8364; // @[sequencer-master.scala 154:24]
  wire  _GEN_8621 = _T_180 ? _GEN_8613 : _GEN_8365; // @[sequencer-master.scala 154:24]
  wire  _GEN_8622 = _T_180 ? _GEN_8614 : _GEN_8366; // @[sequencer-master.scala 154:24]
  wire  _GEN_8623 = _T_180 ? _GEN_8615 : _GEN_8367; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_8624 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_7958; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8625 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_7959; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8626 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_7960; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8627 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_7961; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8628 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_7962; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8629 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_7963; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8630 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_7964; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8631 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_7965; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8632 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_8152; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8633 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_8153; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8634 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_8154; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8635 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_8155; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8636 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_8156; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8637 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_8157; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8638 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_8158; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8639 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_8159; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8640 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_7966; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8641 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_7967; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8642 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_7968; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8643 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_7969; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8644 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_7970; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8645 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_7971; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8646 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_7972; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8647 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_7973; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8648 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_7974; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8649 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_7975; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8650 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_7976; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8651 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_7977; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8652 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_7978; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8653 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_7979; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8654 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_7980; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8655 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_7981; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8656 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_7982; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8657 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_7983; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8658 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_7984; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8659 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_7985; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8660 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_7986; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8661 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_7987; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8662 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_7988; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8663 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_7989; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8664 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_7990; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8665 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_7991; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8666 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_7992; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8667 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_7993; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8668 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_7994; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8669 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_7995; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8670 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_7996; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8671 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_7997; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_8672 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_7998; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8673 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_7999; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8674 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_8000; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8675 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_8001; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8676 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_8002; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8677 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_8003; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8678 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_8004; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8679 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_8005; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8680 = _T_189 ? _GEN_8672 : _GEN_7998; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8681 = _T_189 ? _GEN_8673 : _GEN_7999; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8682 = _T_189 ? _GEN_8674 : _GEN_8000; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8683 = _T_189 ? _GEN_8675 : _GEN_8001; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8684 = _T_189 ? _GEN_8676 : _GEN_8002; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8685 = _T_189 ? _GEN_8677 : _GEN_8003; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8686 = _T_189 ? _GEN_8678 : _GEN_8004; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8687 = _T_189 ? _GEN_8679 : _GEN_8005; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_8688 = io_op_bits_base_vs1_valid ? _GEN_8624 : _GEN_7958; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8689 = io_op_bits_base_vs1_valid ? _GEN_8625 : _GEN_7959; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8690 = io_op_bits_base_vs1_valid ? _GEN_8626 : _GEN_7960; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8691 = io_op_bits_base_vs1_valid ? _GEN_8627 : _GEN_7961; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8692 = io_op_bits_base_vs1_valid ? _GEN_8628 : _GEN_7962; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8693 = io_op_bits_base_vs1_valid ? _GEN_8629 : _GEN_7963; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8694 = io_op_bits_base_vs1_valid ? _GEN_8630 : _GEN_7964; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8695 = io_op_bits_base_vs1_valid ? _GEN_8631 : _GEN_7965; // @[sequencer-master.scala 328:47]
  wire  _GEN_8696 = io_op_bits_base_vs1_valid ? _GEN_8632 : _GEN_8152; // @[sequencer-master.scala 328:47]
  wire  _GEN_8697 = io_op_bits_base_vs1_valid ? _GEN_8633 : _GEN_8153; // @[sequencer-master.scala 328:47]
  wire  _GEN_8698 = io_op_bits_base_vs1_valid ? _GEN_8634 : _GEN_8154; // @[sequencer-master.scala 328:47]
  wire  _GEN_8699 = io_op_bits_base_vs1_valid ? _GEN_8635 : _GEN_8155; // @[sequencer-master.scala 328:47]
  wire  _GEN_8700 = io_op_bits_base_vs1_valid ? _GEN_8636 : _GEN_8156; // @[sequencer-master.scala 328:47]
  wire  _GEN_8701 = io_op_bits_base_vs1_valid ? _GEN_8637 : _GEN_8157; // @[sequencer-master.scala 328:47]
  wire  _GEN_8702 = io_op_bits_base_vs1_valid ? _GEN_8638 : _GEN_8158; // @[sequencer-master.scala 328:47]
  wire  _GEN_8703 = io_op_bits_base_vs1_valid ? _GEN_8639 : _GEN_8159; // @[sequencer-master.scala 328:47]
  wire  _GEN_8704 = io_op_bits_base_vs1_valid ? _GEN_8640 : _GEN_7966; // @[sequencer-master.scala 328:47]
  wire  _GEN_8705 = io_op_bits_base_vs1_valid ? _GEN_8641 : _GEN_7967; // @[sequencer-master.scala 328:47]
  wire  _GEN_8706 = io_op_bits_base_vs1_valid ? _GEN_8642 : _GEN_7968; // @[sequencer-master.scala 328:47]
  wire  _GEN_8707 = io_op_bits_base_vs1_valid ? _GEN_8643 : _GEN_7969; // @[sequencer-master.scala 328:47]
  wire  _GEN_8708 = io_op_bits_base_vs1_valid ? _GEN_8644 : _GEN_7970; // @[sequencer-master.scala 328:47]
  wire  _GEN_8709 = io_op_bits_base_vs1_valid ? _GEN_8645 : _GEN_7971; // @[sequencer-master.scala 328:47]
  wire  _GEN_8710 = io_op_bits_base_vs1_valid ? _GEN_8646 : _GEN_7972; // @[sequencer-master.scala 328:47]
  wire  _GEN_8711 = io_op_bits_base_vs1_valid ? _GEN_8647 : _GEN_7973; // @[sequencer-master.scala 328:47]
  wire  _GEN_8712 = io_op_bits_base_vs1_valid ? _GEN_8648 : _GEN_7974; // @[sequencer-master.scala 328:47]
  wire  _GEN_8713 = io_op_bits_base_vs1_valid ? _GEN_8649 : _GEN_7975; // @[sequencer-master.scala 328:47]
  wire  _GEN_8714 = io_op_bits_base_vs1_valid ? _GEN_8650 : _GEN_7976; // @[sequencer-master.scala 328:47]
  wire  _GEN_8715 = io_op_bits_base_vs1_valid ? _GEN_8651 : _GEN_7977; // @[sequencer-master.scala 328:47]
  wire  _GEN_8716 = io_op_bits_base_vs1_valid ? _GEN_8652 : _GEN_7978; // @[sequencer-master.scala 328:47]
  wire  _GEN_8717 = io_op_bits_base_vs1_valid ? _GEN_8653 : _GEN_7979; // @[sequencer-master.scala 328:47]
  wire  _GEN_8718 = io_op_bits_base_vs1_valid ? _GEN_8654 : _GEN_7980; // @[sequencer-master.scala 328:47]
  wire  _GEN_8719 = io_op_bits_base_vs1_valid ? _GEN_8655 : _GEN_7981; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8720 = io_op_bits_base_vs1_valid ? _GEN_8656 : _GEN_7982; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8721 = io_op_bits_base_vs1_valid ? _GEN_8657 : _GEN_7983; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8722 = io_op_bits_base_vs1_valid ? _GEN_8658 : _GEN_7984; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8723 = io_op_bits_base_vs1_valid ? _GEN_8659 : _GEN_7985; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8724 = io_op_bits_base_vs1_valid ? _GEN_8660 : _GEN_7986; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8725 = io_op_bits_base_vs1_valid ? _GEN_8661 : _GEN_7987; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8726 = io_op_bits_base_vs1_valid ? _GEN_8662 : _GEN_7988; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8727 = io_op_bits_base_vs1_valid ? _GEN_8663 : _GEN_7989; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8728 = io_op_bits_base_vs1_valid ? _GEN_8664 : _GEN_7990; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8729 = io_op_bits_base_vs1_valid ? _GEN_8665 : _GEN_7991; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8730 = io_op_bits_base_vs1_valid ? _GEN_8666 : _GEN_7992; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8731 = io_op_bits_base_vs1_valid ? _GEN_8667 : _GEN_7993; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8732 = io_op_bits_base_vs1_valid ? _GEN_8668 : _GEN_7994; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8733 = io_op_bits_base_vs1_valid ? _GEN_8669 : _GEN_7995; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8734 = io_op_bits_base_vs1_valid ? _GEN_8670 : _GEN_7996; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8735 = io_op_bits_base_vs1_valid ? _GEN_8671 : _GEN_7997; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8736 = io_op_bits_base_vs1_valid ? _GEN_8680 : _GEN_7998; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8737 = io_op_bits_base_vs1_valid ? _GEN_8681 : _GEN_7999; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8738 = io_op_bits_base_vs1_valid ? _GEN_8682 : _GEN_8000; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8739 = io_op_bits_base_vs1_valid ? _GEN_8683 : _GEN_8001; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8740 = io_op_bits_base_vs1_valid ? _GEN_8684 : _GEN_8002; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8741 = io_op_bits_base_vs1_valid ? _GEN_8685 : _GEN_8003; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8742 = io_op_bits_base_vs1_valid ? _GEN_8686 : _GEN_8004; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8743 = io_op_bits_base_vs1_valid ? _GEN_8687 : _GEN_8005; // @[sequencer-master.scala 328:47]
  wire  _GEN_8744 = _GEN_32729 | _GEN_8504; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8745 = _GEN_32730 | _GEN_8505; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8746 = _GEN_32731 | _GEN_8506; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8747 = _GEN_32732 | _GEN_8507; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8748 = _GEN_32733 | _GEN_8508; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8749 = _GEN_32734 | _GEN_8509; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8750 = _GEN_32735 | _GEN_8510; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8751 = _GEN_32736 | _GEN_8511; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8752 = _T_203 ? _GEN_8744 : _GEN_8504; // @[sequencer-master.scala 154:24]
  wire  _GEN_8753 = _T_203 ? _GEN_8745 : _GEN_8505; // @[sequencer-master.scala 154:24]
  wire  _GEN_8754 = _T_203 ? _GEN_8746 : _GEN_8506; // @[sequencer-master.scala 154:24]
  wire  _GEN_8755 = _T_203 ? _GEN_8747 : _GEN_8507; // @[sequencer-master.scala 154:24]
  wire  _GEN_8756 = _T_203 ? _GEN_8748 : _GEN_8508; // @[sequencer-master.scala 154:24]
  wire  _GEN_8757 = _T_203 ? _GEN_8749 : _GEN_8509; // @[sequencer-master.scala 154:24]
  wire  _GEN_8758 = _T_203 ? _GEN_8750 : _GEN_8510; // @[sequencer-master.scala 154:24]
  wire  _GEN_8759 = _T_203 ? _GEN_8751 : _GEN_8511; // @[sequencer-master.scala 154:24]
  wire  _GEN_8760 = _GEN_32729 | _GEN_8520; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8761 = _GEN_32730 | _GEN_8521; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8762 = _GEN_32731 | _GEN_8522; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8763 = _GEN_32732 | _GEN_8523; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8764 = _GEN_32733 | _GEN_8524; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8765 = _GEN_32734 | _GEN_8525; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8766 = _GEN_32735 | _GEN_8526; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8767 = _GEN_32736 | _GEN_8527; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8768 = _T_225 ? _GEN_8760 : _GEN_8520; // @[sequencer-master.scala 154:24]
  wire  _GEN_8769 = _T_225 ? _GEN_8761 : _GEN_8521; // @[sequencer-master.scala 154:24]
  wire  _GEN_8770 = _T_225 ? _GEN_8762 : _GEN_8522; // @[sequencer-master.scala 154:24]
  wire  _GEN_8771 = _T_225 ? _GEN_8763 : _GEN_8523; // @[sequencer-master.scala 154:24]
  wire  _GEN_8772 = _T_225 ? _GEN_8764 : _GEN_8524; // @[sequencer-master.scala 154:24]
  wire  _GEN_8773 = _T_225 ? _GEN_8765 : _GEN_8525; // @[sequencer-master.scala 154:24]
  wire  _GEN_8774 = _T_225 ? _GEN_8766 : _GEN_8526; // @[sequencer-master.scala 154:24]
  wire  _GEN_8775 = _T_225 ? _GEN_8767 : _GEN_8527; // @[sequencer-master.scala 154:24]
  wire  _GEN_8776 = _GEN_32729 | _GEN_8536; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8777 = _GEN_32730 | _GEN_8537; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8778 = _GEN_32731 | _GEN_8538; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8779 = _GEN_32732 | _GEN_8539; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8780 = _GEN_32733 | _GEN_8540; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8781 = _GEN_32734 | _GEN_8541; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8782 = _GEN_32735 | _GEN_8542; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8783 = _GEN_32736 | _GEN_8543; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8784 = _T_247 ? _GEN_8776 : _GEN_8536; // @[sequencer-master.scala 154:24]
  wire  _GEN_8785 = _T_247 ? _GEN_8777 : _GEN_8537; // @[sequencer-master.scala 154:24]
  wire  _GEN_8786 = _T_247 ? _GEN_8778 : _GEN_8538; // @[sequencer-master.scala 154:24]
  wire  _GEN_8787 = _T_247 ? _GEN_8779 : _GEN_8539; // @[sequencer-master.scala 154:24]
  wire  _GEN_8788 = _T_247 ? _GEN_8780 : _GEN_8540; // @[sequencer-master.scala 154:24]
  wire  _GEN_8789 = _T_247 ? _GEN_8781 : _GEN_8541; // @[sequencer-master.scala 154:24]
  wire  _GEN_8790 = _T_247 ? _GEN_8782 : _GEN_8542; // @[sequencer-master.scala 154:24]
  wire  _GEN_8791 = _T_247 ? _GEN_8783 : _GEN_8543; // @[sequencer-master.scala 154:24]
  wire  _GEN_8792 = _GEN_32729 | _GEN_8552; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8793 = _GEN_32730 | _GEN_8553; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8794 = _GEN_32731 | _GEN_8554; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8795 = _GEN_32732 | _GEN_8555; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8796 = _GEN_32733 | _GEN_8556; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8797 = _GEN_32734 | _GEN_8557; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8798 = _GEN_32735 | _GEN_8558; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8799 = _GEN_32736 | _GEN_8559; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8800 = _T_269 ? _GEN_8792 : _GEN_8552; // @[sequencer-master.scala 154:24]
  wire  _GEN_8801 = _T_269 ? _GEN_8793 : _GEN_8553; // @[sequencer-master.scala 154:24]
  wire  _GEN_8802 = _T_269 ? _GEN_8794 : _GEN_8554; // @[sequencer-master.scala 154:24]
  wire  _GEN_8803 = _T_269 ? _GEN_8795 : _GEN_8555; // @[sequencer-master.scala 154:24]
  wire  _GEN_8804 = _T_269 ? _GEN_8796 : _GEN_8556; // @[sequencer-master.scala 154:24]
  wire  _GEN_8805 = _T_269 ? _GEN_8797 : _GEN_8557; // @[sequencer-master.scala 154:24]
  wire  _GEN_8806 = _T_269 ? _GEN_8798 : _GEN_8558; // @[sequencer-master.scala 154:24]
  wire  _GEN_8807 = _T_269 ? _GEN_8799 : _GEN_8559; // @[sequencer-master.scala 154:24]
  wire  _GEN_8808 = _GEN_32729 | _GEN_8568; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8809 = _GEN_32730 | _GEN_8569; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8810 = _GEN_32731 | _GEN_8570; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8811 = _GEN_32732 | _GEN_8571; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8812 = _GEN_32733 | _GEN_8572; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8813 = _GEN_32734 | _GEN_8573; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8814 = _GEN_32735 | _GEN_8574; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8815 = _GEN_32736 | _GEN_8575; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8816 = _T_291 ? _GEN_8808 : _GEN_8568; // @[sequencer-master.scala 154:24]
  wire  _GEN_8817 = _T_291 ? _GEN_8809 : _GEN_8569; // @[sequencer-master.scala 154:24]
  wire  _GEN_8818 = _T_291 ? _GEN_8810 : _GEN_8570; // @[sequencer-master.scala 154:24]
  wire  _GEN_8819 = _T_291 ? _GEN_8811 : _GEN_8571; // @[sequencer-master.scala 154:24]
  wire  _GEN_8820 = _T_291 ? _GEN_8812 : _GEN_8572; // @[sequencer-master.scala 154:24]
  wire  _GEN_8821 = _T_291 ? _GEN_8813 : _GEN_8573; // @[sequencer-master.scala 154:24]
  wire  _GEN_8822 = _T_291 ? _GEN_8814 : _GEN_8574; // @[sequencer-master.scala 154:24]
  wire  _GEN_8823 = _T_291 ? _GEN_8815 : _GEN_8575; // @[sequencer-master.scala 154:24]
  wire  _GEN_8824 = _GEN_32729 | _GEN_8584; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8825 = _GEN_32730 | _GEN_8585; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8826 = _GEN_32731 | _GEN_8586; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8827 = _GEN_32732 | _GEN_8587; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8828 = _GEN_32733 | _GEN_8588; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8829 = _GEN_32734 | _GEN_8589; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8830 = _GEN_32735 | _GEN_8590; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8831 = _GEN_32736 | _GEN_8591; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8832 = _T_313 ? _GEN_8824 : _GEN_8584; // @[sequencer-master.scala 154:24]
  wire  _GEN_8833 = _T_313 ? _GEN_8825 : _GEN_8585; // @[sequencer-master.scala 154:24]
  wire  _GEN_8834 = _T_313 ? _GEN_8826 : _GEN_8586; // @[sequencer-master.scala 154:24]
  wire  _GEN_8835 = _T_313 ? _GEN_8827 : _GEN_8587; // @[sequencer-master.scala 154:24]
  wire  _GEN_8836 = _T_313 ? _GEN_8828 : _GEN_8588; // @[sequencer-master.scala 154:24]
  wire  _GEN_8837 = _T_313 ? _GEN_8829 : _GEN_8589; // @[sequencer-master.scala 154:24]
  wire  _GEN_8838 = _T_313 ? _GEN_8830 : _GEN_8590; // @[sequencer-master.scala 154:24]
  wire  _GEN_8839 = _T_313 ? _GEN_8831 : _GEN_8591; // @[sequencer-master.scala 154:24]
  wire  _GEN_8840 = _GEN_32729 | _GEN_8600; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8841 = _GEN_32730 | _GEN_8601; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8842 = _GEN_32731 | _GEN_8602; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8843 = _GEN_32732 | _GEN_8603; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8844 = _GEN_32733 | _GEN_8604; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8845 = _GEN_32734 | _GEN_8605; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8846 = _GEN_32735 | _GEN_8606; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8847 = _GEN_32736 | _GEN_8607; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8848 = _T_335 ? _GEN_8840 : _GEN_8600; // @[sequencer-master.scala 154:24]
  wire  _GEN_8849 = _T_335 ? _GEN_8841 : _GEN_8601; // @[sequencer-master.scala 154:24]
  wire  _GEN_8850 = _T_335 ? _GEN_8842 : _GEN_8602; // @[sequencer-master.scala 154:24]
  wire  _GEN_8851 = _T_335 ? _GEN_8843 : _GEN_8603; // @[sequencer-master.scala 154:24]
  wire  _GEN_8852 = _T_335 ? _GEN_8844 : _GEN_8604; // @[sequencer-master.scala 154:24]
  wire  _GEN_8853 = _T_335 ? _GEN_8845 : _GEN_8605; // @[sequencer-master.scala 154:24]
  wire  _GEN_8854 = _T_335 ? _GEN_8846 : _GEN_8606; // @[sequencer-master.scala 154:24]
  wire  _GEN_8855 = _T_335 ? _GEN_8847 : _GEN_8607; // @[sequencer-master.scala 154:24]
  wire  _GEN_8856 = _GEN_32729 | _GEN_8616; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8857 = _GEN_32730 | _GEN_8617; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8858 = _GEN_32731 | _GEN_8618; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8859 = _GEN_32732 | _GEN_8619; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8860 = _GEN_32733 | _GEN_8620; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8861 = _GEN_32734 | _GEN_8621; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8862 = _GEN_32735 | _GEN_8622; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8863 = _GEN_32736 | _GEN_8623; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8864 = _T_357 ? _GEN_8856 : _GEN_8616; // @[sequencer-master.scala 154:24]
  wire  _GEN_8865 = _T_357 ? _GEN_8857 : _GEN_8617; // @[sequencer-master.scala 154:24]
  wire  _GEN_8866 = _T_357 ? _GEN_8858 : _GEN_8618; // @[sequencer-master.scala 154:24]
  wire  _GEN_8867 = _T_357 ? _GEN_8859 : _GEN_8619; // @[sequencer-master.scala 154:24]
  wire  _GEN_8868 = _T_357 ? _GEN_8860 : _GEN_8620; // @[sequencer-master.scala 154:24]
  wire  _GEN_8869 = _T_357 ? _GEN_8861 : _GEN_8621; // @[sequencer-master.scala 154:24]
  wire  _GEN_8870 = _T_357 ? _GEN_8862 : _GEN_8622; // @[sequencer-master.scala 154:24]
  wire  _GEN_8871 = _T_357 ? _GEN_8863 : _GEN_8623; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_8872 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_8006; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8873 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_8007; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8874 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_8008; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8875 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_8009; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8876 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_8010; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8877 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_8011; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8878 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_8012; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8879 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_8013; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8880 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_8160; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8881 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_8161; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8882 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_8162; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8883 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_8163; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8884 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_8164; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8885 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_8165; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8886 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_8166; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8887 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_8167; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8888 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_8014; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8889 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_8015; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8890 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_8016; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8891 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_8017; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8892 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_8018; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8893 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_8019; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8894 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_8020; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8895 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_8021; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8896 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_8022; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8897 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_8023; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8898 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_8024; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8899 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_8025; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8900 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_8026; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8901 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_8027; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8902 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_8028; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_8903 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_8029; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8904 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_8030; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8905 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_8031; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8906 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_8032; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8907 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_8033; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8908 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_8034; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8909 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_8035; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8910 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_8036; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_8911 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_8037; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_8912 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_8038; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8913 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_8039; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8914 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_8040; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8915 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_8041; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8916 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_8042; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8917 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_8043; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8918 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_8044; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_8919 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_8045; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_8920 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_8046; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8921 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_8047; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8922 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_8048; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8923 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_8049; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8924 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_8050; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8925 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_8051; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8926 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_8052; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8927 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_8053; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_8928 = _T_366 ? _GEN_8920 : _GEN_8046; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8929 = _T_366 ? _GEN_8921 : _GEN_8047; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8930 = _T_366 ? _GEN_8922 : _GEN_8048; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8931 = _T_366 ? _GEN_8923 : _GEN_8049; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8932 = _T_366 ? _GEN_8924 : _GEN_8050; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8933 = _T_366 ? _GEN_8925 : _GEN_8051; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8934 = _T_366 ? _GEN_8926 : _GEN_8052; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_8935 = _T_366 ? _GEN_8927 : _GEN_8053; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_8936 = io_op_bits_base_vs2_valid ? _GEN_8872 : _GEN_8006; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8937 = io_op_bits_base_vs2_valid ? _GEN_8873 : _GEN_8007; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8938 = io_op_bits_base_vs2_valid ? _GEN_8874 : _GEN_8008; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8939 = io_op_bits_base_vs2_valid ? _GEN_8875 : _GEN_8009; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8940 = io_op_bits_base_vs2_valid ? _GEN_8876 : _GEN_8010; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8941 = io_op_bits_base_vs2_valid ? _GEN_8877 : _GEN_8011; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8942 = io_op_bits_base_vs2_valid ? _GEN_8878 : _GEN_8012; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8943 = io_op_bits_base_vs2_valid ? _GEN_8879 : _GEN_8013; // @[sequencer-master.scala 328:47]
  wire  _GEN_8944 = io_op_bits_base_vs2_valid ? _GEN_8880 : _GEN_8160; // @[sequencer-master.scala 328:47]
  wire  _GEN_8945 = io_op_bits_base_vs2_valid ? _GEN_8881 : _GEN_8161; // @[sequencer-master.scala 328:47]
  wire  _GEN_8946 = io_op_bits_base_vs2_valid ? _GEN_8882 : _GEN_8162; // @[sequencer-master.scala 328:47]
  wire  _GEN_8947 = io_op_bits_base_vs2_valid ? _GEN_8883 : _GEN_8163; // @[sequencer-master.scala 328:47]
  wire  _GEN_8948 = io_op_bits_base_vs2_valid ? _GEN_8884 : _GEN_8164; // @[sequencer-master.scala 328:47]
  wire  _GEN_8949 = io_op_bits_base_vs2_valid ? _GEN_8885 : _GEN_8165; // @[sequencer-master.scala 328:47]
  wire  _GEN_8950 = io_op_bits_base_vs2_valid ? _GEN_8886 : _GEN_8166; // @[sequencer-master.scala 328:47]
  wire  _GEN_8951 = io_op_bits_base_vs2_valid ? _GEN_8887 : _GEN_8167; // @[sequencer-master.scala 328:47]
  wire  _GEN_8952 = io_op_bits_base_vs2_valid ? _GEN_8888 : _GEN_8014; // @[sequencer-master.scala 328:47]
  wire  _GEN_8953 = io_op_bits_base_vs2_valid ? _GEN_8889 : _GEN_8015; // @[sequencer-master.scala 328:47]
  wire  _GEN_8954 = io_op_bits_base_vs2_valid ? _GEN_8890 : _GEN_8016; // @[sequencer-master.scala 328:47]
  wire  _GEN_8955 = io_op_bits_base_vs2_valid ? _GEN_8891 : _GEN_8017; // @[sequencer-master.scala 328:47]
  wire  _GEN_8956 = io_op_bits_base_vs2_valid ? _GEN_8892 : _GEN_8018; // @[sequencer-master.scala 328:47]
  wire  _GEN_8957 = io_op_bits_base_vs2_valid ? _GEN_8893 : _GEN_8019; // @[sequencer-master.scala 328:47]
  wire  _GEN_8958 = io_op_bits_base_vs2_valid ? _GEN_8894 : _GEN_8020; // @[sequencer-master.scala 328:47]
  wire  _GEN_8959 = io_op_bits_base_vs2_valid ? _GEN_8895 : _GEN_8021; // @[sequencer-master.scala 328:47]
  wire  _GEN_8960 = io_op_bits_base_vs2_valid ? _GEN_8896 : _GEN_8022; // @[sequencer-master.scala 328:47]
  wire  _GEN_8961 = io_op_bits_base_vs2_valid ? _GEN_8897 : _GEN_8023; // @[sequencer-master.scala 328:47]
  wire  _GEN_8962 = io_op_bits_base_vs2_valid ? _GEN_8898 : _GEN_8024; // @[sequencer-master.scala 328:47]
  wire  _GEN_8963 = io_op_bits_base_vs2_valid ? _GEN_8899 : _GEN_8025; // @[sequencer-master.scala 328:47]
  wire  _GEN_8964 = io_op_bits_base_vs2_valid ? _GEN_8900 : _GEN_8026; // @[sequencer-master.scala 328:47]
  wire  _GEN_8965 = io_op_bits_base_vs2_valid ? _GEN_8901 : _GEN_8027; // @[sequencer-master.scala 328:47]
  wire  _GEN_8966 = io_op_bits_base_vs2_valid ? _GEN_8902 : _GEN_8028; // @[sequencer-master.scala 328:47]
  wire  _GEN_8967 = io_op_bits_base_vs2_valid ? _GEN_8903 : _GEN_8029; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8968 = io_op_bits_base_vs2_valid ? _GEN_8904 : _GEN_8030; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8969 = io_op_bits_base_vs2_valid ? _GEN_8905 : _GEN_8031; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8970 = io_op_bits_base_vs2_valid ? _GEN_8906 : _GEN_8032; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8971 = io_op_bits_base_vs2_valid ? _GEN_8907 : _GEN_8033; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8972 = io_op_bits_base_vs2_valid ? _GEN_8908 : _GEN_8034; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8973 = io_op_bits_base_vs2_valid ? _GEN_8909 : _GEN_8035; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8974 = io_op_bits_base_vs2_valid ? _GEN_8910 : _GEN_8036; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_8975 = io_op_bits_base_vs2_valid ? _GEN_8911 : _GEN_8037; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8976 = io_op_bits_base_vs2_valid ? _GEN_8912 : _GEN_8038; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8977 = io_op_bits_base_vs2_valid ? _GEN_8913 : _GEN_8039; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8978 = io_op_bits_base_vs2_valid ? _GEN_8914 : _GEN_8040; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8979 = io_op_bits_base_vs2_valid ? _GEN_8915 : _GEN_8041; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8980 = io_op_bits_base_vs2_valid ? _GEN_8916 : _GEN_8042; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8981 = io_op_bits_base_vs2_valid ? _GEN_8917 : _GEN_8043; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8982 = io_op_bits_base_vs2_valid ? _GEN_8918 : _GEN_8044; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_8983 = io_op_bits_base_vs2_valid ? _GEN_8919 : _GEN_8045; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8984 = io_op_bits_base_vs2_valid ? _GEN_8928 : _GEN_8046; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8985 = io_op_bits_base_vs2_valid ? _GEN_8929 : _GEN_8047; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8986 = io_op_bits_base_vs2_valid ? _GEN_8930 : _GEN_8048; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8987 = io_op_bits_base_vs2_valid ? _GEN_8931 : _GEN_8049; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8988 = io_op_bits_base_vs2_valid ? _GEN_8932 : _GEN_8050; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8989 = io_op_bits_base_vs2_valid ? _GEN_8933 : _GEN_8051; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8990 = io_op_bits_base_vs2_valid ? _GEN_8934 : _GEN_8052; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_8991 = io_op_bits_base_vs2_valid ? _GEN_8935 : _GEN_8053; // @[sequencer-master.scala 328:47]
  wire  _GEN_8992 = _GEN_32729 | _GEN_8752; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8993 = _GEN_32730 | _GEN_8753; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8994 = _GEN_32731 | _GEN_8754; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8995 = _GEN_32732 | _GEN_8755; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8996 = _GEN_32733 | _GEN_8756; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8997 = _GEN_32734 | _GEN_8757; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8998 = _GEN_32735 | _GEN_8758; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_8999 = _GEN_32736 | _GEN_8759; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9000 = _T_380 ? _GEN_8992 : _GEN_8752; // @[sequencer-master.scala 154:24]
  wire  _GEN_9001 = _T_380 ? _GEN_8993 : _GEN_8753; // @[sequencer-master.scala 154:24]
  wire  _GEN_9002 = _T_380 ? _GEN_8994 : _GEN_8754; // @[sequencer-master.scala 154:24]
  wire  _GEN_9003 = _T_380 ? _GEN_8995 : _GEN_8755; // @[sequencer-master.scala 154:24]
  wire  _GEN_9004 = _T_380 ? _GEN_8996 : _GEN_8756; // @[sequencer-master.scala 154:24]
  wire  _GEN_9005 = _T_380 ? _GEN_8997 : _GEN_8757; // @[sequencer-master.scala 154:24]
  wire  _GEN_9006 = _T_380 ? _GEN_8998 : _GEN_8758; // @[sequencer-master.scala 154:24]
  wire  _GEN_9007 = _T_380 ? _GEN_8999 : _GEN_8759; // @[sequencer-master.scala 154:24]
  wire  _GEN_9008 = _GEN_32729 | _GEN_8768; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9009 = _GEN_32730 | _GEN_8769; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9010 = _GEN_32731 | _GEN_8770; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9011 = _GEN_32732 | _GEN_8771; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9012 = _GEN_32733 | _GEN_8772; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9013 = _GEN_32734 | _GEN_8773; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9014 = _GEN_32735 | _GEN_8774; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9015 = _GEN_32736 | _GEN_8775; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9016 = _T_402 ? _GEN_9008 : _GEN_8768; // @[sequencer-master.scala 154:24]
  wire  _GEN_9017 = _T_402 ? _GEN_9009 : _GEN_8769; // @[sequencer-master.scala 154:24]
  wire  _GEN_9018 = _T_402 ? _GEN_9010 : _GEN_8770; // @[sequencer-master.scala 154:24]
  wire  _GEN_9019 = _T_402 ? _GEN_9011 : _GEN_8771; // @[sequencer-master.scala 154:24]
  wire  _GEN_9020 = _T_402 ? _GEN_9012 : _GEN_8772; // @[sequencer-master.scala 154:24]
  wire  _GEN_9021 = _T_402 ? _GEN_9013 : _GEN_8773; // @[sequencer-master.scala 154:24]
  wire  _GEN_9022 = _T_402 ? _GEN_9014 : _GEN_8774; // @[sequencer-master.scala 154:24]
  wire  _GEN_9023 = _T_402 ? _GEN_9015 : _GEN_8775; // @[sequencer-master.scala 154:24]
  wire  _GEN_9024 = _GEN_32729 | _GEN_8784; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9025 = _GEN_32730 | _GEN_8785; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9026 = _GEN_32731 | _GEN_8786; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9027 = _GEN_32732 | _GEN_8787; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9028 = _GEN_32733 | _GEN_8788; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9029 = _GEN_32734 | _GEN_8789; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9030 = _GEN_32735 | _GEN_8790; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9031 = _GEN_32736 | _GEN_8791; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9032 = _T_424 ? _GEN_9024 : _GEN_8784; // @[sequencer-master.scala 154:24]
  wire  _GEN_9033 = _T_424 ? _GEN_9025 : _GEN_8785; // @[sequencer-master.scala 154:24]
  wire  _GEN_9034 = _T_424 ? _GEN_9026 : _GEN_8786; // @[sequencer-master.scala 154:24]
  wire  _GEN_9035 = _T_424 ? _GEN_9027 : _GEN_8787; // @[sequencer-master.scala 154:24]
  wire  _GEN_9036 = _T_424 ? _GEN_9028 : _GEN_8788; // @[sequencer-master.scala 154:24]
  wire  _GEN_9037 = _T_424 ? _GEN_9029 : _GEN_8789; // @[sequencer-master.scala 154:24]
  wire  _GEN_9038 = _T_424 ? _GEN_9030 : _GEN_8790; // @[sequencer-master.scala 154:24]
  wire  _GEN_9039 = _T_424 ? _GEN_9031 : _GEN_8791; // @[sequencer-master.scala 154:24]
  wire  _GEN_9040 = _GEN_32729 | _GEN_8800; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9041 = _GEN_32730 | _GEN_8801; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9042 = _GEN_32731 | _GEN_8802; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9043 = _GEN_32732 | _GEN_8803; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9044 = _GEN_32733 | _GEN_8804; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9045 = _GEN_32734 | _GEN_8805; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9046 = _GEN_32735 | _GEN_8806; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9047 = _GEN_32736 | _GEN_8807; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9048 = _T_446 ? _GEN_9040 : _GEN_8800; // @[sequencer-master.scala 154:24]
  wire  _GEN_9049 = _T_446 ? _GEN_9041 : _GEN_8801; // @[sequencer-master.scala 154:24]
  wire  _GEN_9050 = _T_446 ? _GEN_9042 : _GEN_8802; // @[sequencer-master.scala 154:24]
  wire  _GEN_9051 = _T_446 ? _GEN_9043 : _GEN_8803; // @[sequencer-master.scala 154:24]
  wire  _GEN_9052 = _T_446 ? _GEN_9044 : _GEN_8804; // @[sequencer-master.scala 154:24]
  wire  _GEN_9053 = _T_446 ? _GEN_9045 : _GEN_8805; // @[sequencer-master.scala 154:24]
  wire  _GEN_9054 = _T_446 ? _GEN_9046 : _GEN_8806; // @[sequencer-master.scala 154:24]
  wire  _GEN_9055 = _T_446 ? _GEN_9047 : _GEN_8807; // @[sequencer-master.scala 154:24]
  wire  _GEN_9056 = _GEN_32729 | _GEN_8816; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9057 = _GEN_32730 | _GEN_8817; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9058 = _GEN_32731 | _GEN_8818; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9059 = _GEN_32732 | _GEN_8819; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9060 = _GEN_32733 | _GEN_8820; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9061 = _GEN_32734 | _GEN_8821; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9062 = _GEN_32735 | _GEN_8822; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9063 = _GEN_32736 | _GEN_8823; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9064 = _T_468 ? _GEN_9056 : _GEN_8816; // @[sequencer-master.scala 154:24]
  wire  _GEN_9065 = _T_468 ? _GEN_9057 : _GEN_8817; // @[sequencer-master.scala 154:24]
  wire  _GEN_9066 = _T_468 ? _GEN_9058 : _GEN_8818; // @[sequencer-master.scala 154:24]
  wire  _GEN_9067 = _T_468 ? _GEN_9059 : _GEN_8819; // @[sequencer-master.scala 154:24]
  wire  _GEN_9068 = _T_468 ? _GEN_9060 : _GEN_8820; // @[sequencer-master.scala 154:24]
  wire  _GEN_9069 = _T_468 ? _GEN_9061 : _GEN_8821; // @[sequencer-master.scala 154:24]
  wire  _GEN_9070 = _T_468 ? _GEN_9062 : _GEN_8822; // @[sequencer-master.scala 154:24]
  wire  _GEN_9071 = _T_468 ? _GEN_9063 : _GEN_8823; // @[sequencer-master.scala 154:24]
  wire  _GEN_9072 = _GEN_32729 | _GEN_8832; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9073 = _GEN_32730 | _GEN_8833; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9074 = _GEN_32731 | _GEN_8834; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9075 = _GEN_32732 | _GEN_8835; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9076 = _GEN_32733 | _GEN_8836; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9077 = _GEN_32734 | _GEN_8837; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9078 = _GEN_32735 | _GEN_8838; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9079 = _GEN_32736 | _GEN_8839; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9080 = _T_490 ? _GEN_9072 : _GEN_8832; // @[sequencer-master.scala 154:24]
  wire  _GEN_9081 = _T_490 ? _GEN_9073 : _GEN_8833; // @[sequencer-master.scala 154:24]
  wire  _GEN_9082 = _T_490 ? _GEN_9074 : _GEN_8834; // @[sequencer-master.scala 154:24]
  wire  _GEN_9083 = _T_490 ? _GEN_9075 : _GEN_8835; // @[sequencer-master.scala 154:24]
  wire  _GEN_9084 = _T_490 ? _GEN_9076 : _GEN_8836; // @[sequencer-master.scala 154:24]
  wire  _GEN_9085 = _T_490 ? _GEN_9077 : _GEN_8837; // @[sequencer-master.scala 154:24]
  wire  _GEN_9086 = _T_490 ? _GEN_9078 : _GEN_8838; // @[sequencer-master.scala 154:24]
  wire  _GEN_9087 = _T_490 ? _GEN_9079 : _GEN_8839; // @[sequencer-master.scala 154:24]
  wire  _GEN_9088 = _GEN_32729 | _GEN_8848; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9089 = _GEN_32730 | _GEN_8849; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9090 = _GEN_32731 | _GEN_8850; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9091 = _GEN_32732 | _GEN_8851; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9092 = _GEN_32733 | _GEN_8852; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9093 = _GEN_32734 | _GEN_8853; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9094 = _GEN_32735 | _GEN_8854; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9095 = _GEN_32736 | _GEN_8855; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9096 = _T_512 ? _GEN_9088 : _GEN_8848; // @[sequencer-master.scala 154:24]
  wire  _GEN_9097 = _T_512 ? _GEN_9089 : _GEN_8849; // @[sequencer-master.scala 154:24]
  wire  _GEN_9098 = _T_512 ? _GEN_9090 : _GEN_8850; // @[sequencer-master.scala 154:24]
  wire  _GEN_9099 = _T_512 ? _GEN_9091 : _GEN_8851; // @[sequencer-master.scala 154:24]
  wire  _GEN_9100 = _T_512 ? _GEN_9092 : _GEN_8852; // @[sequencer-master.scala 154:24]
  wire  _GEN_9101 = _T_512 ? _GEN_9093 : _GEN_8853; // @[sequencer-master.scala 154:24]
  wire  _GEN_9102 = _T_512 ? _GEN_9094 : _GEN_8854; // @[sequencer-master.scala 154:24]
  wire  _GEN_9103 = _T_512 ? _GEN_9095 : _GEN_8855; // @[sequencer-master.scala 154:24]
  wire  _GEN_9104 = _GEN_32729 | _GEN_8864; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9105 = _GEN_32730 | _GEN_8865; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9106 = _GEN_32731 | _GEN_8866; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9107 = _GEN_32732 | _GEN_8867; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9108 = _GEN_32733 | _GEN_8868; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9109 = _GEN_32734 | _GEN_8869; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9110 = _GEN_32735 | _GEN_8870; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9111 = _GEN_32736 | _GEN_8871; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9112 = _T_534 ? _GEN_9104 : _GEN_8864; // @[sequencer-master.scala 154:24]
  wire  _GEN_9113 = _T_534 ? _GEN_9105 : _GEN_8865; // @[sequencer-master.scala 154:24]
  wire  _GEN_9114 = _T_534 ? _GEN_9106 : _GEN_8866; // @[sequencer-master.scala 154:24]
  wire  _GEN_9115 = _T_534 ? _GEN_9107 : _GEN_8867; // @[sequencer-master.scala 154:24]
  wire  _GEN_9116 = _T_534 ? _GEN_9108 : _GEN_8868; // @[sequencer-master.scala 154:24]
  wire  _GEN_9117 = _T_534 ? _GEN_9109 : _GEN_8869; // @[sequencer-master.scala 154:24]
  wire  _GEN_9118 = _T_534 ? _GEN_9110 : _GEN_8870; // @[sequencer-master.scala 154:24]
  wire  _GEN_9119 = _T_534 ? _GEN_9111 : _GEN_8871; // @[sequencer-master.scala 154:24]
  wire  _GEN_9128 = 3'h0 == tail ? io_op_bits_base_vs3_valid : _GEN_8168; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9129 = 3'h1 == tail ? io_op_bits_base_vs3_valid : _GEN_8169; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9130 = 3'h2 == tail ? io_op_bits_base_vs3_valid : _GEN_8170; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9131 = 3'h3 == tail ? io_op_bits_base_vs3_valid : _GEN_8171; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9132 = 3'h4 == tail ? io_op_bits_base_vs3_valid : _GEN_8172; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9133 = 3'h5 == tail ? io_op_bits_base_vs3_valid : _GEN_8173; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9134 = 3'h6 == tail ? io_op_bits_base_vs3_valid : _GEN_8174; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_9135 = 3'h7 == tail ? io_op_bits_base_vs3_valid : _GEN_8175; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_9160 = 3'h0 == tail ? io_op_bits_reg_vs3_id : _GEN_3738; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9161 = 3'h1 == tail ? io_op_bits_reg_vs3_id : _GEN_3739; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9162 = 3'h2 == tail ? io_op_bits_reg_vs3_id : _GEN_3740; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9163 = 3'h3 == tail ? io_op_bits_reg_vs3_id : _GEN_3741; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9164 = 3'h4 == tail ? io_op_bits_reg_vs3_id : _GEN_3742; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9165 = 3'h5 == tail ? io_op_bits_reg_vs3_id : _GEN_3743; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9166 = 3'h6 == tail ? io_op_bits_reg_vs3_id : _GEN_3744; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_9167 = 3'h7 == tail ? io_op_bits_reg_vs3_id : _GEN_3745; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_9168 = 3'h0 == tail ? io_op_bits_sreg_ss3 : _GEN_3746; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9169 = 3'h1 == tail ? io_op_bits_sreg_ss3 : _GEN_3747; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9170 = 3'h2 == tail ? io_op_bits_sreg_ss3 : _GEN_3748; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9171 = 3'h3 == tail ? io_op_bits_sreg_ss3 : _GEN_3749; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9172 = 3'h4 == tail ? io_op_bits_sreg_ss3 : _GEN_3750; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9173 = 3'h5 == tail ? io_op_bits_sreg_ss3 : _GEN_3751; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9174 = 3'h6 == tail ? io_op_bits_sreg_ss3 : _GEN_3752; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_9175 = 3'h7 == tail ? io_op_bits_sreg_ss3 : _GEN_3753; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire  _GEN_9192 = io_op_bits_base_vs3_valid ? _GEN_9128 : _GEN_8168; // @[sequencer-master.scala 328:47]
  wire  _GEN_9193 = io_op_bits_base_vs3_valid ? _GEN_9129 : _GEN_8169; // @[sequencer-master.scala 328:47]
  wire  _GEN_9194 = io_op_bits_base_vs3_valid ? _GEN_9130 : _GEN_8170; // @[sequencer-master.scala 328:47]
  wire  _GEN_9195 = io_op_bits_base_vs3_valid ? _GEN_9131 : _GEN_8171; // @[sequencer-master.scala 328:47]
  wire  _GEN_9196 = io_op_bits_base_vs3_valid ? _GEN_9132 : _GEN_8172; // @[sequencer-master.scala 328:47]
  wire  _GEN_9197 = io_op_bits_base_vs3_valid ? _GEN_9133 : _GEN_8173; // @[sequencer-master.scala 328:47]
  wire  _GEN_9198 = io_op_bits_base_vs3_valid ? _GEN_9134 : _GEN_8174; // @[sequencer-master.scala 328:47]
  wire  _GEN_9199 = io_op_bits_base_vs3_valid ? _GEN_9135 : _GEN_8175; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9224 = io_op_bits_base_vs3_valid ? _GEN_9160 : _GEN_3738; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9225 = io_op_bits_base_vs3_valid ? _GEN_9161 : _GEN_3739; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9226 = io_op_bits_base_vs3_valid ? _GEN_9162 : _GEN_3740; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9227 = io_op_bits_base_vs3_valid ? _GEN_9163 : _GEN_3741; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9228 = io_op_bits_base_vs3_valid ? _GEN_9164 : _GEN_3742; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9229 = io_op_bits_base_vs3_valid ? _GEN_9165 : _GEN_3743; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9230 = io_op_bits_base_vs3_valid ? _GEN_9166 : _GEN_3744; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_9231 = io_op_bits_base_vs3_valid ? _GEN_9167 : _GEN_3745; // @[sequencer-master.scala 328:47]
  wire  _GEN_9240 = _GEN_32729 | _GEN_9000; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9241 = _GEN_32730 | _GEN_9001; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9242 = _GEN_32731 | _GEN_9002; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9243 = _GEN_32732 | _GEN_9003; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9244 = _GEN_32733 | _GEN_9004; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9245 = _GEN_32734 | _GEN_9005; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9246 = _GEN_32735 | _GEN_9006; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9247 = _GEN_32736 | _GEN_9007; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9248 = _T_557 ? _GEN_9240 : _GEN_9000; // @[sequencer-master.scala 154:24]
  wire  _GEN_9249 = _T_557 ? _GEN_9241 : _GEN_9001; // @[sequencer-master.scala 154:24]
  wire  _GEN_9250 = _T_557 ? _GEN_9242 : _GEN_9002; // @[sequencer-master.scala 154:24]
  wire  _GEN_9251 = _T_557 ? _GEN_9243 : _GEN_9003; // @[sequencer-master.scala 154:24]
  wire  _GEN_9252 = _T_557 ? _GEN_9244 : _GEN_9004; // @[sequencer-master.scala 154:24]
  wire  _GEN_9253 = _T_557 ? _GEN_9245 : _GEN_9005; // @[sequencer-master.scala 154:24]
  wire  _GEN_9254 = _T_557 ? _GEN_9246 : _GEN_9006; // @[sequencer-master.scala 154:24]
  wire  _GEN_9255 = _T_557 ? _GEN_9247 : _GEN_9007; // @[sequencer-master.scala 154:24]
  wire  _GEN_9256 = _GEN_32729 | _GEN_9016; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9257 = _GEN_32730 | _GEN_9017; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9258 = _GEN_32731 | _GEN_9018; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9259 = _GEN_32732 | _GEN_9019; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9260 = _GEN_32733 | _GEN_9020; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9261 = _GEN_32734 | _GEN_9021; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9262 = _GEN_32735 | _GEN_9022; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9263 = _GEN_32736 | _GEN_9023; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9264 = _T_579 ? _GEN_9256 : _GEN_9016; // @[sequencer-master.scala 154:24]
  wire  _GEN_9265 = _T_579 ? _GEN_9257 : _GEN_9017; // @[sequencer-master.scala 154:24]
  wire  _GEN_9266 = _T_579 ? _GEN_9258 : _GEN_9018; // @[sequencer-master.scala 154:24]
  wire  _GEN_9267 = _T_579 ? _GEN_9259 : _GEN_9019; // @[sequencer-master.scala 154:24]
  wire  _GEN_9268 = _T_579 ? _GEN_9260 : _GEN_9020; // @[sequencer-master.scala 154:24]
  wire  _GEN_9269 = _T_579 ? _GEN_9261 : _GEN_9021; // @[sequencer-master.scala 154:24]
  wire  _GEN_9270 = _T_579 ? _GEN_9262 : _GEN_9022; // @[sequencer-master.scala 154:24]
  wire  _GEN_9271 = _T_579 ? _GEN_9263 : _GEN_9023; // @[sequencer-master.scala 154:24]
  wire  _GEN_9272 = _GEN_32729 | _GEN_9032; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9273 = _GEN_32730 | _GEN_9033; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9274 = _GEN_32731 | _GEN_9034; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9275 = _GEN_32732 | _GEN_9035; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9276 = _GEN_32733 | _GEN_9036; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9277 = _GEN_32734 | _GEN_9037; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9278 = _GEN_32735 | _GEN_9038; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9279 = _GEN_32736 | _GEN_9039; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9280 = _T_601 ? _GEN_9272 : _GEN_9032; // @[sequencer-master.scala 154:24]
  wire  _GEN_9281 = _T_601 ? _GEN_9273 : _GEN_9033; // @[sequencer-master.scala 154:24]
  wire  _GEN_9282 = _T_601 ? _GEN_9274 : _GEN_9034; // @[sequencer-master.scala 154:24]
  wire  _GEN_9283 = _T_601 ? _GEN_9275 : _GEN_9035; // @[sequencer-master.scala 154:24]
  wire  _GEN_9284 = _T_601 ? _GEN_9276 : _GEN_9036; // @[sequencer-master.scala 154:24]
  wire  _GEN_9285 = _T_601 ? _GEN_9277 : _GEN_9037; // @[sequencer-master.scala 154:24]
  wire  _GEN_9286 = _T_601 ? _GEN_9278 : _GEN_9038; // @[sequencer-master.scala 154:24]
  wire  _GEN_9287 = _T_601 ? _GEN_9279 : _GEN_9039; // @[sequencer-master.scala 154:24]
  wire  _GEN_9288 = _GEN_32729 | _GEN_9048; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9289 = _GEN_32730 | _GEN_9049; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9290 = _GEN_32731 | _GEN_9050; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9291 = _GEN_32732 | _GEN_9051; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9292 = _GEN_32733 | _GEN_9052; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9293 = _GEN_32734 | _GEN_9053; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9294 = _GEN_32735 | _GEN_9054; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9295 = _GEN_32736 | _GEN_9055; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9296 = _T_623 ? _GEN_9288 : _GEN_9048; // @[sequencer-master.scala 154:24]
  wire  _GEN_9297 = _T_623 ? _GEN_9289 : _GEN_9049; // @[sequencer-master.scala 154:24]
  wire  _GEN_9298 = _T_623 ? _GEN_9290 : _GEN_9050; // @[sequencer-master.scala 154:24]
  wire  _GEN_9299 = _T_623 ? _GEN_9291 : _GEN_9051; // @[sequencer-master.scala 154:24]
  wire  _GEN_9300 = _T_623 ? _GEN_9292 : _GEN_9052; // @[sequencer-master.scala 154:24]
  wire  _GEN_9301 = _T_623 ? _GEN_9293 : _GEN_9053; // @[sequencer-master.scala 154:24]
  wire  _GEN_9302 = _T_623 ? _GEN_9294 : _GEN_9054; // @[sequencer-master.scala 154:24]
  wire  _GEN_9303 = _T_623 ? _GEN_9295 : _GEN_9055; // @[sequencer-master.scala 154:24]
  wire  _GEN_9304 = _GEN_32729 | _GEN_9064; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9305 = _GEN_32730 | _GEN_9065; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9306 = _GEN_32731 | _GEN_9066; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9307 = _GEN_32732 | _GEN_9067; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9308 = _GEN_32733 | _GEN_9068; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9309 = _GEN_32734 | _GEN_9069; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9310 = _GEN_32735 | _GEN_9070; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9311 = _GEN_32736 | _GEN_9071; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9312 = _T_645 ? _GEN_9304 : _GEN_9064; // @[sequencer-master.scala 154:24]
  wire  _GEN_9313 = _T_645 ? _GEN_9305 : _GEN_9065; // @[sequencer-master.scala 154:24]
  wire  _GEN_9314 = _T_645 ? _GEN_9306 : _GEN_9066; // @[sequencer-master.scala 154:24]
  wire  _GEN_9315 = _T_645 ? _GEN_9307 : _GEN_9067; // @[sequencer-master.scala 154:24]
  wire  _GEN_9316 = _T_645 ? _GEN_9308 : _GEN_9068; // @[sequencer-master.scala 154:24]
  wire  _GEN_9317 = _T_645 ? _GEN_9309 : _GEN_9069; // @[sequencer-master.scala 154:24]
  wire  _GEN_9318 = _T_645 ? _GEN_9310 : _GEN_9070; // @[sequencer-master.scala 154:24]
  wire  _GEN_9319 = _T_645 ? _GEN_9311 : _GEN_9071; // @[sequencer-master.scala 154:24]
  wire  _GEN_9320 = _GEN_32729 | _GEN_9080; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9321 = _GEN_32730 | _GEN_9081; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9322 = _GEN_32731 | _GEN_9082; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9323 = _GEN_32732 | _GEN_9083; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9324 = _GEN_32733 | _GEN_9084; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9325 = _GEN_32734 | _GEN_9085; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9326 = _GEN_32735 | _GEN_9086; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9327 = _GEN_32736 | _GEN_9087; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9328 = _T_667 ? _GEN_9320 : _GEN_9080; // @[sequencer-master.scala 154:24]
  wire  _GEN_9329 = _T_667 ? _GEN_9321 : _GEN_9081; // @[sequencer-master.scala 154:24]
  wire  _GEN_9330 = _T_667 ? _GEN_9322 : _GEN_9082; // @[sequencer-master.scala 154:24]
  wire  _GEN_9331 = _T_667 ? _GEN_9323 : _GEN_9083; // @[sequencer-master.scala 154:24]
  wire  _GEN_9332 = _T_667 ? _GEN_9324 : _GEN_9084; // @[sequencer-master.scala 154:24]
  wire  _GEN_9333 = _T_667 ? _GEN_9325 : _GEN_9085; // @[sequencer-master.scala 154:24]
  wire  _GEN_9334 = _T_667 ? _GEN_9326 : _GEN_9086; // @[sequencer-master.scala 154:24]
  wire  _GEN_9335 = _T_667 ? _GEN_9327 : _GEN_9087; // @[sequencer-master.scala 154:24]
  wire  _GEN_9336 = _GEN_32729 | _GEN_9096; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9337 = _GEN_32730 | _GEN_9097; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9338 = _GEN_32731 | _GEN_9098; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9339 = _GEN_32732 | _GEN_9099; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9340 = _GEN_32733 | _GEN_9100; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9341 = _GEN_32734 | _GEN_9101; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9342 = _GEN_32735 | _GEN_9102; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9343 = _GEN_32736 | _GEN_9103; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9344 = _T_689 ? _GEN_9336 : _GEN_9096; // @[sequencer-master.scala 154:24]
  wire  _GEN_9345 = _T_689 ? _GEN_9337 : _GEN_9097; // @[sequencer-master.scala 154:24]
  wire  _GEN_9346 = _T_689 ? _GEN_9338 : _GEN_9098; // @[sequencer-master.scala 154:24]
  wire  _GEN_9347 = _T_689 ? _GEN_9339 : _GEN_9099; // @[sequencer-master.scala 154:24]
  wire  _GEN_9348 = _T_689 ? _GEN_9340 : _GEN_9100; // @[sequencer-master.scala 154:24]
  wire  _GEN_9349 = _T_689 ? _GEN_9341 : _GEN_9101; // @[sequencer-master.scala 154:24]
  wire  _GEN_9350 = _T_689 ? _GEN_9342 : _GEN_9102; // @[sequencer-master.scala 154:24]
  wire  _GEN_9351 = _T_689 ? _GEN_9343 : _GEN_9103; // @[sequencer-master.scala 154:24]
  wire  _GEN_9352 = _GEN_32729 | _GEN_9112; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9353 = _GEN_32730 | _GEN_9113; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9354 = _GEN_32731 | _GEN_9114; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9355 = _GEN_32732 | _GEN_9115; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9356 = _GEN_32733 | _GEN_9116; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9357 = _GEN_32734 | _GEN_9117; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9358 = _GEN_32735 | _GEN_9118; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9359 = _GEN_32736 | _GEN_9119; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_9360 = _T_711 ? _GEN_9352 : _GEN_9112; // @[sequencer-master.scala 154:24]
  wire  _GEN_9361 = _T_711 ? _GEN_9353 : _GEN_9113; // @[sequencer-master.scala 154:24]
  wire  _GEN_9362 = _T_711 ? _GEN_9354 : _GEN_9114; // @[sequencer-master.scala 154:24]
  wire  _GEN_9363 = _T_711 ? _GEN_9355 : _GEN_9115; // @[sequencer-master.scala 154:24]
  wire  _GEN_9364 = _T_711 ? _GEN_9356 : _GEN_9116; // @[sequencer-master.scala 154:24]
  wire  _GEN_9365 = _T_711 ? _GEN_9357 : _GEN_9117; // @[sequencer-master.scala 154:24]
  wire  _GEN_9366 = _T_711 ? _GEN_9358 : _GEN_9118; // @[sequencer-master.scala 154:24]
  wire  _GEN_9367 = _T_711 ? _GEN_9359 : _GEN_9119; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_9368 = 3'h0 == tail ? io_op_bits_base_vd_id : _GEN_8086; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9369 = 3'h1 == tail ? io_op_bits_base_vd_id : _GEN_8087; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9370 = 3'h2 == tail ? io_op_bits_base_vd_id : _GEN_8088; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9371 = 3'h3 == tail ? io_op_bits_base_vd_id : _GEN_8089; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9372 = 3'h4 == tail ? io_op_bits_base_vd_id : _GEN_8090; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9373 = 3'h5 == tail ? io_op_bits_base_vd_id : _GEN_8091; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9374 = 3'h6 == tail ? io_op_bits_base_vd_id : _GEN_8092; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9375 = 3'h7 == tail ? io_op_bits_base_vd_id : _GEN_8093; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9376 = 3'h0 == tail ? io_op_bits_base_vd_valid : _GEN_8176; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9377 = 3'h1 == tail ? io_op_bits_base_vd_valid : _GEN_8177; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9378 = 3'h2 == tail ? io_op_bits_base_vd_valid : _GEN_8178; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9379 = 3'h3 == tail ? io_op_bits_base_vd_valid : _GEN_8179; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9380 = 3'h4 == tail ? io_op_bits_base_vd_valid : _GEN_8180; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9381 = 3'h5 == tail ? io_op_bits_base_vd_valid : _GEN_8181; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9382 = 3'h6 == tail ? io_op_bits_base_vd_valid : _GEN_8182; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9383 = 3'h7 == tail ? io_op_bits_base_vd_valid : _GEN_8183; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9384 = 3'h0 == tail ? io_op_bits_base_vd_scalar : _GEN_8094; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9385 = 3'h1 == tail ? io_op_bits_base_vd_scalar : _GEN_8095; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9386 = 3'h2 == tail ? io_op_bits_base_vd_scalar : _GEN_8096; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9387 = 3'h3 == tail ? io_op_bits_base_vd_scalar : _GEN_8097; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9388 = 3'h4 == tail ? io_op_bits_base_vd_scalar : _GEN_8098; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9389 = 3'h5 == tail ? io_op_bits_base_vd_scalar : _GEN_8099; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9390 = 3'h6 == tail ? io_op_bits_base_vd_scalar : _GEN_8100; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9391 = 3'h7 == tail ? io_op_bits_base_vd_scalar : _GEN_8101; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9392 = 3'h0 == tail ? io_op_bits_base_vd_pred : _GEN_8102; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9393 = 3'h1 == tail ? io_op_bits_base_vd_pred : _GEN_8103; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9394 = 3'h2 == tail ? io_op_bits_base_vd_pred : _GEN_8104; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9395 = 3'h3 == tail ? io_op_bits_base_vd_pred : _GEN_8105; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9396 = 3'h4 == tail ? io_op_bits_base_vd_pred : _GEN_8106; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9397 = 3'h5 == tail ? io_op_bits_base_vd_pred : _GEN_8107; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9398 = 3'h6 == tail ? io_op_bits_base_vd_pred : _GEN_8108; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_9399 = 3'h7 == tail ? io_op_bits_base_vd_pred : _GEN_8109; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9400 = 3'h0 == tail ? io_op_bits_base_vd_prec : _GEN_8110; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9401 = 3'h1 == tail ? io_op_bits_base_vd_prec : _GEN_8111; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9402 = 3'h2 == tail ? io_op_bits_base_vd_prec : _GEN_8112; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9403 = 3'h3 == tail ? io_op_bits_base_vd_prec : _GEN_8113; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9404 = 3'h4 == tail ? io_op_bits_base_vd_prec : _GEN_8114; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9405 = 3'h5 == tail ? io_op_bits_base_vd_prec : _GEN_8115; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9406 = 3'h6 == tail ? io_op_bits_base_vd_prec : _GEN_8116; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_9407 = 3'h7 == tail ? io_op_bits_base_vd_prec : _GEN_8117; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_9408 = 3'h0 == tail ? io_op_bits_reg_vd_id : _GEN_8118; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9409 = 3'h1 == tail ? io_op_bits_reg_vd_id : _GEN_8119; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9410 = 3'h2 == tail ? io_op_bits_reg_vd_id : _GEN_8120; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9411 = 3'h3 == tail ? io_op_bits_reg_vd_id : _GEN_8121; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9412 = 3'h4 == tail ? io_op_bits_reg_vd_id : _GEN_8122; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9413 = 3'h5 == tail ? io_op_bits_reg_vd_id : _GEN_8123; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9414 = 3'h6 == tail ? io_op_bits_reg_vd_id : _GEN_8124; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9415 = 3'h7 == tail ? io_op_bits_reg_vd_id : _GEN_8125; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_9416 = io_op_bits_base_vd_valid ? _GEN_9368 : _GEN_8086; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9417 = io_op_bits_base_vd_valid ? _GEN_9369 : _GEN_8087; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9418 = io_op_bits_base_vd_valid ? _GEN_9370 : _GEN_8088; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9419 = io_op_bits_base_vd_valid ? _GEN_9371 : _GEN_8089; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9420 = io_op_bits_base_vd_valid ? _GEN_9372 : _GEN_8090; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9421 = io_op_bits_base_vd_valid ? _GEN_9373 : _GEN_8091; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9422 = io_op_bits_base_vd_valid ? _GEN_9374 : _GEN_8092; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9423 = io_op_bits_base_vd_valid ? _GEN_9375 : _GEN_8093; // @[sequencer-master.scala 362:41]
  wire  _GEN_9424 = io_op_bits_base_vd_valid ? _GEN_9376 : _GEN_8176; // @[sequencer-master.scala 362:41]
  wire  _GEN_9425 = io_op_bits_base_vd_valid ? _GEN_9377 : _GEN_8177; // @[sequencer-master.scala 362:41]
  wire  _GEN_9426 = io_op_bits_base_vd_valid ? _GEN_9378 : _GEN_8178; // @[sequencer-master.scala 362:41]
  wire  _GEN_9427 = io_op_bits_base_vd_valid ? _GEN_9379 : _GEN_8179; // @[sequencer-master.scala 362:41]
  wire  _GEN_9428 = io_op_bits_base_vd_valid ? _GEN_9380 : _GEN_8180; // @[sequencer-master.scala 362:41]
  wire  _GEN_9429 = io_op_bits_base_vd_valid ? _GEN_9381 : _GEN_8181; // @[sequencer-master.scala 362:41]
  wire  _GEN_9430 = io_op_bits_base_vd_valid ? _GEN_9382 : _GEN_8182; // @[sequencer-master.scala 362:41]
  wire  _GEN_9431 = io_op_bits_base_vd_valid ? _GEN_9383 : _GEN_8183; // @[sequencer-master.scala 362:41]
  wire  _GEN_9432 = io_op_bits_base_vd_valid ? _GEN_9384 : _GEN_8094; // @[sequencer-master.scala 362:41]
  wire  _GEN_9433 = io_op_bits_base_vd_valid ? _GEN_9385 : _GEN_8095; // @[sequencer-master.scala 362:41]
  wire  _GEN_9434 = io_op_bits_base_vd_valid ? _GEN_9386 : _GEN_8096; // @[sequencer-master.scala 362:41]
  wire  _GEN_9435 = io_op_bits_base_vd_valid ? _GEN_9387 : _GEN_8097; // @[sequencer-master.scala 362:41]
  wire  _GEN_9436 = io_op_bits_base_vd_valid ? _GEN_9388 : _GEN_8098; // @[sequencer-master.scala 362:41]
  wire  _GEN_9437 = io_op_bits_base_vd_valid ? _GEN_9389 : _GEN_8099; // @[sequencer-master.scala 362:41]
  wire  _GEN_9438 = io_op_bits_base_vd_valid ? _GEN_9390 : _GEN_8100; // @[sequencer-master.scala 362:41]
  wire  _GEN_9439 = io_op_bits_base_vd_valid ? _GEN_9391 : _GEN_8101; // @[sequencer-master.scala 362:41]
  wire  _GEN_9440 = io_op_bits_base_vd_valid ? _GEN_9392 : _GEN_8102; // @[sequencer-master.scala 362:41]
  wire  _GEN_9441 = io_op_bits_base_vd_valid ? _GEN_9393 : _GEN_8103; // @[sequencer-master.scala 362:41]
  wire  _GEN_9442 = io_op_bits_base_vd_valid ? _GEN_9394 : _GEN_8104; // @[sequencer-master.scala 362:41]
  wire  _GEN_9443 = io_op_bits_base_vd_valid ? _GEN_9395 : _GEN_8105; // @[sequencer-master.scala 362:41]
  wire  _GEN_9444 = io_op_bits_base_vd_valid ? _GEN_9396 : _GEN_8106; // @[sequencer-master.scala 362:41]
  wire  _GEN_9445 = io_op_bits_base_vd_valid ? _GEN_9397 : _GEN_8107; // @[sequencer-master.scala 362:41]
  wire  _GEN_9446 = io_op_bits_base_vd_valid ? _GEN_9398 : _GEN_8108; // @[sequencer-master.scala 362:41]
  wire  _GEN_9447 = io_op_bits_base_vd_valid ? _GEN_9399 : _GEN_8109; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9448 = io_op_bits_base_vd_valid ? _GEN_9400 : _GEN_8110; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9449 = io_op_bits_base_vd_valid ? _GEN_9401 : _GEN_8111; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9450 = io_op_bits_base_vd_valid ? _GEN_9402 : _GEN_8112; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9451 = io_op_bits_base_vd_valid ? _GEN_9403 : _GEN_8113; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9452 = io_op_bits_base_vd_valid ? _GEN_9404 : _GEN_8114; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9453 = io_op_bits_base_vd_valid ? _GEN_9405 : _GEN_8115; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9454 = io_op_bits_base_vd_valid ? _GEN_9406 : _GEN_8116; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_9455 = io_op_bits_base_vd_valid ? _GEN_9407 : _GEN_8117; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9456 = io_op_bits_base_vd_valid ? _GEN_9408 : _GEN_8118; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9457 = io_op_bits_base_vd_valid ? _GEN_9409 : _GEN_8119; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9458 = io_op_bits_base_vd_valid ? _GEN_9410 : _GEN_8120; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9459 = io_op_bits_base_vd_valid ? _GEN_9411 : _GEN_8121; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9460 = io_op_bits_base_vd_valid ? _GEN_9412 : _GEN_8122; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9461 = io_op_bits_base_vd_valid ? _GEN_9413 : _GEN_8123; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9462 = io_op_bits_base_vd_valid ? _GEN_9414 : _GEN_8124; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_9463 = io_op_bits_base_vd_valid ? _GEN_9415 : _GEN_8125; // @[sequencer-master.scala 362:41]
  wire  _GEN_9464 = _GEN_32729 | _GEN_8200; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9465 = _GEN_32730 | _GEN_8201; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9466 = _GEN_32731 | _GEN_8202; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9467 = _GEN_32732 | _GEN_8203; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9468 = _GEN_32733 | _GEN_8204; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9469 = _GEN_32734 | _GEN_8205; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9470 = _GEN_32735 | _GEN_8206; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9471 = _GEN_32736 | _GEN_8207; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9472 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9464 : _GEN_8200; // @[sequencer-master.scala 161:86]
  wire  _GEN_9473 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9465 : _GEN_8201; // @[sequencer-master.scala 161:86]
  wire  _GEN_9474 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9466 : _GEN_8202; // @[sequencer-master.scala 161:86]
  wire  _GEN_9475 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9467 : _GEN_8203; // @[sequencer-master.scala 161:86]
  wire  _GEN_9476 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9468 : _GEN_8204; // @[sequencer-master.scala 161:86]
  wire  _GEN_9477 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9469 : _GEN_8205; // @[sequencer-master.scala 161:86]
  wire  _GEN_9478 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9470 : _GEN_8206; // @[sequencer-master.scala 161:86]
  wire  _GEN_9479 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_9471 : _GEN_8207; // @[sequencer-master.scala 161:86]
  wire  _GEN_9480 = _GEN_32729 | _GEN_8224; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9481 = _GEN_32730 | _GEN_8225; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9482 = _GEN_32731 | _GEN_8226; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9483 = _GEN_32732 | _GEN_8227; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9484 = _GEN_32733 | _GEN_8228; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9485 = _GEN_32734 | _GEN_8229; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9486 = _GEN_32735 | _GEN_8230; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9487 = _GEN_32736 | _GEN_8231; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9488 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9480 : _GEN_8224; // @[sequencer-master.scala 161:86]
  wire  _GEN_9489 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9481 : _GEN_8225; // @[sequencer-master.scala 161:86]
  wire  _GEN_9490 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9482 : _GEN_8226; // @[sequencer-master.scala 161:86]
  wire  _GEN_9491 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9483 : _GEN_8227; // @[sequencer-master.scala 161:86]
  wire  _GEN_9492 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9484 : _GEN_8228; // @[sequencer-master.scala 161:86]
  wire  _GEN_9493 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9485 : _GEN_8229; // @[sequencer-master.scala 161:86]
  wire  _GEN_9494 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9486 : _GEN_8230; // @[sequencer-master.scala 161:86]
  wire  _GEN_9495 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_9487 : _GEN_8231; // @[sequencer-master.scala 161:86]
  wire  _GEN_9496 = _GEN_32729 | _GEN_8248; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9497 = _GEN_32730 | _GEN_8249; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9498 = _GEN_32731 | _GEN_8250; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9499 = _GEN_32732 | _GEN_8251; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9500 = _GEN_32733 | _GEN_8252; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9501 = _GEN_32734 | _GEN_8253; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9502 = _GEN_32735 | _GEN_8254; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9503 = _GEN_32736 | _GEN_8255; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9504 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9496 : _GEN_8248; // @[sequencer-master.scala 161:86]
  wire  _GEN_9505 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9497 : _GEN_8249; // @[sequencer-master.scala 161:86]
  wire  _GEN_9506 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9498 : _GEN_8250; // @[sequencer-master.scala 161:86]
  wire  _GEN_9507 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9499 : _GEN_8251; // @[sequencer-master.scala 161:86]
  wire  _GEN_9508 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9500 : _GEN_8252; // @[sequencer-master.scala 161:86]
  wire  _GEN_9509 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9501 : _GEN_8253; // @[sequencer-master.scala 161:86]
  wire  _GEN_9510 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9502 : _GEN_8254; // @[sequencer-master.scala 161:86]
  wire  _GEN_9511 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_9503 : _GEN_8255; // @[sequencer-master.scala 161:86]
  wire  _GEN_9512 = _GEN_32729 | _GEN_8272; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9513 = _GEN_32730 | _GEN_8273; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9514 = _GEN_32731 | _GEN_8274; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9515 = _GEN_32732 | _GEN_8275; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9516 = _GEN_32733 | _GEN_8276; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9517 = _GEN_32734 | _GEN_8277; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9518 = _GEN_32735 | _GEN_8278; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9519 = _GEN_32736 | _GEN_8279; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9520 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9512 : _GEN_8272; // @[sequencer-master.scala 161:86]
  wire  _GEN_9521 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9513 : _GEN_8273; // @[sequencer-master.scala 161:86]
  wire  _GEN_9522 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9514 : _GEN_8274; // @[sequencer-master.scala 161:86]
  wire  _GEN_9523 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9515 : _GEN_8275; // @[sequencer-master.scala 161:86]
  wire  _GEN_9524 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9516 : _GEN_8276; // @[sequencer-master.scala 161:86]
  wire  _GEN_9525 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9517 : _GEN_8277; // @[sequencer-master.scala 161:86]
  wire  _GEN_9526 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9518 : _GEN_8278; // @[sequencer-master.scala 161:86]
  wire  _GEN_9527 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_9519 : _GEN_8279; // @[sequencer-master.scala 161:86]
  wire  _GEN_9528 = _GEN_32729 | _GEN_8296; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9529 = _GEN_32730 | _GEN_8297; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9530 = _GEN_32731 | _GEN_8298; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9531 = _GEN_32732 | _GEN_8299; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9532 = _GEN_32733 | _GEN_8300; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9533 = _GEN_32734 | _GEN_8301; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9534 = _GEN_32735 | _GEN_8302; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9535 = _GEN_32736 | _GEN_8303; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9536 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9528 : _GEN_8296; // @[sequencer-master.scala 161:86]
  wire  _GEN_9537 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9529 : _GEN_8297; // @[sequencer-master.scala 161:86]
  wire  _GEN_9538 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9530 : _GEN_8298; // @[sequencer-master.scala 161:86]
  wire  _GEN_9539 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9531 : _GEN_8299; // @[sequencer-master.scala 161:86]
  wire  _GEN_9540 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9532 : _GEN_8300; // @[sequencer-master.scala 161:86]
  wire  _GEN_9541 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9533 : _GEN_8301; // @[sequencer-master.scala 161:86]
  wire  _GEN_9542 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9534 : _GEN_8302; // @[sequencer-master.scala 161:86]
  wire  _GEN_9543 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_9535 : _GEN_8303; // @[sequencer-master.scala 161:86]
  wire  _GEN_9544 = _GEN_32729 | _GEN_8320; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9545 = _GEN_32730 | _GEN_8321; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9546 = _GEN_32731 | _GEN_8322; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9547 = _GEN_32732 | _GEN_8323; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9548 = _GEN_32733 | _GEN_8324; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9549 = _GEN_32734 | _GEN_8325; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9550 = _GEN_32735 | _GEN_8326; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9551 = _GEN_32736 | _GEN_8327; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9552 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9544 : _GEN_8320; // @[sequencer-master.scala 161:86]
  wire  _GEN_9553 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9545 : _GEN_8321; // @[sequencer-master.scala 161:86]
  wire  _GEN_9554 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9546 : _GEN_8322; // @[sequencer-master.scala 161:86]
  wire  _GEN_9555 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9547 : _GEN_8323; // @[sequencer-master.scala 161:86]
  wire  _GEN_9556 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9548 : _GEN_8324; // @[sequencer-master.scala 161:86]
  wire  _GEN_9557 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9549 : _GEN_8325; // @[sequencer-master.scala 161:86]
  wire  _GEN_9558 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9550 : _GEN_8326; // @[sequencer-master.scala 161:86]
  wire  _GEN_9559 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_9551 : _GEN_8327; // @[sequencer-master.scala 161:86]
  wire  _GEN_9560 = _GEN_32729 | _GEN_8344; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9561 = _GEN_32730 | _GEN_8345; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9562 = _GEN_32731 | _GEN_8346; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9563 = _GEN_32732 | _GEN_8347; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9564 = _GEN_32733 | _GEN_8348; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9565 = _GEN_32734 | _GEN_8349; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9566 = _GEN_32735 | _GEN_8350; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9567 = _GEN_32736 | _GEN_8351; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9568 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9560 : _GEN_8344; // @[sequencer-master.scala 161:86]
  wire  _GEN_9569 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9561 : _GEN_8345; // @[sequencer-master.scala 161:86]
  wire  _GEN_9570 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9562 : _GEN_8346; // @[sequencer-master.scala 161:86]
  wire  _GEN_9571 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9563 : _GEN_8347; // @[sequencer-master.scala 161:86]
  wire  _GEN_9572 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9564 : _GEN_8348; // @[sequencer-master.scala 161:86]
  wire  _GEN_9573 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9565 : _GEN_8349; // @[sequencer-master.scala 161:86]
  wire  _GEN_9574 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9566 : _GEN_8350; // @[sequencer-master.scala 161:86]
  wire  _GEN_9575 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_9567 : _GEN_8351; // @[sequencer-master.scala 161:86]
  wire  _GEN_9576 = _GEN_32729 | _GEN_8368; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9577 = _GEN_32730 | _GEN_8369; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9578 = _GEN_32731 | _GEN_8370; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9579 = _GEN_32732 | _GEN_8371; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9580 = _GEN_32733 | _GEN_8372; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9581 = _GEN_32734 | _GEN_8373; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9582 = _GEN_32735 | _GEN_8374; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9583 = _GEN_32736 | _GEN_8375; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_9584 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9576 : _GEN_8368; // @[sequencer-master.scala 161:86]
  wire  _GEN_9585 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9577 : _GEN_8369; // @[sequencer-master.scala 161:86]
  wire  _GEN_9586 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9578 : _GEN_8370; // @[sequencer-master.scala 161:86]
  wire  _GEN_9587 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9579 : _GEN_8371; // @[sequencer-master.scala 161:86]
  wire  _GEN_9588 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9580 : _GEN_8372; // @[sequencer-master.scala 161:86]
  wire  _GEN_9589 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9581 : _GEN_8373; // @[sequencer-master.scala 161:86]
  wire  _GEN_9590 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9582 : _GEN_8374; // @[sequencer-master.scala 161:86]
  wire  _GEN_9591 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_9583 : _GEN_8375; // @[sequencer-master.scala 161:86]
  wire  _GEN_9592 = _GEN_32729 | _GEN_8208; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9593 = _GEN_32730 | _GEN_8209; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9594 = _GEN_32731 | _GEN_8210; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9595 = _GEN_32732 | _GEN_8211; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9596 = _GEN_32733 | _GEN_8212; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9597 = _GEN_32734 | _GEN_8213; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9598 = _GEN_32735 | _GEN_8214; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9599 = _GEN_32736 | _GEN_8215; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9600 = _T_1442 ? _GEN_9592 : _GEN_8208; // @[sequencer-master.scala 168:32]
  wire  _GEN_9601 = _T_1442 ? _GEN_9593 : _GEN_8209; // @[sequencer-master.scala 168:32]
  wire  _GEN_9602 = _T_1442 ? _GEN_9594 : _GEN_8210; // @[sequencer-master.scala 168:32]
  wire  _GEN_9603 = _T_1442 ? _GEN_9595 : _GEN_8211; // @[sequencer-master.scala 168:32]
  wire  _GEN_9604 = _T_1442 ? _GEN_9596 : _GEN_8212; // @[sequencer-master.scala 168:32]
  wire  _GEN_9605 = _T_1442 ? _GEN_9597 : _GEN_8213; // @[sequencer-master.scala 168:32]
  wire  _GEN_9606 = _T_1442 ? _GEN_9598 : _GEN_8214; // @[sequencer-master.scala 168:32]
  wire  _GEN_9607 = _T_1442 ? _GEN_9599 : _GEN_8215; // @[sequencer-master.scala 168:32]
  wire  _GEN_9608 = _GEN_32729 | _GEN_8232; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9609 = _GEN_32730 | _GEN_8233; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9610 = _GEN_32731 | _GEN_8234; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9611 = _GEN_32732 | _GEN_8235; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9612 = _GEN_32733 | _GEN_8236; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9613 = _GEN_32734 | _GEN_8237; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9614 = _GEN_32735 | _GEN_8238; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9615 = _GEN_32736 | _GEN_8239; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9616 = _T_1464 ? _GEN_9608 : _GEN_8232; // @[sequencer-master.scala 168:32]
  wire  _GEN_9617 = _T_1464 ? _GEN_9609 : _GEN_8233; // @[sequencer-master.scala 168:32]
  wire  _GEN_9618 = _T_1464 ? _GEN_9610 : _GEN_8234; // @[sequencer-master.scala 168:32]
  wire  _GEN_9619 = _T_1464 ? _GEN_9611 : _GEN_8235; // @[sequencer-master.scala 168:32]
  wire  _GEN_9620 = _T_1464 ? _GEN_9612 : _GEN_8236; // @[sequencer-master.scala 168:32]
  wire  _GEN_9621 = _T_1464 ? _GEN_9613 : _GEN_8237; // @[sequencer-master.scala 168:32]
  wire  _GEN_9622 = _T_1464 ? _GEN_9614 : _GEN_8238; // @[sequencer-master.scala 168:32]
  wire  _GEN_9623 = _T_1464 ? _GEN_9615 : _GEN_8239; // @[sequencer-master.scala 168:32]
  wire  _GEN_9624 = _GEN_32729 | _GEN_8256; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9625 = _GEN_32730 | _GEN_8257; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9626 = _GEN_32731 | _GEN_8258; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9627 = _GEN_32732 | _GEN_8259; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9628 = _GEN_32733 | _GEN_8260; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9629 = _GEN_32734 | _GEN_8261; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9630 = _GEN_32735 | _GEN_8262; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9631 = _GEN_32736 | _GEN_8263; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9632 = _T_1486 ? _GEN_9624 : _GEN_8256; // @[sequencer-master.scala 168:32]
  wire  _GEN_9633 = _T_1486 ? _GEN_9625 : _GEN_8257; // @[sequencer-master.scala 168:32]
  wire  _GEN_9634 = _T_1486 ? _GEN_9626 : _GEN_8258; // @[sequencer-master.scala 168:32]
  wire  _GEN_9635 = _T_1486 ? _GEN_9627 : _GEN_8259; // @[sequencer-master.scala 168:32]
  wire  _GEN_9636 = _T_1486 ? _GEN_9628 : _GEN_8260; // @[sequencer-master.scala 168:32]
  wire  _GEN_9637 = _T_1486 ? _GEN_9629 : _GEN_8261; // @[sequencer-master.scala 168:32]
  wire  _GEN_9638 = _T_1486 ? _GEN_9630 : _GEN_8262; // @[sequencer-master.scala 168:32]
  wire  _GEN_9639 = _T_1486 ? _GEN_9631 : _GEN_8263; // @[sequencer-master.scala 168:32]
  wire  _GEN_9640 = _GEN_32729 | _GEN_8280; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9641 = _GEN_32730 | _GEN_8281; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9642 = _GEN_32731 | _GEN_8282; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9643 = _GEN_32732 | _GEN_8283; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9644 = _GEN_32733 | _GEN_8284; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9645 = _GEN_32734 | _GEN_8285; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9646 = _GEN_32735 | _GEN_8286; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9647 = _GEN_32736 | _GEN_8287; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9648 = _T_1508 ? _GEN_9640 : _GEN_8280; // @[sequencer-master.scala 168:32]
  wire  _GEN_9649 = _T_1508 ? _GEN_9641 : _GEN_8281; // @[sequencer-master.scala 168:32]
  wire  _GEN_9650 = _T_1508 ? _GEN_9642 : _GEN_8282; // @[sequencer-master.scala 168:32]
  wire  _GEN_9651 = _T_1508 ? _GEN_9643 : _GEN_8283; // @[sequencer-master.scala 168:32]
  wire  _GEN_9652 = _T_1508 ? _GEN_9644 : _GEN_8284; // @[sequencer-master.scala 168:32]
  wire  _GEN_9653 = _T_1508 ? _GEN_9645 : _GEN_8285; // @[sequencer-master.scala 168:32]
  wire  _GEN_9654 = _T_1508 ? _GEN_9646 : _GEN_8286; // @[sequencer-master.scala 168:32]
  wire  _GEN_9655 = _T_1508 ? _GEN_9647 : _GEN_8287; // @[sequencer-master.scala 168:32]
  wire  _GEN_9656 = _GEN_32729 | _GEN_8304; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9657 = _GEN_32730 | _GEN_8305; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9658 = _GEN_32731 | _GEN_8306; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9659 = _GEN_32732 | _GEN_8307; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9660 = _GEN_32733 | _GEN_8308; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9661 = _GEN_32734 | _GEN_8309; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9662 = _GEN_32735 | _GEN_8310; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9663 = _GEN_32736 | _GEN_8311; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9664 = _T_1530 ? _GEN_9656 : _GEN_8304; // @[sequencer-master.scala 168:32]
  wire  _GEN_9665 = _T_1530 ? _GEN_9657 : _GEN_8305; // @[sequencer-master.scala 168:32]
  wire  _GEN_9666 = _T_1530 ? _GEN_9658 : _GEN_8306; // @[sequencer-master.scala 168:32]
  wire  _GEN_9667 = _T_1530 ? _GEN_9659 : _GEN_8307; // @[sequencer-master.scala 168:32]
  wire  _GEN_9668 = _T_1530 ? _GEN_9660 : _GEN_8308; // @[sequencer-master.scala 168:32]
  wire  _GEN_9669 = _T_1530 ? _GEN_9661 : _GEN_8309; // @[sequencer-master.scala 168:32]
  wire  _GEN_9670 = _T_1530 ? _GEN_9662 : _GEN_8310; // @[sequencer-master.scala 168:32]
  wire  _GEN_9671 = _T_1530 ? _GEN_9663 : _GEN_8311; // @[sequencer-master.scala 168:32]
  wire  _GEN_9672 = _GEN_32729 | _GEN_8328; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9673 = _GEN_32730 | _GEN_8329; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9674 = _GEN_32731 | _GEN_8330; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9675 = _GEN_32732 | _GEN_8331; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9676 = _GEN_32733 | _GEN_8332; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9677 = _GEN_32734 | _GEN_8333; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9678 = _GEN_32735 | _GEN_8334; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9679 = _GEN_32736 | _GEN_8335; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9680 = _T_1552 ? _GEN_9672 : _GEN_8328; // @[sequencer-master.scala 168:32]
  wire  _GEN_9681 = _T_1552 ? _GEN_9673 : _GEN_8329; // @[sequencer-master.scala 168:32]
  wire  _GEN_9682 = _T_1552 ? _GEN_9674 : _GEN_8330; // @[sequencer-master.scala 168:32]
  wire  _GEN_9683 = _T_1552 ? _GEN_9675 : _GEN_8331; // @[sequencer-master.scala 168:32]
  wire  _GEN_9684 = _T_1552 ? _GEN_9676 : _GEN_8332; // @[sequencer-master.scala 168:32]
  wire  _GEN_9685 = _T_1552 ? _GEN_9677 : _GEN_8333; // @[sequencer-master.scala 168:32]
  wire  _GEN_9686 = _T_1552 ? _GEN_9678 : _GEN_8334; // @[sequencer-master.scala 168:32]
  wire  _GEN_9687 = _T_1552 ? _GEN_9679 : _GEN_8335; // @[sequencer-master.scala 168:32]
  wire  _GEN_9688 = _GEN_32729 | _GEN_8352; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9689 = _GEN_32730 | _GEN_8353; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9690 = _GEN_32731 | _GEN_8354; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9691 = _GEN_32732 | _GEN_8355; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9692 = _GEN_32733 | _GEN_8356; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9693 = _GEN_32734 | _GEN_8357; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9694 = _GEN_32735 | _GEN_8358; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9695 = _GEN_32736 | _GEN_8359; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9696 = _T_1574 ? _GEN_9688 : _GEN_8352; // @[sequencer-master.scala 168:32]
  wire  _GEN_9697 = _T_1574 ? _GEN_9689 : _GEN_8353; // @[sequencer-master.scala 168:32]
  wire  _GEN_9698 = _T_1574 ? _GEN_9690 : _GEN_8354; // @[sequencer-master.scala 168:32]
  wire  _GEN_9699 = _T_1574 ? _GEN_9691 : _GEN_8355; // @[sequencer-master.scala 168:32]
  wire  _GEN_9700 = _T_1574 ? _GEN_9692 : _GEN_8356; // @[sequencer-master.scala 168:32]
  wire  _GEN_9701 = _T_1574 ? _GEN_9693 : _GEN_8357; // @[sequencer-master.scala 168:32]
  wire  _GEN_9702 = _T_1574 ? _GEN_9694 : _GEN_8358; // @[sequencer-master.scala 168:32]
  wire  _GEN_9703 = _T_1574 ? _GEN_9695 : _GEN_8359; // @[sequencer-master.scala 168:32]
  wire  _GEN_9704 = _GEN_32729 | _GEN_8376; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9705 = _GEN_32730 | _GEN_8377; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9706 = _GEN_32731 | _GEN_8378; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9707 = _GEN_32732 | _GEN_8379; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9708 = _GEN_32733 | _GEN_8380; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9709 = _GEN_32734 | _GEN_8381; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9710 = _GEN_32735 | _GEN_8382; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9711 = _GEN_32736 | _GEN_8383; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_9712 = _T_1596 ? _GEN_9704 : _GEN_8376; // @[sequencer-master.scala 168:32]
  wire  _GEN_9713 = _T_1596 ? _GEN_9705 : _GEN_8377; // @[sequencer-master.scala 168:32]
  wire  _GEN_9714 = _T_1596 ? _GEN_9706 : _GEN_8378; // @[sequencer-master.scala 168:32]
  wire  _GEN_9715 = _T_1596 ? _GEN_9707 : _GEN_8379; // @[sequencer-master.scala 168:32]
  wire  _GEN_9716 = _T_1596 ? _GEN_9708 : _GEN_8380; // @[sequencer-master.scala 168:32]
  wire  _GEN_9717 = _T_1596 ? _GEN_9709 : _GEN_8381; // @[sequencer-master.scala 168:32]
  wire  _GEN_9718 = _T_1596 ? _GEN_9710 : _GEN_8382; // @[sequencer-master.scala 168:32]
  wire  _GEN_9719 = _T_1596 ? _GEN_9711 : _GEN_8383; // @[sequencer-master.scala 168:32]
  wire [2:0] _T_2007 = _T_1966 ? 3'h5 : 3'h0; // @[Mux.scala 19:72]
  wire [2:0] _T_2008 = _T_1967 ? 3'h4 : 3'h0; // @[Mux.scala 19:72]
  wire [2:0] _T_2009 = _T_1968 ? 3'h4 : 3'h0; // @[Mux.scala 19:72]
  wire [2:0] _T_2010 = _T_2007 | _T_2008; // @[Mux.scala 19:72]
  wire [2:0] _T_2011 = _T_2010 | _T_2009; // @[Mux.scala 19:72]
  wire [1:0] _GEN_9720 = 3'h0 == tail ? _T_1615[1:0] : _GEN_8054; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9721 = 3'h1 == tail ? _T_1615[1:0] : _GEN_8055; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9722 = 3'h2 == tail ? _T_1615[1:0] : _GEN_8056; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9723 = 3'h3 == tail ? _T_1615[1:0] : _GEN_8057; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9724 = 3'h4 == tail ? _T_1615[1:0] : _GEN_8058; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9725 = 3'h5 == tail ? _T_1615[1:0] : _GEN_8059; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9726 = 3'h6 == tail ? _T_1615[1:0] : _GEN_8060; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_9727 = 3'h7 == tail ? _T_1615[1:0] : _GEN_8061; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_9728 = 3'h0 == tail ? 4'h0 : _GEN_8062; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9729 = 3'h1 == tail ? 4'h0 : _GEN_8063; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9730 = 3'h2 == tail ? 4'h0 : _GEN_8064; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9731 = 3'h3 == tail ? 4'h0 : _GEN_8065; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9732 = 3'h4 == tail ? 4'h0 : _GEN_8066; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9733 = 3'h5 == tail ? 4'h0 : _GEN_8067; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9734 = 3'h6 == tail ? 4'h0 : _GEN_8068; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_9735 = 3'h7 == tail ? 4'h0 : _GEN_8069; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_9736 = 3'h0 == tail ? 3'h0 : _GEN_8070; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9737 = 3'h1 == tail ? 3'h0 : _GEN_8071; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9738 = 3'h2 == tail ? 3'h0 : _GEN_8072; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9739 = 3'h3 == tail ? 3'h0 : _GEN_8073; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9740 = 3'h4 == tail ? 3'h0 : _GEN_8074; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9741 = 3'h5 == tail ? 3'h0 : _GEN_8075; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9742 = 3'h6 == tail ? 3'h0 : _GEN_8076; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_9743 = 3'h7 == tail ? 3'h0 : _GEN_8077; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [3:0] _GEN_34697 = {{1'd0}, _T_2011}; // @[sequencer-master.scala 247:56]
  wire [3:0] _T_2016 = _T_1789[3:0] + _GEN_34697; // @[sequencer-master.scala 247:56]
  wire [3:0] _GEN_9744 = 3'h0 == tail ? _T_2016 : _GEN_9728; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9745 = 3'h1 == tail ? _T_2016 : _GEN_9729; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9746 = 3'h2 == tail ? _T_2016 : _GEN_9730; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9747 = 3'h3 == tail ? _T_2016 : _GEN_9731; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9748 = 3'h4 == tail ? _T_2016 : _GEN_9732; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9749 = 3'h5 == tail ? _T_2016 : _GEN_9733; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9750 = 3'h6 == tail ? _T_2016 : _GEN_9734; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9751 = 3'h7 == tail ? _T_2016 : _GEN_9735; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_9752 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9744 : _GEN_9728; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9753 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9745 : _GEN_9729; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9754 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9746 : _GEN_9730; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9755 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9747 : _GEN_9731; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9756 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9748 : _GEN_9732; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9757 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9749 : _GEN_9733; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9758 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9750 : _GEN_9734; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_9759 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_9751 : _GEN_9735; // @[sequencer-master.scala 235:47]
  wire [2:0] _GEN_9760 = 3'h0 == tail ? _T_2016[2:0] : _GEN_9736; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9761 = 3'h1 == tail ? _T_2016[2:0] : _GEN_9737; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9762 = 3'h2 == tail ? _T_2016[2:0] : _GEN_9738; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9763 = 3'h3 == tail ? _T_2016[2:0] : _GEN_9739; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9764 = 3'h4 == tail ? _T_2016[2:0] : _GEN_9740; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9765 = 3'h5 == tail ? _T_2016[2:0] : _GEN_9741; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9766 = 3'h6 == tail ? _T_2016[2:0] : _GEN_9742; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9767 = 3'h7 == tail ? _T_2016[2:0] : _GEN_9743; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_9768 = io_op_bits_base_vd_pred ? _GEN_9760 : _GEN_9736; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9769 = io_op_bits_base_vd_pred ? _GEN_9761 : _GEN_9737; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9770 = io_op_bits_base_vd_pred ? _GEN_9762 : _GEN_9738; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9771 = io_op_bits_base_vd_pred ? _GEN_9763 : _GEN_9739; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9772 = io_op_bits_base_vd_pred ? _GEN_9764 : _GEN_9740; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9773 = io_op_bits_base_vd_pred ? _GEN_9765 : _GEN_9741; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9774 = io_op_bits_base_vd_pred ? _GEN_9766 : _GEN_9742; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_9775 = io_op_bits_base_vd_pred ? _GEN_9767 : _GEN_9743; // @[sequencer-master.scala 236:45]
  wire  _GEN_9776 = io_op_bits_active_vfma ? _GEN_8128 : _GEN_7638; // @[sequencer-master.scala 644:39]
  wire  _GEN_9777 = io_op_bits_active_vfma ? _GEN_8129 : _GEN_7639; // @[sequencer-master.scala 644:39]
  wire  _GEN_9778 = io_op_bits_active_vfma ? _GEN_8130 : _GEN_7640; // @[sequencer-master.scala 644:39]
  wire  _GEN_9779 = io_op_bits_active_vfma ? _GEN_8131 : _GEN_7641; // @[sequencer-master.scala 644:39]
  wire  _GEN_9780 = io_op_bits_active_vfma ? _GEN_8132 : _GEN_7642; // @[sequencer-master.scala 644:39]
  wire  _GEN_9781 = io_op_bits_active_vfma ? _GEN_8133 : _GEN_7643; // @[sequencer-master.scala 644:39]
  wire  _GEN_9782 = io_op_bits_active_vfma ? _GEN_8134 : _GEN_7644; // @[sequencer-master.scala 644:39]
  wire  _GEN_9783 = io_op_bits_active_vfma ? _GEN_8135 : _GEN_7645; // @[sequencer-master.scala 644:39]
  wire  _GEN_9792 = io_op_bits_active_vfma ? _GEN_8464 : _GEN_7654; // @[sequencer-master.scala 644:39]
  wire  _GEN_9793 = io_op_bits_active_vfma ? _GEN_8465 : _GEN_7655; // @[sequencer-master.scala 644:39]
  wire  _GEN_9794 = io_op_bits_active_vfma ? _GEN_8466 : _GEN_7656; // @[sequencer-master.scala 644:39]
  wire  _GEN_9795 = io_op_bits_active_vfma ? _GEN_8467 : _GEN_7657; // @[sequencer-master.scala 644:39]
  wire  _GEN_9796 = io_op_bits_active_vfma ? _GEN_8468 : _GEN_7658; // @[sequencer-master.scala 644:39]
  wire  _GEN_9797 = io_op_bits_active_vfma ? _GEN_8469 : _GEN_7659; // @[sequencer-master.scala 644:39]
  wire  _GEN_9798 = io_op_bits_active_vfma ? _GEN_8470 : _GEN_7660; // @[sequencer-master.scala 644:39]
  wire  _GEN_9799 = io_op_bits_active_vfma ? _GEN_8471 : _GEN_7661; // @[sequencer-master.scala 644:39]
  wire  _GEN_9800 = io_op_bits_active_vfma ? _GEN_8696 : _GEN_7662; // @[sequencer-master.scala 644:39]
  wire  _GEN_9801 = io_op_bits_active_vfma ? _GEN_8697 : _GEN_7663; // @[sequencer-master.scala 644:39]
  wire  _GEN_9802 = io_op_bits_active_vfma ? _GEN_8698 : _GEN_7664; // @[sequencer-master.scala 644:39]
  wire  _GEN_9803 = io_op_bits_active_vfma ? _GEN_8699 : _GEN_7665; // @[sequencer-master.scala 644:39]
  wire  _GEN_9804 = io_op_bits_active_vfma ? _GEN_8700 : _GEN_7666; // @[sequencer-master.scala 644:39]
  wire  _GEN_9805 = io_op_bits_active_vfma ? _GEN_8701 : _GEN_7667; // @[sequencer-master.scala 644:39]
  wire  _GEN_9806 = io_op_bits_active_vfma ? _GEN_8702 : _GEN_7668; // @[sequencer-master.scala 644:39]
  wire  _GEN_9807 = io_op_bits_active_vfma ? _GEN_8703 : _GEN_7669; // @[sequencer-master.scala 644:39]
  wire  _GEN_9808 = io_op_bits_active_vfma ? _GEN_8944 : _GEN_7670; // @[sequencer-master.scala 644:39]
  wire  _GEN_9809 = io_op_bits_active_vfma ? _GEN_8945 : _GEN_7671; // @[sequencer-master.scala 644:39]
  wire  _GEN_9810 = io_op_bits_active_vfma ? _GEN_8946 : _GEN_7672; // @[sequencer-master.scala 644:39]
  wire  _GEN_9811 = io_op_bits_active_vfma ? _GEN_8947 : _GEN_7673; // @[sequencer-master.scala 644:39]
  wire  _GEN_9812 = io_op_bits_active_vfma ? _GEN_8948 : _GEN_7674; // @[sequencer-master.scala 644:39]
  wire  _GEN_9813 = io_op_bits_active_vfma ? _GEN_8949 : _GEN_7675; // @[sequencer-master.scala 644:39]
  wire  _GEN_9814 = io_op_bits_active_vfma ? _GEN_8950 : _GEN_7676; // @[sequencer-master.scala 644:39]
  wire  _GEN_9815 = io_op_bits_active_vfma ? _GEN_8951 : _GEN_7677; // @[sequencer-master.scala 644:39]
  wire  _GEN_9816 = io_op_bits_active_vfma ? _GEN_9192 : _GEN_7678; // @[sequencer-master.scala 644:39]
  wire  _GEN_9817 = io_op_bits_active_vfma ? _GEN_9193 : _GEN_7679; // @[sequencer-master.scala 644:39]
  wire  _GEN_9818 = io_op_bits_active_vfma ? _GEN_9194 : _GEN_7680; // @[sequencer-master.scala 644:39]
  wire  _GEN_9819 = io_op_bits_active_vfma ? _GEN_9195 : _GEN_7681; // @[sequencer-master.scala 644:39]
  wire  _GEN_9820 = io_op_bits_active_vfma ? _GEN_9196 : _GEN_7682; // @[sequencer-master.scala 644:39]
  wire  _GEN_9821 = io_op_bits_active_vfma ? _GEN_9197 : _GEN_7683; // @[sequencer-master.scala 644:39]
  wire  _GEN_9822 = io_op_bits_active_vfma ? _GEN_9198 : _GEN_7684; // @[sequencer-master.scala 644:39]
  wire  _GEN_9823 = io_op_bits_active_vfma ? _GEN_9199 : _GEN_7685; // @[sequencer-master.scala 644:39]
  wire  _GEN_9824 = io_op_bits_active_vfma ? _GEN_9424 : _GEN_7686; // @[sequencer-master.scala 644:39]
  wire  _GEN_9825 = io_op_bits_active_vfma ? _GEN_9425 : _GEN_7687; // @[sequencer-master.scala 644:39]
  wire  _GEN_9826 = io_op_bits_active_vfma ? _GEN_9426 : _GEN_7688; // @[sequencer-master.scala 644:39]
  wire  _GEN_9827 = io_op_bits_active_vfma ? _GEN_9427 : _GEN_7689; // @[sequencer-master.scala 644:39]
  wire  _GEN_9828 = io_op_bits_active_vfma ? _GEN_9428 : _GEN_7690; // @[sequencer-master.scala 644:39]
  wire  _GEN_9829 = io_op_bits_active_vfma ? _GEN_9429 : _GEN_7691; // @[sequencer-master.scala 644:39]
  wire  _GEN_9830 = io_op_bits_active_vfma ? _GEN_9430 : _GEN_7692; // @[sequencer-master.scala 644:39]
  wire  _GEN_9831 = io_op_bits_active_vfma ? _GEN_9431 : _GEN_7693; // @[sequencer-master.scala 644:39]
  wire  _GEN_9832 = io_op_bits_active_vfma ? _GEN_8184 : _GEN_7694; // @[sequencer-master.scala 644:39]
  wire  _GEN_9833 = io_op_bits_active_vfma ? _GEN_8185 : _GEN_7695; // @[sequencer-master.scala 644:39]
  wire  _GEN_9834 = io_op_bits_active_vfma ? _GEN_8186 : _GEN_7696; // @[sequencer-master.scala 644:39]
  wire  _GEN_9835 = io_op_bits_active_vfma ? _GEN_8187 : _GEN_7697; // @[sequencer-master.scala 644:39]
  wire  _GEN_9836 = io_op_bits_active_vfma ? _GEN_8188 : _GEN_7698; // @[sequencer-master.scala 644:39]
  wire  _GEN_9837 = io_op_bits_active_vfma ? _GEN_8189 : _GEN_7699; // @[sequencer-master.scala 644:39]
  wire  _GEN_9838 = io_op_bits_active_vfma ? _GEN_8190 : _GEN_7700; // @[sequencer-master.scala 644:39]
  wire  _GEN_9839 = io_op_bits_active_vfma ? _GEN_8191 : _GEN_7701; // @[sequencer-master.scala 644:39]
  wire  _GEN_9840 = io_op_bits_active_vfma ? _GEN_9248 : _GEN_7702; // @[sequencer-master.scala 644:39]
  wire  _GEN_9841 = io_op_bits_active_vfma ? _GEN_9249 : _GEN_7703; // @[sequencer-master.scala 644:39]
  wire  _GEN_9842 = io_op_bits_active_vfma ? _GEN_9250 : _GEN_7704; // @[sequencer-master.scala 644:39]
  wire  _GEN_9843 = io_op_bits_active_vfma ? _GEN_9251 : _GEN_7705; // @[sequencer-master.scala 644:39]
  wire  _GEN_9844 = io_op_bits_active_vfma ? _GEN_9252 : _GEN_7706; // @[sequencer-master.scala 644:39]
  wire  _GEN_9845 = io_op_bits_active_vfma ? _GEN_9253 : _GEN_7707; // @[sequencer-master.scala 644:39]
  wire  _GEN_9846 = io_op_bits_active_vfma ? _GEN_9254 : _GEN_7708; // @[sequencer-master.scala 644:39]
  wire  _GEN_9847 = io_op_bits_active_vfma ? _GEN_9255 : _GEN_7709; // @[sequencer-master.scala 644:39]
  wire  _GEN_9848 = io_op_bits_active_vfma ? _GEN_9472 : _GEN_7710; // @[sequencer-master.scala 644:39]
  wire  _GEN_9849 = io_op_bits_active_vfma ? _GEN_9473 : _GEN_7711; // @[sequencer-master.scala 644:39]
  wire  _GEN_9850 = io_op_bits_active_vfma ? _GEN_9474 : _GEN_7712; // @[sequencer-master.scala 644:39]
  wire  _GEN_9851 = io_op_bits_active_vfma ? _GEN_9475 : _GEN_7713; // @[sequencer-master.scala 644:39]
  wire  _GEN_9852 = io_op_bits_active_vfma ? _GEN_9476 : _GEN_7714; // @[sequencer-master.scala 644:39]
  wire  _GEN_9853 = io_op_bits_active_vfma ? _GEN_9477 : _GEN_7715; // @[sequencer-master.scala 644:39]
  wire  _GEN_9854 = io_op_bits_active_vfma ? _GEN_9478 : _GEN_7716; // @[sequencer-master.scala 644:39]
  wire  _GEN_9855 = io_op_bits_active_vfma ? _GEN_9479 : _GEN_7717; // @[sequencer-master.scala 644:39]
  wire  _GEN_9856 = io_op_bits_active_vfma ? _GEN_9600 : _GEN_7718; // @[sequencer-master.scala 644:39]
  wire  _GEN_9857 = io_op_bits_active_vfma ? _GEN_9601 : _GEN_7719; // @[sequencer-master.scala 644:39]
  wire  _GEN_9858 = io_op_bits_active_vfma ? _GEN_9602 : _GEN_7720; // @[sequencer-master.scala 644:39]
  wire  _GEN_9859 = io_op_bits_active_vfma ? _GEN_9603 : _GEN_7721; // @[sequencer-master.scala 644:39]
  wire  _GEN_9860 = io_op_bits_active_vfma ? _GEN_9604 : _GEN_7722; // @[sequencer-master.scala 644:39]
  wire  _GEN_9861 = io_op_bits_active_vfma ? _GEN_9605 : _GEN_7723; // @[sequencer-master.scala 644:39]
  wire  _GEN_9862 = io_op_bits_active_vfma ? _GEN_9606 : _GEN_7724; // @[sequencer-master.scala 644:39]
  wire  _GEN_9863 = io_op_bits_active_vfma ? _GEN_9607 : _GEN_7725; // @[sequencer-master.scala 644:39]
  wire  _GEN_9864 = io_op_bits_active_vfma ? _GEN_9264 : _GEN_7726; // @[sequencer-master.scala 644:39]
  wire  _GEN_9865 = io_op_bits_active_vfma ? _GEN_9265 : _GEN_7727; // @[sequencer-master.scala 644:39]
  wire  _GEN_9866 = io_op_bits_active_vfma ? _GEN_9266 : _GEN_7728; // @[sequencer-master.scala 644:39]
  wire  _GEN_9867 = io_op_bits_active_vfma ? _GEN_9267 : _GEN_7729; // @[sequencer-master.scala 644:39]
  wire  _GEN_9868 = io_op_bits_active_vfma ? _GEN_9268 : _GEN_7730; // @[sequencer-master.scala 644:39]
  wire  _GEN_9869 = io_op_bits_active_vfma ? _GEN_9269 : _GEN_7731; // @[sequencer-master.scala 644:39]
  wire  _GEN_9870 = io_op_bits_active_vfma ? _GEN_9270 : _GEN_7732; // @[sequencer-master.scala 644:39]
  wire  _GEN_9871 = io_op_bits_active_vfma ? _GEN_9271 : _GEN_7733; // @[sequencer-master.scala 644:39]
  wire  _GEN_9872 = io_op_bits_active_vfma ? _GEN_9488 : _GEN_7734; // @[sequencer-master.scala 644:39]
  wire  _GEN_9873 = io_op_bits_active_vfma ? _GEN_9489 : _GEN_7735; // @[sequencer-master.scala 644:39]
  wire  _GEN_9874 = io_op_bits_active_vfma ? _GEN_9490 : _GEN_7736; // @[sequencer-master.scala 644:39]
  wire  _GEN_9875 = io_op_bits_active_vfma ? _GEN_9491 : _GEN_7737; // @[sequencer-master.scala 644:39]
  wire  _GEN_9876 = io_op_bits_active_vfma ? _GEN_9492 : _GEN_7738; // @[sequencer-master.scala 644:39]
  wire  _GEN_9877 = io_op_bits_active_vfma ? _GEN_9493 : _GEN_7739; // @[sequencer-master.scala 644:39]
  wire  _GEN_9878 = io_op_bits_active_vfma ? _GEN_9494 : _GEN_7740; // @[sequencer-master.scala 644:39]
  wire  _GEN_9879 = io_op_bits_active_vfma ? _GEN_9495 : _GEN_7741; // @[sequencer-master.scala 644:39]
  wire  _GEN_9880 = io_op_bits_active_vfma ? _GEN_9616 : _GEN_7742; // @[sequencer-master.scala 644:39]
  wire  _GEN_9881 = io_op_bits_active_vfma ? _GEN_9617 : _GEN_7743; // @[sequencer-master.scala 644:39]
  wire  _GEN_9882 = io_op_bits_active_vfma ? _GEN_9618 : _GEN_7744; // @[sequencer-master.scala 644:39]
  wire  _GEN_9883 = io_op_bits_active_vfma ? _GEN_9619 : _GEN_7745; // @[sequencer-master.scala 644:39]
  wire  _GEN_9884 = io_op_bits_active_vfma ? _GEN_9620 : _GEN_7746; // @[sequencer-master.scala 644:39]
  wire  _GEN_9885 = io_op_bits_active_vfma ? _GEN_9621 : _GEN_7747; // @[sequencer-master.scala 644:39]
  wire  _GEN_9886 = io_op_bits_active_vfma ? _GEN_9622 : _GEN_7748; // @[sequencer-master.scala 644:39]
  wire  _GEN_9887 = io_op_bits_active_vfma ? _GEN_9623 : _GEN_7749; // @[sequencer-master.scala 644:39]
  wire  _GEN_9888 = io_op_bits_active_vfma ? _GEN_9280 : _GEN_7750; // @[sequencer-master.scala 644:39]
  wire  _GEN_9889 = io_op_bits_active_vfma ? _GEN_9281 : _GEN_7751; // @[sequencer-master.scala 644:39]
  wire  _GEN_9890 = io_op_bits_active_vfma ? _GEN_9282 : _GEN_7752; // @[sequencer-master.scala 644:39]
  wire  _GEN_9891 = io_op_bits_active_vfma ? _GEN_9283 : _GEN_7753; // @[sequencer-master.scala 644:39]
  wire  _GEN_9892 = io_op_bits_active_vfma ? _GEN_9284 : _GEN_7754; // @[sequencer-master.scala 644:39]
  wire  _GEN_9893 = io_op_bits_active_vfma ? _GEN_9285 : _GEN_7755; // @[sequencer-master.scala 644:39]
  wire  _GEN_9894 = io_op_bits_active_vfma ? _GEN_9286 : _GEN_7756; // @[sequencer-master.scala 644:39]
  wire  _GEN_9895 = io_op_bits_active_vfma ? _GEN_9287 : _GEN_7757; // @[sequencer-master.scala 644:39]
  wire  _GEN_9896 = io_op_bits_active_vfma ? _GEN_9504 : _GEN_7758; // @[sequencer-master.scala 644:39]
  wire  _GEN_9897 = io_op_bits_active_vfma ? _GEN_9505 : _GEN_7759; // @[sequencer-master.scala 644:39]
  wire  _GEN_9898 = io_op_bits_active_vfma ? _GEN_9506 : _GEN_7760; // @[sequencer-master.scala 644:39]
  wire  _GEN_9899 = io_op_bits_active_vfma ? _GEN_9507 : _GEN_7761; // @[sequencer-master.scala 644:39]
  wire  _GEN_9900 = io_op_bits_active_vfma ? _GEN_9508 : _GEN_7762; // @[sequencer-master.scala 644:39]
  wire  _GEN_9901 = io_op_bits_active_vfma ? _GEN_9509 : _GEN_7763; // @[sequencer-master.scala 644:39]
  wire  _GEN_9902 = io_op_bits_active_vfma ? _GEN_9510 : _GEN_7764; // @[sequencer-master.scala 644:39]
  wire  _GEN_9903 = io_op_bits_active_vfma ? _GEN_9511 : _GEN_7765; // @[sequencer-master.scala 644:39]
  wire  _GEN_9904 = io_op_bits_active_vfma ? _GEN_9632 : _GEN_7766; // @[sequencer-master.scala 644:39]
  wire  _GEN_9905 = io_op_bits_active_vfma ? _GEN_9633 : _GEN_7767; // @[sequencer-master.scala 644:39]
  wire  _GEN_9906 = io_op_bits_active_vfma ? _GEN_9634 : _GEN_7768; // @[sequencer-master.scala 644:39]
  wire  _GEN_9907 = io_op_bits_active_vfma ? _GEN_9635 : _GEN_7769; // @[sequencer-master.scala 644:39]
  wire  _GEN_9908 = io_op_bits_active_vfma ? _GEN_9636 : _GEN_7770; // @[sequencer-master.scala 644:39]
  wire  _GEN_9909 = io_op_bits_active_vfma ? _GEN_9637 : _GEN_7771; // @[sequencer-master.scala 644:39]
  wire  _GEN_9910 = io_op_bits_active_vfma ? _GEN_9638 : _GEN_7772; // @[sequencer-master.scala 644:39]
  wire  _GEN_9911 = io_op_bits_active_vfma ? _GEN_9639 : _GEN_7773; // @[sequencer-master.scala 644:39]
  wire  _GEN_9912 = io_op_bits_active_vfma ? _GEN_9296 : _GEN_7774; // @[sequencer-master.scala 644:39]
  wire  _GEN_9913 = io_op_bits_active_vfma ? _GEN_9297 : _GEN_7775; // @[sequencer-master.scala 644:39]
  wire  _GEN_9914 = io_op_bits_active_vfma ? _GEN_9298 : _GEN_7776; // @[sequencer-master.scala 644:39]
  wire  _GEN_9915 = io_op_bits_active_vfma ? _GEN_9299 : _GEN_7777; // @[sequencer-master.scala 644:39]
  wire  _GEN_9916 = io_op_bits_active_vfma ? _GEN_9300 : _GEN_7778; // @[sequencer-master.scala 644:39]
  wire  _GEN_9917 = io_op_bits_active_vfma ? _GEN_9301 : _GEN_7779; // @[sequencer-master.scala 644:39]
  wire  _GEN_9918 = io_op_bits_active_vfma ? _GEN_9302 : _GEN_7780; // @[sequencer-master.scala 644:39]
  wire  _GEN_9919 = io_op_bits_active_vfma ? _GEN_9303 : _GEN_7781; // @[sequencer-master.scala 644:39]
  wire  _GEN_9920 = io_op_bits_active_vfma ? _GEN_9520 : _GEN_7782; // @[sequencer-master.scala 644:39]
  wire  _GEN_9921 = io_op_bits_active_vfma ? _GEN_9521 : _GEN_7783; // @[sequencer-master.scala 644:39]
  wire  _GEN_9922 = io_op_bits_active_vfma ? _GEN_9522 : _GEN_7784; // @[sequencer-master.scala 644:39]
  wire  _GEN_9923 = io_op_bits_active_vfma ? _GEN_9523 : _GEN_7785; // @[sequencer-master.scala 644:39]
  wire  _GEN_9924 = io_op_bits_active_vfma ? _GEN_9524 : _GEN_7786; // @[sequencer-master.scala 644:39]
  wire  _GEN_9925 = io_op_bits_active_vfma ? _GEN_9525 : _GEN_7787; // @[sequencer-master.scala 644:39]
  wire  _GEN_9926 = io_op_bits_active_vfma ? _GEN_9526 : _GEN_7788; // @[sequencer-master.scala 644:39]
  wire  _GEN_9927 = io_op_bits_active_vfma ? _GEN_9527 : _GEN_7789; // @[sequencer-master.scala 644:39]
  wire  _GEN_9928 = io_op_bits_active_vfma ? _GEN_9648 : _GEN_7790; // @[sequencer-master.scala 644:39]
  wire  _GEN_9929 = io_op_bits_active_vfma ? _GEN_9649 : _GEN_7791; // @[sequencer-master.scala 644:39]
  wire  _GEN_9930 = io_op_bits_active_vfma ? _GEN_9650 : _GEN_7792; // @[sequencer-master.scala 644:39]
  wire  _GEN_9931 = io_op_bits_active_vfma ? _GEN_9651 : _GEN_7793; // @[sequencer-master.scala 644:39]
  wire  _GEN_9932 = io_op_bits_active_vfma ? _GEN_9652 : _GEN_7794; // @[sequencer-master.scala 644:39]
  wire  _GEN_9933 = io_op_bits_active_vfma ? _GEN_9653 : _GEN_7795; // @[sequencer-master.scala 644:39]
  wire  _GEN_9934 = io_op_bits_active_vfma ? _GEN_9654 : _GEN_7796; // @[sequencer-master.scala 644:39]
  wire  _GEN_9935 = io_op_bits_active_vfma ? _GEN_9655 : _GEN_7797; // @[sequencer-master.scala 644:39]
  wire  _GEN_9936 = io_op_bits_active_vfma ? _GEN_9312 : _GEN_7798; // @[sequencer-master.scala 644:39]
  wire  _GEN_9937 = io_op_bits_active_vfma ? _GEN_9313 : _GEN_7799; // @[sequencer-master.scala 644:39]
  wire  _GEN_9938 = io_op_bits_active_vfma ? _GEN_9314 : _GEN_7800; // @[sequencer-master.scala 644:39]
  wire  _GEN_9939 = io_op_bits_active_vfma ? _GEN_9315 : _GEN_7801; // @[sequencer-master.scala 644:39]
  wire  _GEN_9940 = io_op_bits_active_vfma ? _GEN_9316 : _GEN_7802; // @[sequencer-master.scala 644:39]
  wire  _GEN_9941 = io_op_bits_active_vfma ? _GEN_9317 : _GEN_7803; // @[sequencer-master.scala 644:39]
  wire  _GEN_9942 = io_op_bits_active_vfma ? _GEN_9318 : _GEN_7804; // @[sequencer-master.scala 644:39]
  wire  _GEN_9943 = io_op_bits_active_vfma ? _GEN_9319 : _GEN_7805; // @[sequencer-master.scala 644:39]
  wire  _GEN_9944 = io_op_bits_active_vfma ? _GEN_9536 : _GEN_7806; // @[sequencer-master.scala 644:39]
  wire  _GEN_9945 = io_op_bits_active_vfma ? _GEN_9537 : _GEN_7807; // @[sequencer-master.scala 644:39]
  wire  _GEN_9946 = io_op_bits_active_vfma ? _GEN_9538 : _GEN_7808; // @[sequencer-master.scala 644:39]
  wire  _GEN_9947 = io_op_bits_active_vfma ? _GEN_9539 : _GEN_7809; // @[sequencer-master.scala 644:39]
  wire  _GEN_9948 = io_op_bits_active_vfma ? _GEN_9540 : _GEN_7810; // @[sequencer-master.scala 644:39]
  wire  _GEN_9949 = io_op_bits_active_vfma ? _GEN_9541 : _GEN_7811; // @[sequencer-master.scala 644:39]
  wire  _GEN_9950 = io_op_bits_active_vfma ? _GEN_9542 : _GEN_7812; // @[sequencer-master.scala 644:39]
  wire  _GEN_9951 = io_op_bits_active_vfma ? _GEN_9543 : _GEN_7813; // @[sequencer-master.scala 644:39]
  wire  _GEN_9952 = io_op_bits_active_vfma ? _GEN_9664 : _GEN_7814; // @[sequencer-master.scala 644:39]
  wire  _GEN_9953 = io_op_bits_active_vfma ? _GEN_9665 : _GEN_7815; // @[sequencer-master.scala 644:39]
  wire  _GEN_9954 = io_op_bits_active_vfma ? _GEN_9666 : _GEN_7816; // @[sequencer-master.scala 644:39]
  wire  _GEN_9955 = io_op_bits_active_vfma ? _GEN_9667 : _GEN_7817; // @[sequencer-master.scala 644:39]
  wire  _GEN_9956 = io_op_bits_active_vfma ? _GEN_9668 : _GEN_7818; // @[sequencer-master.scala 644:39]
  wire  _GEN_9957 = io_op_bits_active_vfma ? _GEN_9669 : _GEN_7819; // @[sequencer-master.scala 644:39]
  wire  _GEN_9958 = io_op_bits_active_vfma ? _GEN_9670 : _GEN_7820; // @[sequencer-master.scala 644:39]
  wire  _GEN_9959 = io_op_bits_active_vfma ? _GEN_9671 : _GEN_7821; // @[sequencer-master.scala 644:39]
  wire  _GEN_9960 = io_op_bits_active_vfma ? _GEN_9328 : _GEN_7822; // @[sequencer-master.scala 644:39]
  wire  _GEN_9961 = io_op_bits_active_vfma ? _GEN_9329 : _GEN_7823; // @[sequencer-master.scala 644:39]
  wire  _GEN_9962 = io_op_bits_active_vfma ? _GEN_9330 : _GEN_7824; // @[sequencer-master.scala 644:39]
  wire  _GEN_9963 = io_op_bits_active_vfma ? _GEN_9331 : _GEN_7825; // @[sequencer-master.scala 644:39]
  wire  _GEN_9964 = io_op_bits_active_vfma ? _GEN_9332 : _GEN_7826; // @[sequencer-master.scala 644:39]
  wire  _GEN_9965 = io_op_bits_active_vfma ? _GEN_9333 : _GEN_7827; // @[sequencer-master.scala 644:39]
  wire  _GEN_9966 = io_op_bits_active_vfma ? _GEN_9334 : _GEN_7828; // @[sequencer-master.scala 644:39]
  wire  _GEN_9967 = io_op_bits_active_vfma ? _GEN_9335 : _GEN_7829; // @[sequencer-master.scala 644:39]
  wire  _GEN_9968 = io_op_bits_active_vfma ? _GEN_9552 : _GEN_7830; // @[sequencer-master.scala 644:39]
  wire  _GEN_9969 = io_op_bits_active_vfma ? _GEN_9553 : _GEN_7831; // @[sequencer-master.scala 644:39]
  wire  _GEN_9970 = io_op_bits_active_vfma ? _GEN_9554 : _GEN_7832; // @[sequencer-master.scala 644:39]
  wire  _GEN_9971 = io_op_bits_active_vfma ? _GEN_9555 : _GEN_7833; // @[sequencer-master.scala 644:39]
  wire  _GEN_9972 = io_op_bits_active_vfma ? _GEN_9556 : _GEN_7834; // @[sequencer-master.scala 644:39]
  wire  _GEN_9973 = io_op_bits_active_vfma ? _GEN_9557 : _GEN_7835; // @[sequencer-master.scala 644:39]
  wire  _GEN_9974 = io_op_bits_active_vfma ? _GEN_9558 : _GEN_7836; // @[sequencer-master.scala 644:39]
  wire  _GEN_9975 = io_op_bits_active_vfma ? _GEN_9559 : _GEN_7837; // @[sequencer-master.scala 644:39]
  wire  _GEN_9976 = io_op_bits_active_vfma ? _GEN_9680 : _GEN_7838; // @[sequencer-master.scala 644:39]
  wire  _GEN_9977 = io_op_bits_active_vfma ? _GEN_9681 : _GEN_7839; // @[sequencer-master.scala 644:39]
  wire  _GEN_9978 = io_op_bits_active_vfma ? _GEN_9682 : _GEN_7840; // @[sequencer-master.scala 644:39]
  wire  _GEN_9979 = io_op_bits_active_vfma ? _GEN_9683 : _GEN_7841; // @[sequencer-master.scala 644:39]
  wire  _GEN_9980 = io_op_bits_active_vfma ? _GEN_9684 : _GEN_7842; // @[sequencer-master.scala 644:39]
  wire  _GEN_9981 = io_op_bits_active_vfma ? _GEN_9685 : _GEN_7843; // @[sequencer-master.scala 644:39]
  wire  _GEN_9982 = io_op_bits_active_vfma ? _GEN_9686 : _GEN_7844; // @[sequencer-master.scala 644:39]
  wire  _GEN_9983 = io_op_bits_active_vfma ? _GEN_9687 : _GEN_7845; // @[sequencer-master.scala 644:39]
  wire  _GEN_9984 = io_op_bits_active_vfma ? _GEN_9344 : _GEN_7846; // @[sequencer-master.scala 644:39]
  wire  _GEN_9985 = io_op_bits_active_vfma ? _GEN_9345 : _GEN_7847; // @[sequencer-master.scala 644:39]
  wire  _GEN_9986 = io_op_bits_active_vfma ? _GEN_9346 : _GEN_7848; // @[sequencer-master.scala 644:39]
  wire  _GEN_9987 = io_op_bits_active_vfma ? _GEN_9347 : _GEN_7849; // @[sequencer-master.scala 644:39]
  wire  _GEN_9988 = io_op_bits_active_vfma ? _GEN_9348 : _GEN_7850; // @[sequencer-master.scala 644:39]
  wire  _GEN_9989 = io_op_bits_active_vfma ? _GEN_9349 : _GEN_7851; // @[sequencer-master.scala 644:39]
  wire  _GEN_9990 = io_op_bits_active_vfma ? _GEN_9350 : _GEN_7852; // @[sequencer-master.scala 644:39]
  wire  _GEN_9991 = io_op_bits_active_vfma ? _GEN_9351 : _GEN_7853; // @[sequencer-master.scala 644:39]
  wire  _GEN_9992 = io_op_bits_active_vfma ? _GEN_9568 : _GEN_7854; // @[sequencer-master.scala 644:39]
  wire  _GEN_9993 = io_op_bits_active_vfma ? _GEN_9569 : _GEN_7855; // @[sequencer-master.scala 644:39]
  wire  _GEN_9994 = io_op_bits_active_vfma ? _GEN_9570 : _GEN_7856; // @[sequencer-master.scala 644:39]
  wire  _GEN_9995 = io_op_bits_active_vfma ? _GEN_9571 : _GEN_7857; // @[sequencer-master.scala 644:39]
  wire  _GEN_9996 = io_op_bits_active_vfma ? _GEN_9572 : _GEN_7858; // @[sequencer-master.scala 644:39]
  wire  _GEN_9997 = io_op_bits_active_vfma ? _GEN_9573 : _GEN_7859; // @[sequencer-master.scala 644:39]
  wire  _GEN_9998 = io_op_bits_active_vfma ? _GEN_9574 : _GEN_7860; // @[sequencer-master.scala 644:39]
  wire  _GEN_9999 = io_op_bits_active_vfma ? _GEN_9575 : _GEN_7861; // @[sequencer-master.scala 644:39]
  wire  _GEN_10000 = io_op_bits_active_vfma ? _GEN_9696 : _GEN_7862; // @[sequencer-master.scala 644:39]
  wire  _GEN_10001 = io_op_bits_active_vfma ? _GEN_9697 : _GEN_7863; // @[sequencer-master.scala 644:39]
  wire  _GEN_10002 = io_op_bits_active_vfma ? _GEN_9698 : _GEN_7864; // @[sequencer-master.scala 644:39]
  wire  _GEN_10003 = io_op_bits_active_vfma ? _GEN_9699 : _GEN_7865; // @[sequencer-master.scala 644:39]
  wire  _GEN_10004 = io_op_bits_active_vfma ? _GEN_9700 : _GEN_7866; // @[sequencer-master.scala 644:39]
  wire  _GEN_10005 = io_op_bits_active_vfma ? _GEN_9701 : _GEN_7867; // @[sequencer-master.scala 644:39]
  wire  _GEN_10006 = io_op_bits_active_vfma ? _GEN_9702 : _GEN_7868; // @[sequencer-master.scala 644:39]
  wire  _GEN_10007 = io_op_bits_active_vfma ? _GEN_9703 : _GEN_7869; // @[sequencer-master.scala 644:39]
  wire  _GEN_10008 = io_op_bits_active_vfma ? _GEN_9360 : _GEN_7870; // @[sequencer-master.scala 644:39]
  wire  _GEN_10009 = io_op_bits_active_vfma ? _GEN_9361 : _GEN_7871; // @[sequencer-master.scala 644:39]
  wire  _GEN_10010 = io_op_bits_active_vfma ? _GEN_9362 : _GEN_7872; // @[sequencer-master.scala 644:39]
  wire  _GEN_10011 = io_op_bits_active_vfma ? _GEN_9363 : _GEN_7873; // @[sequencer-master.scala 644:39]
  wire  _GEN_10012 = io_op_bits_active_vfma ? _GEN_9364 : _GEN_7874; // @[sequencer-master.scala 644:39]
  wire  _GEN_10013 = io_op_bits_active_vfma ? _GEN_9365 : _GEN_7875; // @[sequencer-master.scala 644:39]
  wire  _GEN_10014 = io_op_bits_active_vfma ? _GEN_9366 : _GEN_7876; // @[sequencer-master.scala 644:39]
  wire  _GEN_10015 = io_op_bits_active_vfma ? _GEN_9367 : _GEN_7877; // @[sequencer-master.scala 644:39]
  wire  _GEN_10016 = io_op_bits_active_vfma ? _GEN_9584 : _GEN_7878; // @[sequencer-master.scala 644:39]
  wire  _GEN_10017 = io_op_bits_active_vfma ? _GEN_9585 : _GEN_7879; // @[sequencer-master.scala 644:39]
  wire  _GEN_10018 = io_op_bits_active_vfma ? _GEN_9586 : _GEN_7880; // @[sequencer-master.scala 644:39]
  wire  _GEN_10019 = io_op_bits_active_vfma ? _GEN_9587 : _GEN_7881; // @[sequencer-master.scala 644:39]
  wire  _GEN_10020 = io_op_bits_active_vfma ? _GEN_9588 : _GEN_7882; // @[sequencer-master.scala 644:39]
  wire  _GEN_10021 = io_op_bits_active_vfma ? _GEN_9589 : _GEN_7883; // @[sequencer-master.scala 644:39]
  wire  _GEN_10022 = io_op_bits_active_vfma ? _GEN_9590 : _GEN_7884; // @[sequencer-master.scala 644:39]
  wire  _GEN_10023 = io_op_bits_active_vfma ? _GEN_9591 : _GEN_7885; // @[sequencer-master.scala 644:39]
  wire  _GEN_10024 = io_op_bits_active_vfma ? _GEN_9712 : _GEN_7886; // @[sequencer-master.scala 644:39]
  wire  _GEN_10025 = io_op_bits_active_vfma ? _GEN_9713 : _GEN_7887; // @[sequencer-master.scala 644:39]
  wire  _GEN_10026 = io_op_bits_active_vfma ? _GEN_9714 : _GEN_7888; // @[sequencer-master.scala 644:39]
  wire  _GEN_10027 = io_op_bits_active_vfma ? _GEN_9715 : _GEN_7889; // @[sequencer-master.scala 644:39]
  wire  _GEN_10028 = io_op_bits_active_vfma ? _GEN_9716 : _GEN_7890; // @[sequencer-master.scala 644:39]
  wire  _GEN_10029 = io_op_bits_active_vfma ? _GEN_9717 : _GEN_7891; // @[sequencer-master.scala 644:39]
  wire  _GEN_10030 = io_op_bits_active_vfma ? _GEN_9718 : _GEN_7892; // @[sequencer-master.scala 644:39]
  wire  _GEN_10031 = io_op_bits_active_vfma ? _GEN_9719 : _GEN_7893; // @[sequencer-master.scala 644:39]
  wire  _GEN_10032 = io_op_bits_active_vfma ? _GEN_8384 : _GEN_7894; // @[sequencer-master.scala 644:39]
  wire  _GEN_10033 = io_op_bits_active_vfma ? _GEN_8385 : _GEN_7895; // @[sequencer-master.scala 644:39]
  wire  _GEN_10034 = io_op_bits_active_vfma ? _GEN_8386 : _GEN_7896; // @[sequencer-master.scala 644:39]
  wire  _GEN_10035 = io_op_bits_active_vfma ? _GEN_8387 : _GEN_7897; // @[sequencer-master.scala 644:39]
  wire  _GEN_10036 = io_op_bits_active_vfma ? _GEN_8388 : _GEN_7898; // @[sequencer-master.scala 644:39]
  wire  _GEN_10037 = io_op_bits_active_vfma ? _GEN_8389 : _GEN_7899; // @[sequencer-master.scala 644:39]
  wire  _GEN_10038 = io_op_bits_active_vfma ? _GEN_8390 : _GEN_7900; // @[sequencer-master.scala 644:39]
  wire  _GEN_10039 = io_op_bits_active_vfma ? _GEN_8391 : _GEN_7901; // @[sequencer-master.scala 644:39]
  wire  _GEN_10048 = io_op_bits_active_vfma ? _GEN_8400 : e_0_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10049 = io_op_bits_active_vfma ? _GEN_8401 : e_1_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10050 = io_op_bits_active_vfma ? _GEN_8402 : e_2_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10051 = io_op_bits_active_vfma ? _GEN_8403 : e_3_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10052 = io_op_bits_active_vfma ? _GEN_8404 : e_4_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10053 = io_op_bits_active_vfma ? _GEN_8405 : e_5_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10054 = io_op_bits_active_vfma ? _GEN_8406 : e_6_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire  _GEN_10055 = io_op_bits_active_vfma ? _GEN_8407 : e_7_active_vfmu; // @[sequencer-master.scala 644:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_10056 = io_op_bits_active_vfma ? _GEN_8408 : _GEN_7918; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10057 = io_op_bits_active_vfma ? _GEN_8409 : _GEN_7919; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10058 = io_op_bits_active_vfma ? _GEN_8410 : _GEN_7920; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10059 = io_op_bits_active_vfma ? _GEN_8411 : _GEN_7921; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10060 = io_op_bits_active_vfma ? _GEN_8412 : _GEN_7922; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10061 = io_op_bits_active_vfma ? _GEN_8413 : _GEN_7923; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10062 = io_op_bits_active_vfma ? _GEN_8414 : _GEN_7924; // @[sequencer-master.scala 644:39]
  wire [9:0] _GEN_10063 = io_op_bits_active_vfma ? _GEN_8415 : _GEN_7925; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10064 = io_op_bits_active_vfma ? _GEN_8456 : _GEN_7926; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10065 = io_op_bits_active_vfma ? _GEN_8457 : _GEN_7927; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10066 = io_op_bits_active_vfma ? _GEN_8458 : _GEN_7928; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10067 = io_op_bits_active_vfma ? _GEN_8459 : _GEN_7929; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10068 = io_op_bits_active_vfma ? _GEN_8460 : _GEN_7930; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10069 = io_op_bits_active_vfma ? _GEN_8461 : _GEN_7931; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10070 = io_op_bits_active_vfma ? _GEN_8462 : _GEN_7932; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10071 = io_op_bits_active_vfma ? _GEN_8463 : _GEN_7933; // @[sequencer-master.scala 644:39]
  wire  _GEN_10072 = io_op_bits_active_vfma ? _GEN_8472 : _GEN_7934; // @[sequencer-master.scala 644:39]
  wire  _GEN_10073 = io_op_bits_active_vfma ? _GEN_8473 : _GEN_7935; // @[sequencer-master.scala 644:39]
  wire  _GEN_10074 = io_op_bits_active_vfma ? _GEN_8474 : _GEN_7936; // @[sequencer-master.scala 644:39]
  wire  _GEN_10075 = io_op_bits_active_vfma ? _GEN_8475 : _GEN_7937; // @[sequencer-master.scala 644:39]
  wire  _GEN_10076 = io_op_bits_active_vfma ? _GEN_8476 : _GEN_7938; // @[sequencer-master.scala 644:39]
  wire  _GEN_10077 = io_op_bits_active_vfma ? _GEN_8477 : _GEN_7939; // @[sequencer-master.scala 644:39]
  wire  _GEN_10078 = io_op_bits_active_vfma ? _GEN_8478 : _GEN_7940; // @[sequencer-master.scala 644:39]
  wire  _GEN_10079 = io_op_bits_active_vfma ? _GEN_8479 : _GEN_7941; // @[sequencer-master.scala 644:39]
  wire  _GEN_10080 = io_op_bits_active_vfma ? _GEN_8480 : _GEN_7942; // @[sequencer-master.scala 644:39]
  wire  _GEN_10081 = io_op_bits_active_vfma ? _GEN_8481 : _GEN_7943; // @[sequencer-master.scala 644:39]
  wire  _GEN_10082 = io_op_bits_active_vfma ? _GEN_8482 : _GEN_7944; // @[sequencer-master.scala 644:39]
  wire  _GEN_10083 = io_op_bits_active_vfma ? _GEN_8483 : _GEN_7945; // @[sequencer-master.scala 644:39]
  wire  _GEN_10084 = io_op_bits_active_vfma ? _GEN_8484 : _GEN_7946; // @[sequencer-master.scala 644:39]
  wire  _GEN_10085 = io_op_bits_active_vfma ? _GEN_8485 : _GEN_7947; // @[sequencer-master.scala 644:39]
  wire  _GEN_10086 = io_op_bits_active_vfma ? _GEN_8486 : _GEN_7948; // @[sequencer-master.scala 644:39]
  wire  _GEN_10087 = io_op_bits_active_vfma ? _GEN_8487 : _GEN_7949; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10088 = io_op_bits_active_vfma ? _GEN_8488 : _GEN_7950; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10089 = io_op_bits_active_vfma ? _GEN_8489 : _GEN_7951; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10090 = io_op_bits_active_vfma ? _GEN_8490 : _GEN_7952; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10091 = io_op_bits_active_vfma ? _GEN_8491 : _GEN_7953; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10092 = io_op_bits_active_vfma ? _GEN_8492 : _GEN_7954; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10093 = io_op_bits_active_vfma ? _GEN_8493 : _GEN_7955; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10094 = io_op_bits_active_vfma ? _GEN_8494 : _GEN_7956; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10095 = io_op_bits_active_vfma ? _GEN_8495 : _GEN_7957; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10096 = io_op_bits_active_vfma ? _GEN_8688 : _GEN_7958; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10097 = io_op_bits_active_vfma ? _GEN_8689 : _GEN_7959; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10098 = io_op_bits_active_vfma ? _GEN_8690 : _GEN_7960; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10099 = io_op_bits_active_vfma ? _GEN_8691 : _GEN_7961; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10100 = io_op_bits_active_vfma ? _GEN_8692 : _GEN_7962; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10101 = io_op_bits_active_vfma ? _GEN_8693 : _GEN_7963; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10102 = io_op_bits_active_vfma ? _GEN_8694 : _GEN_7964; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10103 = io_op_bits_active_vfma ? _GEN_8695 : _GEN_7965; // @[sequencer-master.scala 644:39]
  wire  _GEN_10104 = io_op_bits_active_vfma ? _GEN_8704 : _GEN_7966; // @[sequencer-master.scala 644:39]
  wire  _GEN_10105 = io_op_bits_active_vfma ? _GEN_8705 : _GEN_7967; // @[sequencer-master.scala 644:39]
  wire  _GEN_10106 = io_op_bits_active_vfma ? _GEN_8706 : _GEN_7968; // @[sequencer-master.scala 644:39]
  wire  _GEN_10107 = io_op_bits_active_vfma ? _GEN_8707 : _GEN_7969; // @[sequencer-master.scala 644:39]
  wire  _GEN_10108 = io_op_bits_active_vfma ? _GEN_8708 : _GEN_7970; // @[sequencer-master.scala 644:39]
  wire  _GEN_10109 = io_op_bits_active_vfma ? _GEN_8709 : _GEN_7971; // @[sequencer-master.scala 644:39]
  wire  _GEN_10110 = io_op_bits_active_vfma ? _GEN_8710 : _GEN_7972; // @[sequencer-master.scala 644:39]
  wire  _GEN_10111 = io_op_bits_active_vfma ? _GEN_8711 : _GEN_7973; // @[sequencer-master.scala 644:39]
  wire  _GEN_10112 = io_op_bits_active_vfma ? _GEN_8712 : _GEN_7974; // @[sequencer-master.scala 644:39]
  wire  _GEN_10113 = io_op_bits_active_vfma ? _GEN_8713 : _GEN_7975; // @[sequencer-master.scala 644:39]
  wire  _GEN_10114 = io_op_bits_active_vfma ? _GEN_8714 : _GEN_7976; // @[sequencer-master.scala 644:39]
  wire  _GEN_10115 = io_op_bits_active_vfma ? _GEN_8715 : _GEN_7977; // @[sequencer-master.scala 644:39]
  wire  _GEN_10116 = io_op_bits_active_vfma ? _GEN_8716 : _GEN_7978; // @[sequencer-master.scala 644:39]
  wire  _GEN_10117 = io_op_bits_active_vfma ? _GEN_8717 : _GEN_7979; // @[sequencer-master.scala 644:39]
  wire  _GEN_10118 = io_op_bits_active_vfma ? _GEN_8718 : _GEN_7980; // @[sequencer-master.scala 644:39]
  wire  _GEN_10119 = io_op_bits_active_vfma ? _GEN_8719 : _GEN_7981; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10120 = io_op_bits_active_vfma ? _GEN_8720 : _GEN_7982; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10121 = io_op_bits_active_vfma ? _GEN_8721 : _GEN_7983; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10122 = io_op_bits_active_vfma ? _GEN_8722 : _GEN_7984; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10123 = io_op_bits_active_vfma ? _GEN_8723 : _GEN_7985; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10124 = io_op_bits_active_vfma ? _GEN_8724 : _GEN_7986; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10125 = io_op_bits_active_vfma ? _GEN_8725 : _GEN_7987; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10126 = io_op_bits_active_vfma ? _GEN_8726 : _GEN_7988; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10127 = io_op_bits_active_vfma ? _GEN_8727 : _GEN_7989; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10128 = io_op_bits_active_vfma ? _GEN_8728 : _GEN_7990; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10129 = io_op_bits_active_vfma ? _GEN_8729 : _GEN_7991; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10130 = io_op_bits_active_vfma ? _GEN_8730 : _GEN_7992; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10131 = io_op_bits_active_vfma ? _GEN_8731 : _GEN_7993; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10132 = io_op_bits_active_vfma ? _GEN_8732 : _GEN_7994; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10133 = io_op_bits_active_vfma ? _GEN_8733 : _GEN_7995; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10134 = io_op_bits_active_vfma ? _GEN_8734 : _GEN_7996; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10135 = io_op_bits_active_vfma ? _GEN_8735 : _GEN_7997; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10136 = io_op_bits_active_vfma ? _GEN_8736 : _GEN_7998; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10137 = io_op_bits_active_vfma ? _GEN_8737 : _GEN_7999; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10138 = io_op_bits_active_vfma ? _GEN_8738 : _GEN_8000; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10139 = io_op_bits_active_vfma ? _GEN_8739 : _GEN_8001; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10140 = io_op_bits_active_vfma ? _GEN_8740 : _GEN_8002; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10141 = io_op_bits_active_vfma ? _GEN_8741 : _GEN_8003; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10142 = io_op_bits_active_vfma ? _GEN_8742 : _GEN_8004; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10143 = io_op_bits_active_vfma ? _GEN_8743 : _GEN_8005; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10144 = io_op_bits_active_vfma ? _GEN_8936 : _GEN_8006; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10145 = io_op_bits_active_vfma ? _GEN_8937 : _GEN_8007; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10146 = io_op_bits_active_vfma ? _GEN_8938 : _GEN_8008; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10147 = io_op_bits_active_vfma ? _GEN_8939 : _GEN_8009; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10148 = io_op_bits_active_vfma ? _GEN_8940 : _GEN_8010; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10149 = io_op_bits_active_vfma ? _GEN_8941 : _GEN_8011; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10150 = io_op_bits_active_vfma ? _GEN_8942 : _GEN_8012; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10151 = io_op_bits_active_vfma ? _GEN_8943 : _GEN_8013; // @[sequencer-master.scala 644:39]
  wire  _GEN_10152 = io_op_bits_active_vfma ? _GEN_8952 : _GEN_8014; // @[sequencer-master.scala 644:39]
  wire  _GEN_10153 = io_op_bits_active_vfma ? _GEN_8953 : _GEN_8015; // @[sequencer-master.scala 644:39]
  wire  _GEN_10154 = io_op_bits_active_vfma ? _GEN_8954 : _GEN_8016; // @[sequencer-master.scala 644:39]
  wire  _GEN_10155 = io_op_bits_active_vfma ? _GEN_8955 : _GEN_8017; // @[sequencer-master.scala 644:39]
  wire  _GEN_10156 = io_op_bits_active_vfma ? _GEN_8956 : _GEN_8018; // @[sequencer-master.scala 644:39]
  wire  _GEN_10157 = io_op_bits_active_vfma ? _GEN_8957 : _GEN_8019; // @[sequencer-master.scala 644:39]
  wire  _GEN_10158 = io_op_bits_active_vfma ? _GEN_8958 : _GEN_8020; // @[sequencer-master.scala 644:39]
  wire  _GEN_10159 = io_op_bits_active_vfma ? _GEN_8959 : _GEN_8021; // @[sequencer-master.scala 644:39]
  wire  _GEN_10160 = io_op_bits_active_vfma ? _GEN_8960 : _GEN_8022; // @[sequencer-master.scala 644:39]
  wire  _GEN_10161 = io_op_bits_active_vfma ? _GEN_8961 : _GEN_8023; // @[sequencer-master.scala 644:39]
  wire  _GEN_10162 = io_op_bits_active_vfma ? _GEN_8962 : _GEN_8024; // @[sequencer-master.scala 644:39]
  wire  _GEN_10163 = io_op_bits_active_vfma ? _GEN_8963 : _GEN_8025; // @[sequencer-master.scala 644:39]
  wire  _GEN_10164 = io_op_bits_active_vfma ? _GEN_8964 : _GEN_8026; // @[sequencer-master.scala 644:39]
  wire  _GEN_10165 = io_op_bits_active_vfma ? _GEN_8965 : _GEN_8027; // @[sequencer-master.scala 644:39]
  wire  _GEN_10166 = io_op_bits_active_vfma ? _GEN_8966 : _GEN_8028; // @[sequencer-master.scala 644:39]
  wire  _GEN_10167 = io_op_bits_active_vfma ? _GEN_8967 : _GEN_8029; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10168 = io_op_bits_active_vfma ? _GEN_8968 : _GEN_8030; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10169 = io_op_bits_active_vfma ? _GEN_8969 : _GEN_8031; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10170 = io_op_bits_active_vfma ? _GEN_8970 : _GEN_8032; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10171 = io_op_bits_active_vfma ? _GEN_8971 : _GEN_8033; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10172 = io_op_bits_active_vfma ? _GEN_8972 : _GEN_8034; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10173 = io_op_bits_active_vfma ? _GEN_8973 : _GEN_8035; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10174 = io_op_bits_active_vfma ? _GEN_8974 : _GEN_8036; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10175 = io_op_bits_active_vfma ? _GEN_8975 : _GEN_8037; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10176 = io_op_bits_active_vfma ? _GEN_8976 : _GEN_8038; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10177 = io_op_bits_active_vfma ? _GEN_8977 : _GEN_8039; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10178 = io_op_bits_active_vfma ? _GEN_8978 : _GEN_8040; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10179 = io_op_bits_active_vfma ? _GEN_8979 : _GEN_8041; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10180 = io_op_bits_active_vfma ? _GEN_8980 : _GEN_8042; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10181 = io_op_bits_active_vfma ? _GEN_8981 : _GEN_8043; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10182 = io_op_bits_active_vfma ? _GEN_8982 : _GEN_8044; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10183 = io_op_bits_active_vfma ? _GEN_8983 : _GEN_8045; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10184 = io_op_bits_active_vfma ? _GEN_8984 : _GEN_8046; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10185 = io_op_bits_active_vfma ? _GEN_8985 : _GEN_8047; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10186 = io_op_bits_active_vfma ? _GEN_8986 : _GEN_8048; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10187 = io_op_bits_active_vfma ? _GEN_8987 : _GEN_8049; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10188 = io_op_bits_active_vfma ? _GEN_8988 : _GEN_8050; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10189 = io_op_bits_active_vfma ? _GEN_8989 : _GEN_8051; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10190 = io_op_bits_active_vfma ? _GEN_8990 : _GEN_8052; // @[sequencer-master.scala 644:39]
  wire [63:0] _GEN_10191 = io_op_bits_active_vfma ? _GEN_8991 : _GEN_8053; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10224 = io_op_bits_active_vfma ? _GEN_9224 : _GEN_3738; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10225 = io_op_bits_active_vfma ? _GEN_9225 : _GEN_3739; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10226 = io_op_bits_active_vfma ? _GEN_9226 : _GEN_3740; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10227 = io_op_bits_active_vfma ? _GEN_9227 : _GEN_3741; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10228 = io_op_bits_active_vfma ? _GEN_9228 : _GEN_3742; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10229 = io_op_bits_active_vfma ? _GEN_9229 : _GEN_3743; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10230 = io_op_bits_active_vfma ? _GEN_9230 : _GEN_3744; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10231 = io_op_bits_active_vfma ? _GEN_9231 : _GEN_3745; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10240 = io_op_bits_active_vfma ? _GEN_9416 : _GEN_8086; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10241 = io_op_bits_active_vfma ? _GEN_9417 : _GEN_8087; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10242 = io_op_bits_active_vfma ? _GEN_9418 : _GEN_8088; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10243 = io_op_bits_active_vfma ? _GEN_9419 : _GEN_8089; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10244 = io_op_bits_active_vfma ? _GEN_9420 : _GEN_8090; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10245 = io_op_bits_active_vfma ? _GEN_9421 : _GEN_8091; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10246 = io_op_bits_active_vfma ? _GEN_9422 : _GEN_8092; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10247 = io_op_bits_active_vfma ? _GEN_9423 : _GEN_8093; // @[sequencer-master.scala 644:39]
  wire  _GEN_10248 = io_op_bits_active_vfma ? _GEN_9432 : _GEN_8094; // @[sequencer-master.scala 644:39]
  wire  _GEN_10249 = io_op_bits_active_vfma ? _GEN_9433 : _GEN_8095; // @[sequencer-master.scala 644:39]
  wire  _GEN_10250 = io_op_bits_active_vfma ? _GEN_9434 : _GEN_8096; // @[sequencer-master.scala 644:39]
  wire  _GEN_10251 = io_op_bits_active_vfma ? _GEN_9435 : _GEN_8097; // @[sequencer-master.scala 644:39]
  wire  _GEN_10252 = io_op_bits_active_vfma ? _GEN_9436 : _GEN_8098; // @[sequencer-master.scala 644:39]
  wire  _GEN_10253 = io_op_bits_active_vfma ? _GEN_9437 : _GEN_8099; // @[sequencer-master.scala 644:39]
  wire  _GEN_10254 = io_op_bits_active_vfma ? _GEN_9438 : _GEN_8100; // @[sequencer-master.scala 644:39]
  wire  _GEN_10255 = io_op_bits_active_vfma ? _GEN_9439 : _GEN_8101; // @[sequencer-master.scala 644:39]
  wire  _GEN_10256 = io_op_bits_active_vfma ? _GEN_9440 : _GEN_8102; // @[sequencer-master.scala 644:39]
  wire  _GEN_10257 = io_op_bits_active_vfma ? _GEN_9441 : _GEN_8103; // @[sequencer-master.scala 644:39]
  wire  _GEN_10258 = io_op_bits_active_vfma ? _GEN_9442 : _GEN_8104; // @[sequencer-master.scala 644:39]
  wire  _GEN_10259 = io_op_bits_active_vfma ? _GEN_9443 : _GEN_8105; // @[sequencer-master.scala 644:39]
  wire  _GEN_10260 = io_op_bits_active_vfma ? _GEN_9444 : _GEN_8106; // @[sequencer-master.scala 644:39]
  wire  _GEN_10261 = io_op_bits_active_vfma ? _GEN_9445 : _GEN_8107; // @[sequencer-master.scala 644:39]
  wire  _GEN_10262 = io_op_bits_active_vfma ? _GEN_9446 : _GEN_8108; // @[sequencer-master.scala 644:39]
  wire  _GEN_10263 = io_op_bits_active_vfma ? _GEN_9447 : _GEN_8109; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10264 = io_op_bits_active_vfma ? _GEN_9448 : _GEN_8110; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10265 = io_op_bits_active_vfma ? _GEN_9449 : _GEN_8111; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10266 = io_op_bits_active_vfma ? _GEN_9450 : _GEN_8112; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10267 = io_op_bits_active_vfma ? _GEN_9451 : _GEN_8113; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10268 = io_op_bits_active_vfma ? _GEN_9452 : _GEN_8114; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10269 = io_op_bits_active_vfma ? _GEN_9453 : _GEN_8115; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10270 = io_op_bits_active_vfma ? _GEN_9454 : _GEN_8116; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10271 = io_op_bits_active_vfma ? _GEN_9455 : _GEN_8117; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10272 = io_op_bits_active_vfma ? _GEN_9456 : _GEN_8118; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10273 = io_op_bits_active_vfma ? _GEN_9457 : _GEN_8119; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10274 = io_op_bits_active_vfma ? _GEN_9458 : _GEN_8120; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10275 = io_op_bits_active_vfma ? _GEN_9459 : _GEN_8121; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10276 = io_op_bits_active_vfma ? _GEN_9460 : _GEN_8122; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10277 = io_op_bits_active_vfma ? _GEN_9461 : _GEN_8123; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10278 = io_op_bits_active_vfma ? _GEN_9462 : _GEN_8124; // @[sequencer-master.scala 644:39]
  wire [7:0] _GEN_10279 = io_op_bits_active_vfma ? _GEN_9463 : _GEN_8125; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10280 = io_op_bits_active_vfma ? _GEN_9720 : _GEN_8054; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10281 = io_op_bits_active_vfma ? _GEN_9721 : _GEN_8055; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10282 = io_op_bits_active_vfma ? _GEN_9722 : _GEN_8056; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10283 = io_op_bits_active_vfma ? _GEN_9723 : _GEN_8057; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10284 = io_op_bits_active_vfma ? _GEN_9724 : _GEN_8058; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10285 = io_op_bits_active_vfma ? _GEN_9725 : _GEN_8059; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10286 = io_op_bits_active_vfma ? _GEN_9726 : _GEN_8060; // @[sequencer-master.scala 644:39]
  wire [1:0] _GEN_10287 = io_op_bits_active_vfma ? _GEN_9727 : _GEN_8061; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10288 = io_op_bits_active_vfma ? _GEN_9752 : _GEN_8062; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10289 = io_op_bits_active_vfma ? _GEN_9753 : _GEN_8063; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10290 = io_op_bits_active_vfma ? _GEN_9754 : _GEN_8064; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10291 = io_op_bits_active_vfma ? _GEN_9755 : _GEN_8065; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10292 = io_op_bits_active_vfma ? _GEN_9756 : _GEN_8066; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10293 = io_op_bits_active_vfma ? _GEN_9757 : _GEN_8067; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10294 = io_op_bits_active_vfma ? _GEN_9758 : _GEN_8068; // @[sequencer-master.scala 644:39]
  wire [3:0] _GEN_10295 = io_op_bits_active_vfma ? _GEN_9759 : _GEN_8069; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10296 = io_op_bits_active_vfma ? _GEN_9768 : _GEN_8070; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10297 = io_op_bits_active_vfma ? _GEN_9769 : _GEN_8071; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10298 = io_op_bits_active_vfma ? _GEN_9770 : _GEN_8072; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10299 = io_op_bits_active_vfma ? _GEN_9771 : _GEN_8073; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10300 = io_op_bits_active_vfma ? _GEN_9772 : _GEN_8074; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10301 = io_op_bits_active_vfma ? _GEN_9773 : _GEN_8075; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10302 = io_op_bits_active_vfma ? _GEN_9774 : _GEN_8076; // @[sequencer-master.scala 644:39]
  wire [2:0] _GEN_10303 = io_op_bits_active_vfma ? _GEN_9775 : _GEN_8077; // @[sequencer-master.scala 644:39]
  wire  _GEN_10304 = io_op_bits_active_vfma | _GEN_8126; // @[sequencer-master.scala 644:39 sequencer-master.scala 265:41]
  wire [2:0] _GEN_10305 = io_op_bits_active_vfma ? _T_1645 : _GEN_8127; // @[sequencer-master.scala 644:39 sequencer-master.scala 265:66]
  wire  _GEN_10322 = 3'h0 == tail ? 1'h0 : _GEN_9792; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10323 = 3'h1 == tail ? 1'h0 : _GEN_9793; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10324 = 3'h2 == tail ? 1'h0 : _GEN_9794; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10325 = 3'h3 == tail ? 1'h0 : _GEN_9795; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10326 = 3'h4 == tail ? 1'h0 : _GEN_9796; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10327 = 3'h5 == tail ? 1'h0 : _GEN_9797; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10328 = 3'h6 == tail ? 1'h0 : _GEN_9798; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10329 = 3'h7 == tail ? 1'h0 : _GEN_9799; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_10330 = 3'h0 == tail ? 1'h0 : _GEN_9800; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10331 = 3'h1 == tail ? 1'h0 : _GEN_9801; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10332 = 3'h2 == tail ? 1'h0 : _GEN_9802; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10333 = 3'h3 == tail ? 1'h0 : _GEN_9803; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10334 = 3'h4 == tail ? 1'h0 : _GEN_9804; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10335 = 3'h5 == tail ? 1'h0 : _GEN_9805; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10336 = 3'h6 == tail ? 1'h0 : _GEN_9806; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10337 = 3'h7 == tail ? 1'h0 : _GEN_9807; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_10338 = 3'h0 == tail ? 1'h0 : _GEN_9808; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10339 = 3'h1 == tail ? 1'h0 : _GEN_9809; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10340 = 3'h2 == tail ? 1'h0 : _GEN_9810; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10341 = 3'h3 == tail ? 1'h0 : _GEN_9811; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10342 = 3'h4 == tail ? 1'h0 : _GEN_9812; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10343 = 3'h5 == tail ? 1'h0 : _GEN_9813; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10344 = 3'h6 == tail ? 1'h0 : _GEN_9814; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10345 = 3'h7 == tail ? 1'h0 : _GEN_9815; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_10346 = 3'h0 == tail ? 1'h0 : _GEN_9816; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10347 = 3'h1 == tail ? 1'h0 : _GEN_9817; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10348 = 3'h2 == tail ? 1'h0 : _GEN_9818; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10349 = 3'h3 == tail ? 1'h0 : _GEN_9819; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10350 = 3'h4 == tail ? 1'h0 : _GEN_9820; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10351 = 3'h5 == tail ? 1'h0 : _GEN_9821; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10352 = 3'h6 == tail ? 1'h0 : _GEN_9822; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10353 = 3'h7 == tail ? 1'h0 : _GEN_9823; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_10354 = 3'h0 == tail ? 1'h0 : _GEN_9824; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10355 = 3'h1 == tail ? 1'h0 : _GEN_9825; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10356 = 3'h2 == tail ? 1'h0 : _GEN_9826; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10357 = 3'h3 == tail ? 1'h0 : _GEN_9827; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10358 = 3'h4 == tail ? 1'h0 : _GEN_9828; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10359 = 3'h5 == tail ? 1'h0 : _GEN_9829; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10360 = 3'h6 == tail ? 1'h0 : _GEN_9830; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10361 = 3'h7 == tail ? 1'h0 : _GEN_9831; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_10370 = 3'h0 == tail ? 1'h0 : _GEN_9840; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10371 = 3'h1 == tail ? 1'h0 : _GEN_9841; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10372 = 3'h2 == tail ? 1'h0 : _GEN_9842; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10373 = 3'h3 == tail ? 1'h0 : _GEN_9843; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10374 = 3'h4 == tail ? 1'h0 : _GEN_9844; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10375 = 3'h5 == tail ? 1'h0 : _GEN_9845; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10376 = 3'h6 == tail ? 1'h0 : _GEN_9846; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10377 = 3'h7 == tail ? 1'h0 : _GEN_9847; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10378 = 3'h0 == tail ? 1'h0 : _GEN_9848; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10379 = 3'h1 == tail ? 1'h0 : _GEN_9849; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10380 = 3'h2 == tail ? 1'h0 : _GEN_9850; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10381 = 3'h3 == tail ? 1'h0 : _GEN_9851; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10382 = 3'h4 == tail ? 1'h0 : _GEN_9852; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10383 = 3'h5 == tail ? 1'h0 : _GEN_9853; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10384 = 3'h6 == tail ? 1'h0 : _GEN_9854; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10385 = 3'h7 == tail ? 1'h0 : _GEN_9855; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10386 = 3'h0 == tail ? 1'h0 : _GEN_9856; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10387 = 3'h1 == tail ? 1'h0 : _GEN_9857; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10388 = 3'h2 == tail ? 1'h0 : _GEN_9858; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10389 = 3'h3 == tail ? 1'h0 : _GEN_9859; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10390 = 3'h4 == tail ? 1'h0 : _GEN_9860; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10391 = 3'h5 == tail ? 1'h0 : _GEN_9861; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10392 = 3'h6 == tail ? 1'h0 : _GEN_9862; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10393 = 3'h7 == tail ? 1'h0 : _GEN_9863; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10394 = 3'h0 == tail ? 1'h0 : _GEN_9864; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10395 = 3'h1 == tail ? 1'h0 : _GEN_9865; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10396 = 3'h2 == tail ? 1'h0 : _GEN_9866; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10397 = 3'h3 == tail ? 1'h0 : _GEN_9867; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10398 = 3'h4 == tail ? 1'h0 : _GEN_9868; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10399 = 3'h5 == tail ? 1'h0 : _GEN_9869; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10400 = 3'h6 == tail ? 1'h0 : _GEN_9870; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10401 = 3'h7 == tail ? 1'h0 : _GEN_9871; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10402 = 3'h0 == tail ? 1'h0 : _GEN_9872; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10403 = 3'h1 == tail ? 1'h0 : _GEN_9873; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10404 = 3'h2 == tail ? 1'h0 : _GEN_9874; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10405 = 3'h3 == tail ? 1'h0 : _GEN_9875; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10406 = 3'h4 == tail ? 1'h0 : _GEN_9876; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10407 = 3'h5 == tail ? 1'h0 : _GEN_9877; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10408 = 3'h6 == tail ? 1'h0 : _GEN_9878; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10409 = 3'h7 == tail ? 1'h0 : _GEN_9879; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10410 = 3'h0 == tail ? 1'h0 : _GEN_9880; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10411 = 3'h1 == tail ? 1'h0 : _GEN_9881; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10412 = 3'h2 == tail ? 1'h0 : _GEN_9882; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10413 = 3'h3 == tail ? 1'h0 : _GEN_9883; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10414 = 3'h4 == tail ? 1'h0 : _GEN_9884; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10415 = 3'h5 == tail ? 1'h0 : _GEN_9885; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10416 = 3'h6 == tail ? 1'h0 : _GEN_9886; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10417 = 3'h7 == tail ? 1'h0 : _GEN_9887; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10418 = 3'h0 == tail ? 1'h0 : _GEN_9888; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10419 = 3'h1 == tail ? 1'h0 : _GEN_9889; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10420 = 3'h2 == tail ? 1'h0 : _GEN_9890; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10421 = 3'h3 == tail ? 1'h0 : _GEN_9891; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10422 = 3'h4 == tail ? 1'h0 : _GEN_9892; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10423 = 3'h5 == tail ? 1'h0 : _GEN_9893; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10424 = 3'h6 == tail ? 1'h0 : _GEN_9894; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10425 = 3'h7 == tail ? 1'h0 : _GEN_9895; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10426 = 3'h0 == tail ? 1'h0 : _GEN_9896; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10427 = 3'h1 == tail ? 1'h0 : _GEN_9897; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10428 = 3'h2 == tail ? 1'h0 : _GEN_9898; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10429 = 3'h3 == tail ? 1'h0 : _GEN_9899; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10430 = 3'h4 == tail ? 1'h0 : _GEN_9900; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10431 = 3'h5 == tail ? 1'h0 : _GEN_9901; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10432 = 3'h6 == tail ? 1'h0 : _GEN_9902; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10433 = 3'h7 == tail ? 1'h0 : _GEN_9903; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10434 = 3'h0 == tail ? 1'h0 : _GEN_9904; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10435 = 3'h1 == tail ? 1'h0 : _GEN_9905; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10436 = 3'h2 == tail ? 1'h0 : _GEN_9906; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10437 = 3'h3 == tail ? 1'h0 : _GEN_9907; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10438 = 3'h4 == tail ? 1'h0 : _GEN_9908; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10439 = 3'h5 == tail ? 1'h0 : _GEN_9909; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10440 = 3'h6 == tail ? 1'h0 : _GEN_9910; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10441 = 3'h7 == tail ? 1'h0 : _GEN_9911; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10442 = 3'h0 == tail ? 1'h0 : _GEN_9912; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10443 = 3'h1 == tail ? 1'h0 : _GEN_9913; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10444 = 3'h2 == tail ? 1'h0 : _GEN_9914; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10445 = 3'h3 == tail ? 1'h0 : _GEN_9915; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10446 = 3'h4 == tail ? 1'h0 : _GEN_9916; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10447 = 3'h5 == tail ? 1'h0 : _GEN_9917; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10448 = 3'h6 == tail ? 1'h0 : _GEN_9918; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10449 = 3'h7 == tail ? 1'h0 : _GEN_9919; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10450 = 3'h0 == tail ? 1'h0 : _GEN_9920; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10451 = 3'h1 == tail ? 1'h0 : _GEN_9921; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10452 = 3'h2 == tail ? 1'h0 : _GEN_9922; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10453 = 3'h3 == tail ? 1'h0 : _GEN_9923; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10454 = 3'h4 == tail ? 1'h0 : _GEN_9924; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10455 = 3'h5 == tail ? 1'h0 : _GEN_9925; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10456 = 3'h6 == tail ? 1'h0 : _GEN_9926; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10457 = 3'h7 == tail ? 1'h0 : _GEN_9927; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10458 = 3'h0 == tail ? 1'h0 : _GEN_9928; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10459 = 3'h1 == tail ? 1'h0 : _GEN_9929; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10460 = 3'h2 == tail ? 1'h0 : _GEN_9930; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10461 = 3'h3 == tail ? 1'h0 : _GEN_9931; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10462 = 3'h4 == tail ? 1'h0 : _GEN_9932; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10463 = 3'h5 == tail ? 1'h0 : _GEN_9933; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10464 = 3'h6 == tail ? 1'h0 : _GEN_9934; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10465 = 3'h7 == tail ? 1'h0 : _GEN_9935; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10466 = 3'h0 == tail ? 1'h0 : _GEN_9936; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10467 = 3'h1 == tail ? 1'h0 : _GEN_9937; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10468 = 3'h2 == tail ? 1'h0 : _GEN_9938; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10469 = 3'h3 == tail ? 1'h0 : _GEN_9939; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10470 = 3'h4 == tail ? 1'h0 : _GEN_9940; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10471 = 3'h5 == tail ? 1'h0 : _GEN_9941; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10472 = 3'h6 == tail ? 1'h0 : _GEN_9942; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10473 = 3'h7 == tail ? 1'h0 : _GEN_9943; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10474 = 3'h0 == tail ? 1'h0 : _GEN_9944; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10475 = 3'h1 == tail ? 1'h0 : _GEN_9945; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10476 = 3'h2 == tail ? 1'h0 : _GEN_9946; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10477 = 3'h3 == tail ? 1'h0 : _GEN_9947; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10478 = 3'h4 == tail ? 1'h0 : _GEN_9948; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10479 = 3'h5 == tail ? 1'h0 : _GEN_9949; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10480 = 3'h6 == tail ? 1'h0 : _GEN_9950; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10481 = 3'h7 == tail ? 1'h0 : _GEN_9951; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10482 = 3'h0 == tail ? 1'h0 : _GEN_9952; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10483 = 3'h1 == tail ? 1'h0 : _GEN_9953; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10484 = 3'h2 == tail ? 1'h0 : _GEN_9954; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10485 = 3'h3 == tail ? 1'h0 : _GEN_9955; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10486 = 3'h4 == tail ? 1'h0 : _GEN_9956; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10487 = 3'h5 == tail ? 1'h0 : _GEN_9957; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10488 = 3'h6 == tail ? 1'h0 : _GEN_9958; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10489 = 3'h7 == tail ? 1'h0 : _GEN_9959; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10490 = 3'h0 == tail ? 1'h0 : _GEN_9960; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10491 = 3'h1 == tail ? 1'h0 : _GEN_9961; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10492 = 3'h2 == tail ? 1'h0 : _GEN_9962; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10493 = 3'h3 == tail ? 1'h0 : _GEN_9963; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10494 = 3'h4 == tail ? 1'h0 : _GEN_9964; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10495 = 3'h5 == tail ? 1'h0 : _GEN_9965; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10496 = 3'h6 == tail ? 1'h0 : _GEN_9966; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10497 = 3'h7 == tail ? 1'h0 : _GEN_9967; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10498 = 3'h0 == tail ? 1'h0 : _GEN_9968; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10499 = 3'h1 == tail ? 1'h0 : _GEN_9969; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10500 = 3'h2 == tail ? 1'h0 : _GEN_9970; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10501 = 3'h3 == tail ? 1'h0 : _GEN_9971; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10502 = 3'h4 == tail ? 1'h0 : _GEN_9972; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10503 = 3'h5 == tail ? 1'h0 : _GEN_9973; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10504 = 3'h6 == tail ? 1'h0 : _GEN_9974; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10505 = 3'h7 == tail ? 1'h0 : _GEN_9975; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10506 = 3'h0 == tail ? 1'h0 : _GEN_9976; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10507 = 3'h1 == tail ? 1'h0 : _GEN_9977; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10508 = 3'h2 == tail ? 1'h0 : _GEN_9978; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10509 = 3'h3 == tail ? 1'h0 : _GEN_9979; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10510 = 3'h4 == tail ? 1'h0 : _GEN_9980; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10511 = 3'h5 == tail ? 1'h0 : _GEN_9981; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10512 = 3'h6 == tail ? 1'h0 : _GEN_9982; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10513 = 3'h7 == tail ? 1'h0 : _GEN_9983; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10514 = 3'h0 == tail ? 1'h0 : _GEN_9984; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10515 = 3'h1 == tail ? 1'h0 : _GEN_9985; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10516 = 3'h2 == tail ? 1'h0 : _GEN_9986; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10517 = 3'h3 == tail ? 1'h0 : _GEN_9987; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10518 = 3'h4 == tail ? 1'h0 : _GEN_9988; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10519 = 3'h5 == tail ? 1'h0 : _GEN_9989; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10520 = 3'h6 == tail ? 1'h0 : _GEN_9990; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10521 = 3'h7 == tail ? 1'h0 : _GEN_9991; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10522 = 3'h0 == tail ? 1'h0 : _GEN_9992; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10523 = 3'h1 == tail ? 1'h0 : _GEN_9993; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10524 = 3'h2 == tail ? 1'h0 : _GEN_9994; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10525 = 3'h3 == tail ? 1'h0 : _GEN_9995; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10526 = 3'h4 == tail ? 1'h0 : _GEN_9996; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10527 = 3'h5 == tail ? 1'h0 : _GEN_9997; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10528 = 3'h6 == tail ? 1'h0 : _GEN_9998; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10529 = 3'h7 == tail ? 1'h0 : _GEN_9999; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10530 = 3'h0 == tail ? 1'h0 : _GEN_10000; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10531 = 3'h1 == tail ? 1'h0 : _GEN_10001; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10532 = 3'h2 == tail ? 1'h0 : _GEN_10002; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10533 = 3'h3 == tail ? 1'h0 : _GEN_10003; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10534 = 3'h4 == tail ? 1'h0 : _GEN_10004; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10535 = 3'h5 == tail ? 1'h0 : _GEN_10005; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10536 = 3'h6 == tail ? 1'h0 : _GEN_10006; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10537 = 3'h7 == tail ? 1'h0 : _GEN_10007; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10538 = 3'h0 == tail ? 1'h0 : _GEN_10008; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10539 = 3'h1 == tail ? 1'h0 : _GEN_10009; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10540 = 3'h2 == tail ? 1'h0 : _GEN_10010; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10541 = 3'h3 == tail ? 1'h0 : _GEN_10011; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10542 = 3'h4 == tail ? 1'h0 : _GEN_10012; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10543 = 3'h5 == tail ? 1'h0 : _GEN_10013; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10544 = 3'h6 == tail ? 1'h0 : _GEN_10014; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10545 = 3'h7 == tail ? 1'h0 : _GEN_10015; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_10546 = 3'h0 == tail ? 1'h0 : _GEN_10016; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10547 = 3'h1 == tail ? 1'h0 : _GEN_10017; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10548 = 3'h2 == tail ? 1'h0 : _GEN_10018; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10549 = 3'h3 == tail ? 1'h0 : _GEN_10019; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10550 = 3'h4 == tail ? 1'h0 : _GEN_10020; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10551 = 3'h5 == tail ? 1'h0 : _GEN_10021; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10552 = 3'h6 == tail ? 1'h0 : _GEN_10022; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10553 = 3'h7 == tail ? 1'h0 : _GEN_10023; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_10554 = 3'h0 == tail ? 1'h0 : _GEN_10024; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10555 = 3'h1 == tail ? 1'h0 : _GEN_10025; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10556 = 3'h2 == tail ? 1'h0 : _GEN_10026; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10557 = 3'h3 == tail ? 1'h0 : _GEN_10027; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10558 = 3'h4 == tail ? 1'h0 : _GEN_10028; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10559 = 3'h5 == tail ? 1'h0 : _GEN_10029; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10560 = 3'h6 == tail ? 1'h0 : _GEN_10030; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10561 = 3'h7 == tail ? 1'h0 : _GEN_10031; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_10562 = 3'h0 == tail ? 1'h0 : _GEN_10032; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10563 = 3'h1 == tail ? 1'h0 : _GEN_10033; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10564 = 3'h2 == tail ? 1'h0 : _GEN_10034; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10565 = 3'h3 == tail ? 1'h0 : _GEN_10035; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10566 = 3'h4 == tail ? 1'h0 : _GEN_10036; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10567 = 3'h5 == tail ? 1'h0 : _GEN_10037; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10568 = 3'h6 == tail ? 1'h0 : _GEN_10038; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10569 = 3'h7 == tail ? 1'h0 : _GEN_10039; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_10578 = _GEN_32729 | _GEN_7910; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10579 = _GEN_32730 | _GEN_7911; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10580 = _GEN_32731 | _GEN_7912; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10581 = _GEN_32732 | _GEN_7913; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10582 = _GEN_32733 | _GEN_7914; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10583 = _GEN_32734 | _GEN_7915; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10584 = _GEN_32735 | _GEN_7916; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_10585 = _GEN_32736 | _GEN_7917; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_10586 = 3'h0 == tail ? _e_tail_fn_union_2 : _GEN_10056; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10587 = 3'h1 == tail ? _e_tail_fn_union_2 : _GEN_10057; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10588 = 3'h2 == tail ? _e_tail_fn_union_2 : _GEN_10058; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10589 = 3'h3 == tail ? _e_tail_fn_union_2 : _GEN_10059; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10590 = 3'h4 == tail ? _e_tail_fn_union_2 : _GEN_10060; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10591 = 3'h5 == tail ? _e_tail_fn_union_2 : _GEN_10061; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10592 = 3'h6 == tail ? _e_tail_fn_union_2 : _GEN_10062; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_10593 = 3'h7 == tail ? _e_tail_fn_union_2 : _GEN_10063; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_10594 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_10064; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10595 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_10065; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10596 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_10066; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10597 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_10067; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10598 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_10068; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10599 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_10069; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10600 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_10070; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_10601 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_10071; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10602 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_10322; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10603 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_10323; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10604 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_10324; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10605 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_10325; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10606 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_10326; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10607 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_10327; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10608 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_10328; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10609 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_10329; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10610 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_10072; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10611 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_10073; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10612 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_10074; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10613 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_10075; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10614 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_10076; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10615 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_10077; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10616 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_10078; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10617 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_10079; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10618 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_10080; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10619 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_10081; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10620 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_10082; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10621 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_10083; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10622 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_10084; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10623 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_10085; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10624 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_10086; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_10625 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_10087; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_10626 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_10088; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10627 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_10089; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10628 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_10090; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10629 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_10091; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10630 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_10092; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10631 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_10093; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10632 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_10094; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_10633 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_10095; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_10634 = io_op_bits_base_vp_valid ? _GEN_10594 : _GEN_10064; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10635 = io_op_bits_base_vp_valid ? _GEN_10595 : _GEN_10065; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10636 = io_op_bits_base_vp_valid ? _GEN_10596 : _GEN_10066; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10637 = io_op_bits_base_vp_valid ? _GEN_10597 : _GEN_10067; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10638 = io_op_bits_base_vp_valid ? _GEN_10598 : _GEN_10068; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10639 = io_op_bits_base_vp_valid ? _GEN_10599 : _GEN_10069; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10640 = io_op_bits_base_vp_valid ? _GEN_10600 : _GEN_10070; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_10641 = io_op_bits_base_vp_valid ? _GEN_10601 : _GEN_10071; // @[sequencer-master.scala 320:41]
  wire  _GEN_10642 = io_op_bits_base_vp_valid ? _GEN_10602 : _GEN_10322; // @[sequencer-master.scala 320:41]
  wire  _GEN_10643 = io_op_bits_base_vp_valid ? _GEN_10603 : _GEN_10323; // @[sequencer-master.scala 320:41]
  wire  _GEN_10644 = io_op_bits_base_vp_valid ? _GEN_10604 : _GEN_10324; // @[sequencer-master.scala 320:41]
  wire  _GEN_10645 = io_op_bits_base_vp_valid ? _GEN_10605 : _GEN_10325; // @[sequencer-master.scala 320:41]
  wire  _GEN_10646 = io_op_bits_base_vp_valid ? _GEN_10606 : _GEN_10326; // @[sequencer-master.scala 320:41]
  wire  _GEN_10647 = io_op_bits_base_vp_valid ? _GEN_10607 : _GEN_10327; // @[sequencer-master.scala 320:41]
  wire  _GEN_10648 = io_op_bits_base_vp_valid ? _GEN_10608 : _GEN_10328; // @[sequencer-master.scala 320:41]
  wire  _GEN_10649 = io_op_bits_base_vp_valid ? _GEN_10609 : _GEN_10329; // @[sequencer-master.scala 320:41]
  wire  _GEN_10650 = io_op_bits_base_vp_valid ? _GEN_10610 : _GEN_10072; // @[sequencer-master.scala 320:41]
  wire  _GEN_10651 = io_op_bits_base_vp_valid ? _GEN_10611 : _GEN_10073; // @[sequencer-master.scala 320:41]
  wire  _GEN_10652 = io_op_bits_base_vp_valid ? _GEN_10612 : _GEN_10074; // @[sequencer-master.scala 320:41]
  wire  _GEN_10653 = io_op_bits_base_vp_valid ? _GEN_10613 : _GEN_10075; // @[sequencer-master.scala 320:41]
  wire  _GEN_10654 = io_op_bits_base_vp_valid ? _GEN_10614 : _GEN_10076; // @[sequencer-master.scala 320:41]
  wire  _GEN_10655 = io_op_bits_base_vp_valid ? _GEN_10615 : _GEN_10077; // @[sequencer-master.scala 320:41]
  wire  _GEN_10656 = io_op_bits_base_vp_valid ? _GEN_10616 : _GEN_10078; // @[sequencer-master.scala 320:41]
  wire  _GEN_10657 = io_op_bits_base_vp_valid ? _GEN_10617 : _GEN_10079; // @[sequencer-master.scala 320:41]
  wire  _GEN_10658 = io_op_bits_base_vp_valid ? _GEN_10618 : _GEN_10080; // @[sequencer-master.scala 320:41]
  wire  _GEN_10659 = io_op_bits_base_vp_valid ? _GEN_10619 : _GEN_10081; // @[sequencer-master.scala 320:41]
  wire  _GEN_10660 = io_op_bits_base_vp_valid ? _GEN_10620 : _GEN_10082; // @[sequencer-master.scala 320:41]
  wire  _GEN_10661 = io_op_bits_base_vp_valid ? _GEN_10621 : _GEN_10083; // @[sequencer-master.scala 320:41]
  wire  _GEN_10662 = io_op_bits_base_vp_valid ? _GEN_10622 : _GEN_10084; // @[sequencer-master.scala 320:41]
  wire  _GEN_10663 = io_op_bits_base_vp_valid ? _GEN_10623 : _GEN_10085; // @[sequencer-master.scala 320:41]
  wire  _GEN_10664 = io_op_bits_base_vp_valid ? _GEN_10624 : _GEN_10086; // @[sequencer-master.scala 320:41]
  wire  _GEN_10665 = io_op_bits_base_vp_valid ? _GEN_10625 : _GEN_10087; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10666 = io_op_bits_base_vp_valid ? _GEN_10626 : _GEN_10088; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10667 = io_op_bits_base_vp_valid ? _GEN_10627 : _GEN_10089; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10668 = io_op_bits_base_vp_valid ? _GEN_10628 : _GEN_10090; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10669 = io_op_bits_base_vp_valid ? _GEN_10629 : _GEN_10091; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10670 = io_op_bits_base_vp_valid ? _GEN_10630 : _GEN_10092; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10671 = io_op_bits_base_vp_valid ? _GEN_10631 : _GEN_10093; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10672 = io_op_bits_base_vp_valid ? _GEN_10632 : _GEN_10094; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_10673 = io_op_bits_base_vp_valid ? _GEN_10633 : _GEN_10095; // @[sequencer-master.scala 320:41]
  wire  _GEN_10674 = _GEN_32729 | _GEN_10370; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10675 = _GEN_32730 | _GEN_10371; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10676 = _GEN_32731 | _GEN_10372; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10677 = _GEN_32732 | _GEN_10373; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10678 = _GEN_32733 | _GEN_10374; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10679 = _GEN_32734 | _GEN_10375; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10680 = _GEN_32735 | _GEN_10376; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10681 = _GEN_32736 | _GEN_10377; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10682 = _T_26 ? _GEN_10674 : _GEN_10370; // @[sequencer-master.scala 154:24]
  wire  _GEN_10683 = _T_26 ? _GEN_10675 : _GEN_10371; // @[sequencer-master.scala 154:24]
  wire  _GEN_10684 = _T_26 ? _GEN_10676 : _GEN_10372; // @[sequencer-master.scala 154:24]
  wire  _GEN_10685 = _T_26 ? _GEN_10677 : _GEN_10373; // @[sequencer-master.scala 154:24]
  wire  _GEN_10686 = _T_26 ? _GEN_10678 : _GEN_10374; // @[sequencer-master.scala 154:24]
  wire  _GEN_10687 = _T_26 ? _GEN_10679 : _GEN_10375; // @[sequencer-master.scala 154:24]
  wire  _GEN_10688 = _T_26 ? _GEN_10680 : _GEN_10376; // @[sequencer-master.scala 154:24]
  wire  _GEN_10689 = _T_26 ? _GEN_10681 : _GEN_10377; // @[sequencer-master.scala 154:24]
  wire  _GEN_10690 = _GEN_32729 | _GEN_10394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10691 = _GEN_32730 | _GEN_10395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10692 = _GEN_32731 | _GEN_10396; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10693 = _GEN_32732 | _GEN_10397; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10694 = _GEN_32733 | _GEN_10398; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10695 = _GEN_32734 | _GEN_10399; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10696 = _GEN_32735 | _GEN_10400; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10697 = _GEN_32736 | _GEN_10401; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10698 = _T_48 ? _GEN_10690 : _GEN_10394; // @[sequencer-master.scala 154:24]
  wire  _GEN_10699 = _T_48 ? _GEN_10691 : _GEN_10395; // @[sequencer-master.scala 154:24]
  wire  _GEN_10700 = _T_48 ? _GEN_10692 : _GEN_10396; // @[sequencer-master.scala 154:24]
  wire  _GEN_10701 = _T_48 ? _GEN_10693 : _GEN_10397; // @[sequencer-master.scala 154:24]
  wire  _GEN_10702 = _T_48 ? _GEN_10694 : _GEN_10398; // @[sequencer-master.scala 154:24]
  wire  _GEN_10703 = _T_48 ? _GEN_10695 : _GEN_10399; // @[sequencer-master.scala 154:24]
  wire  _GEN_10704 = _T_48 ? _GEN_10696 : _GEN_10400; // @[sequencer-master.scala 154:24]
  wire  _GEN_10705 = _T_48 ? _GEN_10697 : _GEN_10401; // @[sequencer-master.scala 154:24]
  wire  _GEN_10706 = _GEN_32729 | _GEN_10418; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10707 = _GEN_32730 | _GEN_10419; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10708 = _GEN_32731 | _GEN_10420; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10709 = _GEN_32732 | _GEN_10421; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10710 = _GEN_32733 | _GEN_10422; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10711 = _GEN_32734 | _GEN_10423; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10712 = _GEN_32735 | _GEN_10424; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10713 = _GEN_32736 | _GEN_10425; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10714 = _T_70 ? _GEN_10706 : _GEN_10418; // @[sequencer-master.scala 154:24]
  wire  _GEN_10715 = _T_70 ? _GEN_10707 : _GEN_10419; // @[sequencer-master.scala 154:24]
  wire  _GEN_10716 = _T_70 ? _GEN_10708 : _GEN_10420; // @[sequencer-master.scala 154:24]
  wire  _GEN_10717 = _T_70 ? _GEN_10709 : _GEN_10421; // @[sequencer-master.scala 154:24]
  wire  _GEN_10718 = _T_70 ? _GEN_10710 : _GEN_10422; // @[sequencer-master.scala 154:24]
  wire  _GEN_10719 = _T_70 ? _GEN_10711 : _GEN_10423; // @[sequencer-master.scala 154:24]
  wire  _GEN_10720 = _T_70 ? _GEN_10712 : _GEN_10424; // @[sequencer-master.scala 154:24]
  wire  _GEN_10721 = _T_70 ? _GEN_10713 : _GEN_10425; // @[sequencer-master.scala 154:24]
  wire  _GEN_10722 = _GEN_32729 | _GEN_10442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10723 = _GEN_32730 | _GEN_10443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10724 = _GEN_32731 | _GEN_10444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10725 = _GEN_32732 | _GEN_10445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10726 = _GEN_32733 | _GEN_10446; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10727 = _GEN_32734 | _GEN_10447; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10728 = _GEN_32735 | _GEN_10448; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10729 = _GEN_32736 | _GEN_10449; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10730 = _T_92 ? _GEN_10722 : _GEN_10442; // @[sequencer-master.scala 154:24]
  wire  _GEN_10731 = _T_92 ? _GEN_10723 : _GEN_10443; // @[sequencer-master.scala 154:24]
  wire  _GEN_10732 = _T_92 ? _GEN_10724 : _GEN_10444; // @[sequencer-master.scala 154:24]
  wire  _GEN_10733 = _T_92 ? _GEN_10725 : _GEN_10445; // @[sequencer-master.scala 154:24]
  wire  _GEN_10734 = _T_92 ? _GEN_10726 : _GEN_10446; // @[sequencer-master.scala 154:24]
  wire  _GEN_10735 = _T_92 ? _GEN_10727 : _GEN_10447; // @[sequencer-master.scala 154:24]
  wire  _GEN_10736 = _T_92 ? _GEN_10728 : _GEN_10448; // @[sequencer-master.scala 154:24]
  wire  _GEN_10737 = _T_92 ? _GEN_10729 : _GEN_10449; // @[sequencer-master.scala 154:24]
  wire  _GEN_10738 = _GEN_32729 | _GEN_10466; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10739 = _GEN_32730 | _GEN_10467; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10740 = _GEN_32731 | _GEN_10468; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10741 = _GEN_32732 | _GEN_10469; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10742 = _GEN_32733 | _GEN_10470; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10743 = _GEN_32734 | _GEN_10471; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10744 = _GEN_32735 | _GEN_10472; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10745 = _GEN_32736 | _GEN_10473; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10746 = _T_114 ? _GEN_10738 : _GEN_10466; // @[sequencer-master.scala 154:24]
  wire  _GEN_10747 = _T_114 ? _GEN_10739 : _GEN_10467; // @[sequencer-master.scala 154:24]
  wire  _GEN_10748 = _T_114 ? _GEN_10740 : _GEN_10468; // @[sequencer-master.scala 154:24]
  wire  _GEN_10749 = _T_114 ? _GEN_10741 : _GEN_10469; // @[sequencer-master.scala 154:24]
  wire  _GEN_10750 = _T_114 ? _GEN_10742 : _GEN_10470; // @[sequencer-master.scala 154:24]
  wire  _GEN_10751 = _T_114 ? _GEN_10743 : _GEN_10471; // @[sequencer-master.scala 154:24]
  wire  _GEN_10752 = _T_114 ? _GEN_10744 : _GEN_10472; // @[sequencer-master.scala 154:24]
  wire  _GEN_10753 = _T_114 ? _GEN_10745 : _GEN_10473; // @[sequencer-master.scala 154:24]
  wire  _GEN_10754 = _GEN_32729 | _GEN_10490; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10755 = _GEN_32730 | _GEN_10491; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10756 = _GEN_32731 | _GEN_10492; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10757 = _GEN_32732 | _GEN_10493; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10758 = _GEN_32733 | _GEN_10494; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10759 = _GEN_32734 | _GEN_10495; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10760 = _GEN_32735 | _GEN_10496; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10761 = _GEN_32736 | _GEN_10497; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10762 = _T_136 ? _GEN_10754 : _GEN_10490; // @[sequencer-master.scala 154:24]
  wire  _GEN_10763 = _T_136 ? _GEN_10755 : _GEN_10491; // @[sequencer-master.scala 154:24]
  wire  _GEN_10764 = _T_136 ? _GEN_10756 : _GEN_10492; // @[sequencer-master.scala 154:24]
  wire  _GEN_10765 = _T_136 ? _GEN_10757 : _GEN_10493; // @[sequencer-master.scala 154:24]
  wire  _GEN_10766 = _T_136 ? _GEN_10758 : _GEN_10494; // @[sequencer-master.scala 154:24]
  wire  _GEN_10767 = _T_136 ? _GEN_10759 : _GEN_10495; // @[sequencer-master.scala 154:24]
  wire  _GEN_10768 = _T_136 ? _GEN_10760 : _GEN_10496; // @[sequencer-master.scala 154:24]
  wire  _GEN_10769 = _T_136 ? _GEN_10761 : _GEN_10497; // @[sequencer-master.scala 154:24]
  wire  _GEN_10770 = _GEN_32729 | _GEN_10514; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10771 = _GEN_32730 | _GEN_10515; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10772 = _GEN_32731 | _GEN_10516; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10773 = _GEN_32732 | _GEN_10517; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10774 = _GEN_32733 | _GEN_10518; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10775 = _GEN_32734 | _GEN_10519; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10776 = _GEN_32735 | _GEN_10520; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10777 = _GEN_32736 | _GEN_10521; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10778 = _T_158 ? _GEN_10770 : _GEN_10514; // @[sequencer-master.scala 154:24]
  wire  _GEN_10779 = _T_158 ? _GEN_10771 : _GEN_10515; // @[sequencer-master.scala 154:24]
  wire  _GEN_10780 = _T_158 ? _GEN_10772 : _GEN_10516; // @[sequencer-master.scala 154:24]
  wire  _GEN_10781 = _T_158 ? _GEN_10773 : _GEN_10517; // @[sequencer-master.scala 154:24]
  wire  _GEN_10782 = _T_158 ? _GEN_10774 : _GEN_10518; // @[sequencer-master.scala 154:24]
  wire  _GEN_10783 = _T_158 ? _GEN_10775 : _GEN_10519; // @[sequencer-master.scala 154:24]
  wire  _GEN_10784 = _T_158 ? _GEN_10776 : _GEN_10520; // @[sequencer-master.scala 154:24]
  wire  _GEN_10785 = _T_158 ? _GEN_10777 : _GEN_10521; // @[sequencer-master.scala 154:24]
  wire  _GEN_10786 = _GEN_32729 | _GEN_10538; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10787 = _GEN_32730 | _GEN_10539; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10788 = _GEN_32731 | _GEN_10540; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10789 = _GEN_32732 | _GEN_10541; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10790 = _GEN_32733 | _GEN_10542; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10791 = _GEN_32734 | _GEN_10543; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10792 = _GEN_32735 | _GEN_10544; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10793 = _GEN_32736 | _GEN_10545; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10794 = _T_180 ? _GEN_10786 : _GEN_10538; // @[sequencer-master.scala 154:24]
  wire  _GEN_10795 = _T_180 ? _GEN_10787 : _GEN_10539; // @[sequencer-master.scala 154:24]
  wire  _GEN_10796 = _T_180 ? _GEN_10788 : _GEN_10540; // @[sequencer-master.scala 154:24]
  wire  _GEN_10797 = _T_180 ? _GEN_10789 : _GEN_10541; // @[sequencer-master.scala 154:24]
  wire  _GEN_10798 = _T_180 ? _GEN_10790 : _GEN_10542; // @[sequencer-master.scala 154:24]
  wire  _GEN_10799 = _T_180 ? _GEN_10791 : _GEN_10543; // @[sequencer-master.scala 154:24]
  wire  _GEN_10800 = _T_180 ? _GEN_10792 : _GEN_10544; // @[sequencer-master.scala 154:24]
  wire  _GEN_10801 = _T_180 ? _GEN_10793 : _GEN_10545; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_10802 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_10096; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10803 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_10097; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10804 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_10098; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10805 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_10099; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10806 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_10100; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10807 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_10101; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10808 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_10102; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10809 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_10103; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10810 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_10330; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10811 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_10331; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10812 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_10332; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10813 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_10333; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10814 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_10334; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10815 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_10335; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10816 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_10336; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10817 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_10337; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10818 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_10104; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10819 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_10105; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10820 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_10106; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10821 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_10107; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10822 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_10108; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10823 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_10109; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10824 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_10110; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10825 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_10111; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10826 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_10112; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10827 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_10113; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10828 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_10114; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10829 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_10115; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10830 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_10116; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10831 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_10117; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10832 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_10118; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_10833 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_10119; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10834 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_10120; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10835 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_10121; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10836 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_10122; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10837 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_10123; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10838 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_10124; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10839 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_10125; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10840 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_10126; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_10841 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_10127; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_10842 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_10128; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10843 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_10129; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10844 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_10130; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10845 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_10131; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10846 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_10132; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10847 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_10133; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10848 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_10134; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_10849 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_10135; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_10850 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_10136; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10851 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_10137; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10852 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_10138; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10853 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_10139; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10854 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_10140; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10855 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_10141; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10856 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_10142; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10857 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_10143; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_10858 = _T_189 ? _GEN_10850 : _GEN_10136; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10859 = _T_189 ? _GEN_10851 : _GEN_10137; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10860 = _T_189 ? _GEN_10852 : _GEN_10138; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10861 = _T_189 ? _GEN_10853 : _GEN_10139; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10862 = _T_189 ? _GEN_10854 : _GEN_10140; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10863 = _T_189 ? _GEN_10855 : _GEN_10141; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10864 = _T_189 ? _GEN_10856 : _GEN_10142; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_10865 = _T_189 ? _GEN_10857 : _GEN_10143; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_10866 = io_op_bits_base_vs1_valid ? _GEN_10802 : _GEN_10096; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10867 = io_op_bits_base_vs1_valid ? _GEN_10803 : _GEN_10097; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10868 = io_op_bits_base_vs1_valid ? _GEN_10804 : _GEN_10098; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10869 = io_op_bits_base_vs1_valid ? _GEN_10805 : _GEN_10099; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10870 = io_op_bits_base_vs1_valid ? _GEN_10806 : _GEN_10100; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10871 = io_op_bits_base_vs1_valid ? _GEN_10807 : _GEN_10101; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10872 = io_op_bits_base_vs1_valid ? _GEN_10808 : _GEN_10102; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10873 = io_op_bits_base_vs1_valid ? _GEN_10809 : _GEN_10103; // @[sequencer-master.scala 328:47]
  wire  _GEN_10874 = io_op_bits_base_vs1_valid ? _GEN_10810 : _GEN_10330; // @[sequencer-master.scala 328:47]
  wire  _GEN_10875 = io_op_bits_base_vs1_valid ? _GEN_10811 : _GEN_10331; // @[sequencer-master.scala 328:47]
  wire  _GEN_10876 = io_op_bits_base_vs1_valid ? _GEN_10812 : _GEN_10332; // @[sequencer-master.scala 328:47]
  wire  _GEN_10877 = io_op_bits_base_vs1_valid ? _GEN_10813 : _GEN_10333; // @[sequencer-master.scala 328:47]
  wire  _GEN_10878 = io_op_bits_base_vs1_valid ? _GEN_10814 : _GEN_10334; // @[sequencer-master.scala 328:47]
  wire  _GEN_10879 = io_op_bits_base_vs1_valid ? _GEN_10815 : _GEN_10335; // @[sequencer-master.scala 328:47]
  wire  _GEN_10880 = io_op_bits_base_vs1_valid ? _GEN_10816 : _GEN_10336; // @[sequencer-master.scala 328:47]
  wire  _GEN_10881 = io_op_bits_base_vs1_valid ? _GEN_10817 : _GEN_10337; // @[sequencer-master.scala 328:47]
  wire  _GEN_10882 = io_op_bits_base_vs1_valid ? _GEN_10818 : _GEN_10104; // @[sequencer-master.scala 328:47]
  wire  _GEN_10883 = io_op_bits_base_vs1_valid ? _GEN_10819 : _GEN_10105; // @[sequencer-master.scala 328:47]
  wire  _GEN_10884 = io_op_bits_base_vs1_valid ? _GEN_10820 : _GEN_10106; // @[sequencer-master.scala 328:47]
  wire  _GEN_10885 = io_op_bits_base_vs1_valid ? _GEN_10821 : _GEN_10107; // @[sequencer-master.scala 328:47]
  wire  _GEN_10886 = io_op_bits_base_vs1_valid ? _GEN_10822 : _GEN_10108; // @[sequencer-master.scala 328:47]
  wire  _GEN_10887 = io_op_bits_base_vs1_valid ? _GEN_10823 : _GEN_10109; // @[sequencer-master.scala 328:47]
  wire  _GEN_10888 = io_op_bits_base_vs1_valid ? _GEN_10824 : _GEN_10110; // @[sequencer-master.scala 328:47]
  wire  _GEN_10889 = io_op_bits_base_vs1_valid ? _GEN_10825 : _GEN_10111; // @[sequencer-master.scala 328:47]
  wire  _GEN_10890 = io_op_bits_base_vs1_valid ? _GEN_10826 : _GEN_10112; // @[sequencer-master.scala 328:47]
  wire  _GEN_10891 = io_op_bits_base_vs1_valid ? _GEN_10827 : _GEN_10113; // @[sequencer-master.scala 328:47]
  wire  _GEN_10892 = io_op_bits_base_vs1_valid ? _GEN_10828 : _GEN_10114; // @[sequencer-master.scala 328:47]
  wire  _GEN_10893 = io_op_bits_base_vs1_valid ? _GEN_10829 : _GEN_10115; // @[sequencer-master.scala 328:47]
  wire  _GEN_10894 = io_op_bits_base_vs1_valid ? _GEN_10830 : _GEN_10116; // @[sequencer-master.scala 328:47]
  wire  _GEN_10895 = io_op_bits_base_vs1_valid ? _GEN_10831 : _GEN_10117; // @[sequencer-master.scala 328:47]
  wire  _GEN_10896 = io_op_bits_base_vs1_valid ? _GEN_10832 : _GEN_10118; // @[sequencer-master.scala 328:47]
  wire  _GEN_10897 = io_op_bits_base_vs1_valid ? _GEN_10833 : _GEN_10119; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10898 = io_op_bits_base_vs1_valid ? _GEN_10834 : _GEN_10120; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10899 = io_op_bits_base_vs1_valid ? _GEN_10835 : _GEN_10121; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10900 = io_op_bits_base_vs1_valid ? _GEN_10836 : _GEN_10122; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10901 = io_op_bits_base_vs1_valid ? _GEN_10837 : _GEN_10123; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10902 = io_op_bits_base_vs1_valid ? _GEN_10838 : _GEN_10124; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10903 = io_op_bits_base_vs1_valid ? _GEN_10839 : _GEN_10125; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10904 = io_op_bits_base_vs1_valid ? _GEN_10840 : _GEN_10126; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_10905 = io_op_bits_base_vs1_valid ? _GEN_10841 : _GEN_10127; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10906 = io_op_bits_base_vs1_valid ? _GEN_10842 : _GEN_10128; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10907 = io_op_bits_base_vs1_valid ? _GEN_10843 : _GEN_10129; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10908 = io_op_bits_base_vs1_valid ? _GEN_10844 : _GEN_10130; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10909 = io_op_bits_base_vs1_valid ? _GEN_10845 : _GEN_10131; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10910 = io_op_bits_base_vs1_valid ? _GEN_10846 : _GEN_10132; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10911 = io_op_bits_base_vs1_valid ? _GEN_10847 : _GEN_10133; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10912 = io_op_bits_base_vs1_valid ? _GEN_10848 : _GEN_10134; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_10913 = io_op_bits_base_vs1_valid ? _GEN_10849 : _GEN_10135; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10914 = io_op_bits_base_vs1_valid ? _GEN_10858 : _GEN_10136; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10915 = io_op_bits_base_vs1_valid ? _GEN_10859 : _GEN_10137; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10916 = io_op_bits_base_vs1_valid ? _GEN_10860 : _GEN_10138; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10917 = io_op_bits_base_vs1_valid ? _GEN_10861 : _GEN_10139; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10918 = io_op_bits_base_vs1_valid ? _GEN_10862 : _GEN_10140; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10919 = io_op_bits_base_vs1_valid ? _GEN_10863 : _GEN_10141; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10920 = io_op_bits_base_vs1_valid ? _GEN_10864 : _GEN_10142; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_10921 = io_op_bits_base_vs1_valid ? _GEN_10865 : _GEN_10143; // @[sequencer-master.scala 328:47]
  wire  _GEN_10922 = _GEN_32729 | _GEN_10682; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10923 = _GEN_32730 | _GEN_10683; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10924 = _GEN_32731 | _GEN_10684; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10925 = _GEN_32732 | _GEN_10685; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10926 = _GEN_32733 | _GEN_10686; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10927 = _GEN_32734 | _GEN_10687; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10928 = _GEN_32735 | _GEN_10688; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10929 = _GEN_32736 | _GEN_10689; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10930 = _T_203 ? _GEN_10922 : _GEN_10682; // @[sequencer-master.scala 154:24]
  wire  _GEN_10931 = _T_203 ? _GEN_10923 : _GEN_10683; // @[sequencer-master.scala 154:24]
  wire  _GEN_10932 = _T_203 ? _GEN_10924 : _GEN_10684; // @[sequencer-master.scala 154:24]
  wire  _GEN_10933 = _T_203 ? _GEN_10925 : _GEN_10685; // @[sequencer-master.scala 154:24]
  wire  _GEN_10934 = _T_203 ? _GEN_10926 : _GEN_10686; // @[sequencer-master.scala 154:24]
  wire  _GEN_10935 = _T_203 ? _GEN_10927 : _GEN_10687; // @[sequencer-master.scala 154:24]
  wire  _GEN_10936 = _T_203 ? _GEN_10928 : _GEN_10688; // @[sequencer-master.scala 154:24]
  wire  _GEN_10937 = _T_203 ? _GEN_10929 : _GEN_10689; // @[sequencer-master.scala 154:24]
  wire  _GEN_10938 = _GEN_32729 | _GEN_10698; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10939 = _GEN_32730 | _GEN_10699; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10940 = _GEN_32731 | _GEN_10700; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10941 = _GEN_32732 | _GEN_10701; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10942 = _GEN_32733 | _GEN_10702; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10943 = _GEN_32734 | _GEN_10703; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10944 = _GEN_32735 | _GEN_10704; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10945 = _GEN_32736 | _GEN_10705; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10946 = _T_225 ? _GEN_10938 : _GEN_10698; // @[sequencer-master.scala 154:24]
  wire  _GEN_10947 = _T_225 ? _GEN_10939 : _GEN_10699; // @[sequencer-master.scala 154:24]
  wire  _GEN_10948 = _T_225 ? _GEN_10940 : _GEN_10700; // @[sequencer-master.scala 154:24]
  wire  _GEN_10949 = _T_225 ? _GEN_10941 : _GEN_10701; // @[sequencer-master.scala 154:24]
  wire  _GEN_10950 = _T_225 ? _GEN_10942 : _GEN_10702; // @[sequencer-master.scala 154:24]
  wire  _GEN_10951 = _T_225 ? _GEN_10943 : _GEN_10703; // @[sequencer-master.scala 154:24]
  wire  _GEN_10952 = _T_225 ? _GEN_10944 : _GEN_10704; // @[sequencer-master.scala 154:24]
  wire  _GEN_10953 = _T_225 ? _GEN_10945 : _GEN_10705; // @[sequencer-master.scala 154:24]
  wire  _GEN_10954 = _GEN_32729 | _GEN_10714; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10955 = _GEN_32730 | _GEN_10715; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10956 = _GEN_32731 | _GEN_10716; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10957 = _GEN_32732 | _GEN_10717; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10958 = _GEN_32733 | _GEN_10718; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10959 = _GEN_32734 | _GEN_10719; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10960 = _GEN_32735 | _GEN_10720; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10961 = _GEN_32736 | _GEN_10721; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10962 = _T_247 ? _GEN_10954 : _GEN_10714; // @[sequencer-master.scala 154:24]
  wire  _GEN_10963 = _T_247 ? _GEN_10955 : _GEN_10715; // @[sequencer-master.scala 154:24]
  wire  _GEN_10964 = _T_247 ? _GEN_10956 : _GEN_10716; // @[sequencer-master.scala 154:24]
  wire  _GEN_10965 = _T_247 ? _GEN_10957 : _GEN_10717; // @[sequencer-master.scala 154:24]
  wire  _GEN_10966 = _T_247 ? _GEN_10958 : _GEN_10718; // @[sequencer-master.scala 154:24]
  wire  _GEN_10967 = _T_247 ? _GEN_10959 : _GEN_10719; // @[sequencer-master.scala 154:24]
  wire  _GEN_10968 = _T_247 ? _GEN_10960 : _GEN_10720; // @[sequencer-master.scala 154:24]
  wire  _GEN_10969 = _T_247 ? _GEN_10961 : _GEN_10721; // @[sequencer-master.scala 154:24]
  wire  _GEN_10970 = _GEN_32729 | _GEN_10730; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10971 = _GEN_32730 | _GEN_10731; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10972 = _GEN_32731 | _GEN_10732; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10973 = _GEN_32732 | _GEN_10733; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10974 = _GEN_32733 | _GEN_10734; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10975 = _GEN_32734 | _GEN_10735; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10976 = _GEN_32735 | _GEN_10736; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10977 = _GEN_32736 | _GEN_10737; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10978 = _T_269 ? _GEN_10970 : _GEN_10730; // @[sequencer-master.scala 154:24]
  wire  _GEN_10979 = _T_269 ? _GEN_10971 : _GEN_10731; // @[sequencer-master.scala 154:24]
  wire  _GEN_10980 = _T_269 ? _GEN_10972 : _GEN_10732; // @[sequencer-master.scala 154:24]
  wire  _GEN_10981 = _T_269 ? _GEN_10973 : _GEN_10733; // @[sequencer-master.scala 154:24]
  wire  _GEN_10982 = _T_269 ? _GEN_10974 : _GEN_10734; // @[sequencer-master.scala 154:24]
  wire  _GEN_10983 = _T_269 ? _GEN_10975 : _GEN_10735; // @[sequencer-master.scala 154:24]
  wire  _GEN_10984 = _T_269 ? _GEN_10976 : _GEN_10736; // @[sequencer-master.scala 154:24]
  wire  _GEN_10985 = _T_269 ? _GEN_10977 : _GEN_10737; // @[sequencer-master.scala 154:24]
  wire  _GEN_10986 = _GEN_32729 | _GEN_10746; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10987 = _GEN_32730 | _GEN_10747; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10988 = _GEN_32731 | _GEN_10748; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10989 = _GEN_32732 | _GEN_10749; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10990 = _GEN_32733 | _GEN_10750; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10991 = _GEN_32734 | _GEN_10751; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10992 = _GEN_32735 | _GEN_10752; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10993 = _GEN_32736 | _GEN_10753; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_10994 = _T_291 ? _GEN_10986 : _GEN_10746; // @[sequencer-master.scala 154:24]
  wire  _GEN_10995 = _T_291 ? _GEN_10987 : _GEN_10747; // @[sequencer-master.scala 154:24]
  wire  _GEN_10996 = _T_291 ? _GEN_10988 : _GEN_10748; // @[sequencer-master.scala 154:24]
  wire  _GEN_10997 = _T_291 ? _GEN_10989 : _GEN_10749; // @[sequencer-master.scala 154:24]
  wire  _GEN_10998 = _T_291 ? _GEN_10990 : _GEN_10750; // @[sequencer-master.scala 154:24]
  wire  _GEN_10999 = _T_291 ? _GEN_10991 : _GEN_10751; // @[sequencer-master.scala 154:24]
  wire  _GEN_11000 = _T_291 ? _GEN_10992 : _GEN_10752; // @[sequencer-master.scala 154:24]
  wire  _GEN_11001 = _T_291 ? _GEN_10993 : _GEN_10753; // @[sequencer-master.scala 154:24]
  wire  _GEN_11002 = _GEN_32729 | _GEN_10762; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11003 = _GEN_32730 | _GEN_10763; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11004 = _GEN_32731 | _GEN_10764; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11005 = _GEN_32732 | _GEN_10765; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11006 = _GEN_32733 | _GEN_10766; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11007 = _GEN_32734 | _GEN_10767; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11008 = _GEN_32735 | _GEN_10768; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11009 = _GEN_32736 | _GEN_10769; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11010 = _T_313 ? _GEN_11002 : _GEN_10762; // @[sequencer-master.scala 154:24]
  wire  _GEN_11011 = _T_313 ? _GEN_11003 : _GEN_10763; // @[sequencer-master.scala 154:24]
  wire  _GEN_11012 = _T_313 ? _GEN_11004 : _GEN_10764; // @[sequencer-master.scala 154:24]
  wire  _GEN_11013 = _T_313 ? _GEN_11005 : _GEN_10765; // @[sequencer-master.scala 154:24]
  wire  _GEN_11014 = _T_313 ? _GEN_11006 : _GEN_10766; // @[sequencer-master.scala 154:24]
  wire  _GEN_11015 = _T_313 ? _GEN_11007 : _GEN_10767; // @[sequencer-master.scala 154:24]
  wire  _GEN_11016 = _T_313 ? _GEN_11008 : _GEN_10768; // @[sequencer-master.scala 154:24]
  wire  _GEN_11017 = _T_313 ? _GEN_11009 : _GEN_10769; // @[sequencer-master.scala 154:24]
  wire  _GEN_11018 = _GEN_32729 | _GEN_10778; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11019 = _GEN_32730 | _GEN_10779; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11020 = _GEN_32731 | _GEN_10780; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11021 = _GEN_32732 | _GEN_10781; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11022 = _GEN_32733 | _GEN_10782; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11023 = _GEN_32734 | _GEN_10783; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11024 = _GEN_32735 | _GEN_10784; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11025 = _GEN_32736 | _GEN_10785; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11026 = _T_335 ? _GEN_11018 : _GEN_10778; // @[sequencer-master.scala 154:24]
  wire  _GEN_11027 = _T_335 ? _GEN_11019 : _GEN_10779; // @[sequencer-master.scala 154:24]
  wire  _GEN_11028 = _T_335 ? _GEN_11020 : _GEN_10780; // @[sequencer-master.scala 154:24]
  wire  _GEN_11029 = _T_335 ? _GEN_11021 : _GEN_10781; // @[sequencer-master.scala 154:24]
  wire  _GEN_11030 = _T_335 ? _GEN_11022 : _GEN_10782; // @[sequencer-master.scala 154:24]
  wire  _GEN_11031 = _T_335 ? _GEN_11023 : _GEN_10783; // @[sequencer-master.scala 154:24]
  wire  _GEN_11032 = _T_335 ? _GEN_11024 : _GEN_10784; // @[sequencer-master.scala 154:24]
  wire  _GEN_11033 = _T_335 ? _GEN_11025 : _GEN_10785; // @[sequencer-master.scala 154:24]
  wire  _GEN_11034 = _GEN_32729 | _GEN_10794; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11035 = _GEN_32730 | _GEN_10795; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11036 = _GEN_32731 | _GEN_10796; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11037 = _GEN_32732 | _GEN_10797; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11038 = _GEN_32733 | _GEN_10798; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11039 = _GEN_32734 | _GEN_10799; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11040 = _GEN_32735 | _GEN_10800; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11041 = _GEN_32736 | _GEN_10801; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11042 = _T_357 ? _GEN_11034 : _GEN_10794; // @[sequencer-master.scala 154:24]
  wire  _GEN_11043 = _T_357 ? _GEN_11035 : _GEN_10795; // @[sequencer-master.scala 154:24]
  wire  _GEN_11044 = _T_357 ? _GEN_11036 : _GEN_10796; // @[sequencer-master.scala 154:24]
  wire  _GEN_11045 = _T_357 ? _GEN_11037 : _GEN_10797; // @[sequencer-master.scala 154:24]
  wire  _GEN_11046 = _T_357 ? _GEN_11038 : _GEN_10798; // @[sequencer-master.scala 154:24]
  wire  _GEN_11047 = _T_357 ? _GEN_11039 : _GEN_10799; // @[sequencer-master.scala 154:24]
  wire  _GEN_11048 = _T_357 ? _GEN_11040 : _GEN_10800; // @[sequencer-master.scala 154:24]
  wire  _GEN_11049 = _T_357 ? _GEN_11041 : _GEN_10801; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_11050 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_10144; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11051 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_10145; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11052 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_10146; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11053 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_10147; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11054 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_10148; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11055 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_10149; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11056 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_10150; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11057 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_10151; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11058 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_10338; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11059 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_10339; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11060 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_10340; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11061 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_10341; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11062 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_10342; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11063 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_10343; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11064 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_10344; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11065 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_10345; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11066 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_10152; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11067 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_10153; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11068 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_10154; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11069 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_10155; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11070 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_10156; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11071 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_10157; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11072 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_10158; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11073 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_10159; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11074 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_10160; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11075 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_10161; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11076 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_10162; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11077 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_10163; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11078 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_10164; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11079 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_10165; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11080 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_10166; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_11081 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_10167; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11082 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_10168; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11083 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_10169; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11084 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_10170; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11085 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_10171; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11086 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_10172; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11087 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_10173; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11088 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_10174; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_11089 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_10175; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_11090 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_10176; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11091 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_10177; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11092 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_10178; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11093 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_10179; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11094 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_10180; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11095 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_10181; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11096 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_10182; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_11097 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_10183; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_11098 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_10184; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11099 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_10185; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11100 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_10186; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11101 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_10187; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11102 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_10188; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11103 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_10189; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11104 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_10190; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11105 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_10191; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_11106 = _T_366 ? _GEN_11098 : _GEN_10184; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11107 = _T_366 ? _GEN_11099 : _GEN_10185; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11108 = _T_366 ? _GEN_11100 : _GEN_10186; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11109 = _T_366 ? _GEN_11101 : _GEN_10187; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11110 = _T_366 ? _GEN_11102 : _GEN_10188; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11111 = _T_366 ? _GEN_11103 : _GEN_10189; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11112 = _T_366 ? _GEN_11104 : _GEN_10190; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_11113 = _T_366 ? _GEN_11105 : _GEN_10191; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_11114 = io_op_bits_base_vs2_valid ? _GEN_11050 : _GEN_10144; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11115 = io_op_bits_base_vs2_valid ? _GEN_11051 : _GEN_10145; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11116 = io_op_bits_base_vs2_valid ? _GEN_11052 : _GEN_10146; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11117 = io_op_bits_base_vs2_valid ? _GEN_11053 : _GEN_10147; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11118 = io_op_bits_base_vs2_valid ? _GEN_11054 : _GEN_10148; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11119 = io_op_bits_base_vs2_valid ? _GEN_11055 : _GEN_10149; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11120 = io_op_bits_base_vs2_valid ? _GEN_11056 : _GEN_10150; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11121 = io_op_bits_base_vs2_valid ? _GEN_11057 : _GEN_10151; // @[sequencer-master.scala 328:47]
  wire  _GEN_11122 = io_op_bits_base_vs2_valid ? _GEN_11058 : _GEN_10338; // @[sequencer-master.scala 328:47]
  wire  _GEN_11123 = io_op_bits_base_vs2_valid ? _GEN_11059 : _GEN_10339; // @[sequencer-master.scala 328:47]
  wire  _GEN_11124 = io_op_bits_base_vs2_valid ? _GEN_11060 : _GEN_10340; // @[sequencer-master.scala 328:47]
  wire  _GEN_11125 = io_op_bits_base_vs2_valid ? _GEN_11061 : _GEN_10341; // @[sequencer-master.scala 328:47]
  wire  _GEN_11126 = io_op_bits_base_vs2_valid ? _GEN_11062 : _GEN_10342; // @[sequencer-master.scala 328:47]
  wire  _GEN_11127 = io_op_bits_base_vs2_valid ? _GEN_11063 : _GEN_10343; // @[sequencer-master.scala 328:47]
  wire  _GEN_11128 = io_op_bits_base_vs2_valid ? _GEN_11064 : _GEN_10344; // @[sequencer-master.scala 328:47]
  wire  _GEN_11129 = io_op_bits_base_vs2_valid ? _GEN_11065 : _GEN_10345; // @[sequencer-master.scala 328:47]
  wire  _GEN_11130 = io_op_bits_base_vs2_valid ? _GEN_11066 : _GEN_10152; // @[sequencer-master.scala 328:47]
  wire  _GEN_11131 = io_op_bits_base_vs2_valid ? _GEN_11067 : _GEN_10153; // @[sequencer-master.scala 328:47]
  wire  _GEN_11132 = io_op_bits_base_vs2_valid ? _GEN_11068 : _GEN_10154; // @[sequencer-master.scala 328:47]
  wire  _GEN_11133 = io_op_bits_base_vs2_valid ? _GEN_11069 : _GEN_10155; // @[sequencer-master.scala 328:47]
  wire  _GEN_11134 = io_op_bits_base_vs2_valid ? _GEN_11070 : _GEN_10156; // @[sequencer-master.scala 328:47]
  wire  _GEN_11135 = io_op_bits_base_vs2_valid ? _GEN_11071 : _GEN_10157; // @[sequencer-master.scala 328:47]
  wire  _GEN_11136 = io_op_bits_base_vs2_valid ? _GEN_11072 : _GEN_10158; // @[sequencer-master.scala 328:47]
  wire  _GEN_11137 = io_op_bits_base_vs2_valid ? _GEN_11073 : _GEN_10159; // @[sequencer-master.scala 328:47]
  wire  _GEN_11138 = io_op_bits_base_vs2_valid ? _GEN_11074 : _GEN_10160; // @[sequencer-master.scala 328:47]
  wire  _GEN_11139 = io_op_bits_base_vs2_valid ? _GEN_11075 : _GEN_10161; // @[sequencer-master.scala 328:47]
  wire  _GEN_11140 = io_op_bits_base_vs2_valid ? _GEN_11076 : _GEN_10162; // @[sequencer-master.scala 328:47]
  wire  _GEN_11141 = io_op_bits_base_vs2_valid ? _GEN_11077 : _GEN_10163; // @[sequencer-master.scala 328:47]
  wire  _GEN_11142 = io_op_bits_base_vs2_valid ? _GEN_11078 : _GEN_10164; // @[sequencer-master.scala 328:47]
  wire  _GEN_11143 = io_op_bits_base_vs2_valid ? _GEN_11079 : _GEN_10165; // @[sequencer-master.scala 328:47]
  wire  _GEN_11144 = io_op_bits_base_vs2_valid ? _GEN_11080 : _GEN_10166; // @[sequencer-master.scala 328:47]
  wire  _GEN_11145 = io_op_bits_base_vs2_valid ? _GEN_11081 : _GEN_10167; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11146 = io_op_bits_base_vs2_valid ? _GEN_11082 : _GEN_10168; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11147 = io_op_bits_base_vs2_valid ? _GEN_11083 : _GEN_10169; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11148 = io_op_bits_base_vs2_valid ? _GEN_11084 : _GEN_10170; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11149 = io_op_bits_base_vs2_valid ? _GEN_11085 : _GEN_10171; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11150 = io_op_bits_base_vs2_valid ? _GEN_11086 : _GEN_10172; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11151 = io_op_bits_base_vs2_valid ? _GEN_11087 : _GEN_10173; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11152 = io_op_bits_base_vs2_valid ? _GEN_11088 : _GEN_10174; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_11153 = io_op_bits_base_vs2_valid ? _GEN_11089 : _GEN_10175; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11154 = io_op_bits_base_vs2_valid ? _GEN_11090 : _GEN_10176; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11155 = io_op_bits_base_vs2_valid ? _GEN_11091 : _GEN_10177; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11156 = io_op_bits_base_vs2_valid ? _GEN_11092 : _GEN_10178; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11157 = io_op_bits_base_vs2_valid ? _GEN_11093 : _GEN_10179; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11158 = io_op_bits_base_vs2_valid ? _GEN_11094 : _GEN_10180; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11159 = io_op_bits_base_vs2_valid ? _GEN_11095 : _GEN_10181; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11160 = io_op_bits_base_vs2_valid ? _GEN_11096 : _GEN_10182; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_11161 = io_op_bits_base_vs2_valid ? _GEN_11097 : _GEN_10183; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11162 = io_op_bits_base_vs2_valid ? _GEN_11106 : _GEN_10184; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11163 = io_op_bits_base_vs2_valid ? _GEN_11107 : _GEN_10185; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11164 = io_op_bits_base_vs2_valid ? _GEN_11108 : _GEN_10186; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11165 = io_op_bits_base_vs2_valid ? _GEN_11109 : _GEN_10187; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11166 = io_op_bits_base_vs2_valid ? _GEN_11110 : _GEN_10188; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11167 = io_op_bits_base_vs2_valid ? _GEN_11111 : _GEN_10189; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11168 = io_op_bits_base_vs2_valid ? _GEN_11112 : _GEN_10190; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_11169 = io_op_bits_base_vs2_valid ? _GEN_11113 : _GEN_10191; // @[sequencer-master.scala 328:47]
  wire  _GEN_11170 = _GEN_32729 | _GEN_10930; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11171 = _GEN_32730 | _GEN_10931; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11172 = _GEN_32731 | _GEN_10932; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11173 = _GEN_32732 | _GEN_10933; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11174 = _GEN_32733 | _GEN_10934; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11175 = _GEN_32734 | _GEN_10935; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11176 = _GEN_32735 | _GEN_10936; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11177 = _GEN_32736 | _GEN_10937; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11178 = _T_380 ? _GEN_11170 : _GEN_10930; // @[sequencer-master.scala 154:24]
  wire  _GEN_11179 = _T_380 ? _GEN_11171 : _GEN_10931; // @[sequencer-master.scala 154:24]
  wire  _GEN_11180 = _T_380 ? _GEN_11172 : _GEN_10932; // @[sequencer-master.scala 154:24]
  wire  _GEN_11181 = _T_380 ? _GEN_11173 : _GEN_10933; // @[sequencer-master.scala 154:24]
  wire  _GEN_11182 = _T_380 ? _GEN_11174 : _GEN_10934; // @[sequencer-master.scala 154:24]
  wire  _GEN_11183 = _T_380 ? _GEN_11175 : _GEN_10935; // @[sequencer-master.scala 154:24]
  wire  _GEN_11184 = _T_380 ? _GEN_11176 : _GEN_10936; // @[sequencer-master.scala 154:24]
  wire  _GEN_11185 = _T_380 ? _GEN_11177 : _GEN_10937; // @[sequencer-master.scala 154:24]
  wire  _GEN_11186 = _GEN_32729 | _GEN_10946; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11187 = _GEN_32730 | _GEN_10947; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11188 = _GEN_32731 | _GEN_10948; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11189 = _GEN_32732 | _GEN_10949; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11190 = _GEN_32733 | _GEN_10950; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11191 = _GEN_32734 | _GEN_10951; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11192 = _GEN_32735 | _GEN_10952; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11193 = _GEN_32736 | _GEN_10953; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11194 = _T_402 ? _GEN_11186 : _GEN_10946; // @[sequencer-master.scala 154:24]
  wire  _GEN_11195 = _T_402 ? _GEN_11187 : _GEN_10947; // @[sequencer-master.scala 154:24]
  wire  _GEN_11196 = _T_402 ? _GEN_11188 : _GEN_10948; // @[sequencer-master.scala 154:24]
  wire  _GEN_11197 = _T_402 ? _GEN_11189 : _GEN_10949; // @[sequencer-master.scala 154:24]
  wire  _GEN_11198 = _T_402 ? _GEN_11190 : _GEN_10950; // @[sequencer-master.scala 154:24]
  wire  _GEN_11199 = _T_402 ? _GEN_11191 : _GEN_10951; // @[sequencer-master.scala 154:24]
  wire  _GEN_11200 = _T_402 ? _GEN_11192 : _GEN_10952; // @[sequencer-master.scala 154:24]
  wire  _GEN_11201 = _T_402 ? _GEN_11193 : _GEN_10953; // @[sequencer-master.scala 154:24]
  wire  _GEN_11202 = _GEN_32729 | _GEN_10962; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11203 = _GEN_32730 | _GEN_10963; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11204 = _GEN_32731 | _GEN_10964; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11205 = _GEN_32732 | _GEN_10965; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11206 = _GEN_32733 | _GEN_10966; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11207 = _GEN_32734 | _GEN_10967; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11208 = _GEN_32735 | _GEN_10968; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11209 = _GEN_32736 | _GEN_10969; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11210 = _T_424 ? _GEN_11202 : _GEN_10962; // @[sequencer-master.scala 154:24]
  wire  _GEN_11211 = _T_424 ? _GEN_11203 : _GEN_10963; // @[sequencer-master.scala 154:24]
  wire  _GEN_11212 = _T_424 ? _GEN_11204 : _GEN_10964; // @[sequencer-master.scala 154:24]
  wire  _GEN_11213 = _T_424 ? _GEN_11205 : _GEN_10965; // @[sequencer-master.scala 154:24]
  wire  _GEN_11214 = _T_424 ? _GEN_11206 : _GEN_10966; // @[sequencer-master.scala 154:24]
  wire  _GEN_11215 = _T_424 ? _GEN_11207 : _GEN_10967; // @[sequencer-master.scala 154:24]
  wire  _GEN_11216 = _T_424 ? _GEN_11208 : _GEN_10968; // @[sequencer-master.scala 154:24]
  wire  _GEN_11217 = _T_424 ? _GEN_11209 : _GEN_10969; // @[sequencer-master.scala 154:24]
  wire  _GEN_11218 = _GEN_32729 | _GEN_10978; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11219 = _GEN_32730 | _GEN_10979; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11220 = _GEN_32731 | _GEN_10980; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11221 = _GEN_32732 | _GEN_10981; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11222 = _GEN_32733 | _GEN_10982; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11223 = _GEN_32734 | _GEN_10983; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11224 = _GEN_32735 | _GEN_10984; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11225 = _GEN_32736 | _GEN_10985; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11226 = _T_446 ? _GEN_11218 : _GEN_10978; // @[sequencer-master.scala 154:24]
  wire  _GEN_11227 = _T_446 ? _GEN_11219 : _GEN_10979; // @[sequencer-master.scala 154:24]
  wire  _GEN_11228 = _T_446 ? _GEN_11220 : _GEN_10980; // @[sequencer-master.scala 154:24]
  wire  _GEN_11229 = _T_446 ? _GEN_11221 : _GEN_10981; // @[sequencer-master.scala 154:24]
  wire  _GEN_11230 = _T_446 ? _GEN_11222 : _GEN_10982; // @[sequencer-master.scala 154:24]
  wire  _GEN_11231 = _T_446 ? _GEN_11223 : _GEN_10983; // @[sequencer-master.scala 154:24]
  wire  _GEN_11232 = _T_446 ? _GEN_11224 : _GEN_10984; // @[sequencer-master.scala 154:24]
  wire  _GEN_11233 = _T_446 ? _GEN_11225 : _GEN_10985; // @[sequencer-master.scala 154:24]
  wire  _GEN_11234 = _GEN_32729 | _GEN_10994; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11235 = _GEN_32730 | _GEN_10995; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11236 = _GEN_32731 | _GEN_10996; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11237 = _GEN_32732 | _GEN_10997; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11238 = _GEN_32733 | _GEN_10998; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11239 = _GEN_32734 | _GEN_10999; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11240 = _GEN_32735 | _GEN_11000; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11241 = _GEN_32736 | _GEN_11001; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11242 = _T_468 ? _GEN_11234 : _GEN_10994; // @[sequencer-master.scala 154:24]
  wire  _GEN_11243 = _T_468 ? _GEN_11235 : _GEN_10995; // @[sequencer-master.scala 154:24]
  wire  _GEN_11244 = _T_468 ? _GEN_11236 : _GEN_10996; // @[sequencer-master.scala 154:24]
  wire  _GEN_11245 = _T_468 ? _GEN_11237 : _GEN_10997; // @[sequencer-master.scala 154:24]
  wire  _GEN_11246 = _T_468 ? _GEN_11238 : _GEN_10998; // @[sequencer-master.scala 154:24]
  wire  _GEN_11247 = _T_468 ? _GEN_11239 : _GEN_10999; // @[sequencer-master.scala 154:24]
  wire  _GEN_11248 = _T_468 ? _GEN_11240 : _GEN_11000; // @[sequencer-master.scala 154:24]
  wire  _GEN_11249 = _T_468 ? _GEN_11241 : _GEN_11001; // @[sequencer-master.scala 154:24]
  wire  _GEN_11250 = _GEN_32729 | _GEN_11010; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11251 = _GEN_32730 | _GEN_11011; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11252 = _GEN_32731 | _GEN_11012; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11253 = _GEN_32732 | _GEN_11013; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11254 = _GEN_32733 | _GEN_11014; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11255 = _GEN_32734 | _GEN_11015; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11256 = _GEN_32735 | _GEN_11016; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11257 = _GEN_32736 | _GEN_11017; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11258 = _T_490 ? _GEN_11250 : _GEN_11010; // @[sequencer-master.scala 154:24]
  wire  _GEN_11259 = _T_490 ? _GEN_11251 : _GEN_11011; // @[sequencer-master.scala 154:24]
  wire  _GEN_11260 = _T_490 ? _GEN_11252 : _GEN_11012; // @[sequencer-master.scala 154:24]
  wire  _GEN_11261 = _T_490 ? _GEN_11253 : _GEN_11013; // @[sequencer-master.scala 154:24]
  wire  _GEN_11262 = _T_490 ? _GEN_11254 : _GEN_11014; // @[sequencer-master.scala 154:24]
  wire  _GEN_11263 = _T_490 ? _GEN_11255 : _GEN_11015; // @[sequencer-master.scala 154:24]
  wire  _GEN_11264 = _T_490 ? _GEN_11256 : _GEN_11016; // @[sequencer-master.scala 154:24]
  wire  _GEN_11265 = _T_490 ? _GEN_11257 : _GEN_11017; // @[sequencer-master.scala 154:24]
  wire  _GEN_11266 = _GEN_32729 | _GEN_11026; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11267 = _GEN_32730 | _GEN_11027; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11268 = _GEN_32731 | _GEN_11028; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11269 = _GEN_32732 | _GEN_11029; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11270 = _GEN_32733 | _GEN_11030; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11271 = _GEN_32734 | _GEN_11031; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11272 = _GEN_32735 | _GEN_11032; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11273 = _GEN_32736 | _GEN_11033; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11274 = _T_512 ? _GEN_11266 : _GEN_11026; // @[sequencer-master.scala 154:24]
  wire  _GEN_11275 = _T_512 ? _GEN_11267 : _GEN_11027; // @[sequencer-master.scala 154:24]
  wire  _GEN_11276 = _T_512 ? _GEN_11268 : _GEN_11028; // @[sequencer-master.scala 154:24]
  wire  _GEN_11277 = _T_512 ? _GEN_11269 : _GEN_11029; // @[sequencer-master.scala 154:24]
  wire  _GEN_11278 = _T_512 ? _GEN_11270 : _GEN_11030; // @[sequencer-master.scala 154:24]
  wire  _GEN_11279 = _T_512 ? _GEN_11271 : _GEN_11031; // @[sequencer-master.scala 154:24]
  wire  _GEN_11280 = _T_512 ? _GEN_11272 : _GEN_11032; // @[sequencer-master.scala 154:24]
  wire  _GEN_11281 = _T_512 ? _GEN_11273 : _GEN_11033; // @[sequencer-master.scala 154:24]
  wire  _GEN_11282 = _GEN_32729 | _GEN_11042; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11283 = _GEN_32730 | _GEN_11043; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11284 = _GEN_32731 | _GEN_11044; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11285 = _GEN_32732 | _GEN_11045; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11286 = _GEN_32733 | _GEN_11046; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11287 = _GEN_32734 | _GEN_11047; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11288 = _GEN_32735 | _GEN_11048; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11289 = _GEN_32736 | _GEN_11049; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_11290 = _T_534 ? _GEN_11282 : _GEN_11042; // @[sequencer-master.scala 154:24]
  wire  _GEN_11291 = _T_534 ? _GEN_11283 : _GEN_11043; // @[sequencer-master.scala 154:24]
  wire  _GEN_11292 = _T_534 ? _GEN_11284 : _GEN_11044; // @[sequencer-master.scala 154:24]
  wire  _GEN_11293 = _T_534 ? _GEN_11285 : _GEN_11045; // @[sequencer-master.scala 154:24]
  wire  _GEN_11294 = _T_534 ? _GEN_11286 : _GEN_11046; // @[sequencer-master.scala 154:24]
  wire  _GEN_11295 = _T_534 ? _GEN_11287 : _GEN_11047; // @[sequencer-master.scala 154:24]
  wire  _GEN_11296 = _T_534 ? _GEN_11288 : _GEN_11048; // @[sequencer-master.scala 154:24]
  wire  _GEN_11297 = _T_534 ? _GEN_11289 : _GEN_11049; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_11298 = 3'h0 == tail ? _T_1615[1:0] : _GEN_10280; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11299 = 3'h1 == tail ? _T_1615[1:0] : _GEN_10281; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11300 = 3'h2 == tail ? _T_1615[1:0] : _GEN_10282; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11301 = 3'h3 == tail ? _T_1615[1:0] : _GEN_10283; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11302 = 3'h4 == tail ? _T_1615[1:0] : _GEN_10284; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11303 = 3'h5 == tail ? _T_1615[1:0] : _GEN_10285; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11304 = 3'h6 == tail ? _T_1615[1:0] : _GEN_10286; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_11305 = 3'h7 == tail ? _T_1615[1:0] : _GEN_10287; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_11306 = 3'h0 == tail ? 4'h0 : _GEN_10288; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11307 = 3'h1 == tail ? 4'h0 : _GEN_10289; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11308 = 3'h2 == tail ? 4'h0 : _GEN_10290; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11309 = 3'h3 == tail ? 4'h0 : _GEN_10291; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11310 = 3'h4 == tail ? 4'h0 : _GEN_10292; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11311 = 3'h5 == tail ? 4'h0 : _GEN_10293; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11312 = 3'h6 == tail ? 4'h0 : _GEN_10294; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_11313 = 3'h7 == tail ? 4'h0 : _GEN_10295; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_11314 = 3'h0 == tail ? 3'h0 : _GEN_10296; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11315 = 3'h1 == tail ? 3'h0 : _GEN_10297; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11316 = 3'h2 == tail ? 3'h0 : _GEN_10298; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11317 = 3'h3 == tail ? 3'h0 : _GEN_10299; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11318 = 3'h4 == tail ? 3'h0 : _GEN_10300; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11319 = 3'h5 == tail ? 3'h0 : _GEN_10301; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11320 = 3'h6 == tail ? 3'h0 : _GEN_10302; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_11321 = 3'h7 == tail ? 3'h0 : _GEN_10303; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_11322 = _GEN_32729 | _GEN_10378; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11323 = _GEN_32730 | _GEN_10379; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11324 = _GEN_32731 | _GEN_10380; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11325 = _GEN_32732 | _GEN_10381; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11326 = _GEN_32733 | _GEN_10382; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11327 = _GEN_32734 | _GEN_10383; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11328 = _GEN_32735 | _GEN_10384; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11329 = _GEN_32736 | _GEN_10385; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11330 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11322 : _GEN_10378; // @[sequencer-master.scala 161:86]
  wire  _GEN_11331 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11323 : _GEN_10379; // @[sequencer-master.scala 161:86]
  wire  _GEN_11332 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11324 : _GEN_10380; // @[sequencer-master.scala 161:86]
  wire  _GEN_11333 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11325 : _GEN_10381; // @[sequencer-master.scala 161:86]
  wire  _GEN_11334 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11326 : _GEN_10382; // @[sequencer-master.scala 161:86]
  wire  _GEN_11335 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11327 : _GEN_10383; // @[sequencer-master.scala 161:86]
  wire  _GEN_11336 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11328 : _GEN_10384; // @[sequencer-master.scala 161:86]
  wire  _GEN_11337 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11329 : _GEN_10385; // @[sequencer-master.scala 161:86]
  wire  _GEN_11338 = _GEN_32729 | _GEN_10402; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11339 = _GEN_32730 | _GEN_10403; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11340 = _GEN_32731 | _GEN_10404; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11341 = _GEN_32732 | _GEN_10405; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11342 = _GEN_32733 | _GEN_10406; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11343 = _GEN_32734 | _GEN_10407; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11344 = _GEN_32735 | _GEN_10408; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11345 = _GEN_32736 | _GEN_10409; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11346 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11338 : _GEN_10402; // @[sequencer-master.scala 161:86]
  wire  _GEN_11347 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11339 : _GEN_10403; // @[sequencer-master.scala 161:86]
  wire  _GEN_11348 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11340 : _GEN_10404; // @[sequencer-master.scala 161:86]
  wire  _GEN_11349 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11341 : _GEN_10405; // @[sequencer-master.scala 161:86]
  wire  _GEN_11350 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11342 : _GEN_10406; // @[sequencer-master.scala 161:86]
  wire  _GEN_11351 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11343 : _GEN_10407; // @[sequencer-master.scala 161:86]
  wire  _GEN_11352 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11344 : _GEN_10408; // @[sequencer-master.scala 161:86]
  wire  _GEN_11353 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11345 : _GEN_10409; // @[sequencer-master.scala 161:86]
  wire  _GEN_11354 = _GEN_32729 | _GEN_10426; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11355 = _GEN_32730 | _GEN_10427; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11356 = _GEN_32731 | _GEN_10428; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11357 = _GEN_32732 | _GEN_10429; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11358 = _GEN_32733 | _GEN_10430; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11359 = _GEN_32734 | _GEN_10431; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11360 = _GEN_32735 | _GEN_10432; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11361 = _GEN_32736 | _GEN_10433; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11362 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11354 : _GEN_10426; // @[sequencer-master.scala 161:86]
  wire  _GEN_11363 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11355 : _GEN_10427; // @[sequencer-master.scala 161:86]
  wire  _GEN_11364 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11356 : _GEN_10428; // @[sequencer-master.scala 161:86]
  wire  _GEN_11365 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11357 : _GEN_10429; // @[sequencer-master.scala 161:86]
  wire  _GEN_11366 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11358 : _GEN_10430; // @[sequencer-master.scala 161:86]
  wire  _GEN_11367 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11359 : _GEN_10431; // @[sequencer-master.scala 161:86]
  wire  _GEN_11368 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11360 : _GEN_10432; // @[sequencer-master.scala 161:86]
  wire  _GEN_11369 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11361 : _GEN_10433; // @[sequencer-master.scala 161:86]
  wire  _GEN_11370 = _GEN_32729 | _GEN_10450; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11371 = _GEN_32730 | _GEN_10451; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11372 = _GEN_32731 | _GEN_10452; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11373 = _GEN_32732 | _GEN_10453; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11374 = _GEN_32733 | _GEN_10454; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11375 = _GEN_32734 | _GEN_10455; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11376 = _GEN_32735 | _GEN_10456; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11377 = _GEN_32736 | _GEN_10457; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11378 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11370 : _GEN_10450; // @[sequencer-master.scala 161:86]
  wire  _GEN_11379 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11371 : _GEN_10451; // @[sequencer-master.scala 161:86]
  wire  _GEN_11380 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11372 : _GEN_10452; // @[sequencer-master.scala 161:86]
  wire  _GEN_11381 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11373 : _GEN_10453; // @[sequencer-master.scala 161:86]
  wire  _GEN_11382 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11374 : _GEN_10454; // @[sequencer-master.scala 161:86]
  wire  _GEN_11383 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11375 : _GEN_10455; // @[sequencer-master.scala 161:86]
  wire  _GEN_11384 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11376 : _GEN_10456; // @[sequencer-master.scala 161:86]
  wire  _GEN_11385 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_11377 : _GEN_10457; // @[sequencer-master.scala 161:86]
  wire  _GEN_11386 = _GEN_32729 | _GEN_10474; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11387 = _GEN_32730 | _GEN_10475; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11388 = _GEN_32731 | _GEN_10476; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11389 = _GEN_32732 | _GEN_10477; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11390 = _GEN_32733 | _GEN_10478; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11391 = _GEN_32734 | _GEN_10479; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11392 = _GEN_32735 | _GEN_10480; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11393 = _GEN_32736 | _GEN_10481; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11394 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11386 : _GEN_10474; // @[sequencer-master.scala 161:86]
  wire  _GEN_11395 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11387 : _GEN_10475; // @[sequencer-master.scala 161:86]
  wire  _GEN_11396 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11388 : _GEN_10476; // @[sequencer-master.scala 161:86]
  wire  _GEN_11397 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11389 : _GEN_10477; // @[sequencer-master.scala 161:86]
  wire  _GEN_11398 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11390 : _GEN_10478; // @[sequencer-master.scala 161:86]
  wire  _GEN_11399 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11391 : _GEN_10479; // @[sequencer-master.scala 161:86]
  wire  _GEN_11400 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11392 : _GEN_10480; // @[sequencer-master.scala 161:86]
  wire  _GEN_11401 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_11393 : _GEN_10481; // @[sequencer-master.scala 161:86]
  wire  _GEN_11402 = _GEN_32729 | _GEN_10498; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11403 = _GEN_32730 | _GEN_10499; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11404 = _GEN_32731 | _GEN_10500; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11405 = _GEN_32732 | _GEN_10501; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11406 = _GEN_32733 | _GEN_10502; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11407 = _GEN_32734 | _GEN_10503; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11408 = _GEN_32735 | _GEN_10504; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11409 = _GEN_32736 | _GEN_10505; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11410 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11402 : _GEN_10498; // @[sequencer-master.scala 161:86]
  wire  _GEN_11411 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11403 : _GEN_10499; // @[sequencer-master.scala 161:86]
  wire  _GEN_11412 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11404 : _GEN_10500; // @[sequencer-master.scala 161:86]
  wire  _GEN_11413 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11405 : _GEN_10501; // @[sequencer-master.scala 161:86]
  wire  _GEN_11414 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11406 : _GEN_10502; // @[sequencer-master.scala 161:86]
  wire  _GEN_11415 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11407 : _GEN_10503; // @[sequencer-master.scala 161:86]
  wire  _GEN_11416 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11408 : _GEN_10504; // @[sequencer-master.scala 161:86]
  wire  _GEN_11417 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_11409 : _GEN_10505; // @[sequencer-master.scala 161:86]
  wire  _GEN_11418 = _GEN_32729 | _GEN_10522; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11419 = _GEN_32730 | _GEN_10523; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11420 = _GEN_32731 | _GEN_10524; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11421 = _GEN_32732 | _GEN_10525; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11422 = _GEN_32733 | _GEN_10526; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11423 = _GEN_32734 | _GEN_10527; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11424 = _GEN_32735 | _GEN_10528; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11425 = _GEN_32736 | _GEN_10529; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11426 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11418 : _GEN_10522; // @[sequencer-master.scala 161:86]
  wire  _GEN_11427 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11419 : _GEN_10523; // @[sequencer-master.scala 161:86]
  wire  _GEN_11428 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11420 : _GEN_10524; // @[sequencer-master.scala 161:86]
  wire  _GEN_11429 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11421 : _GEN_10525; // @[sequencer-master.scala 161:86]
  wire  _GEN_11430 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11422 : _GEN_10526; // @[sequencer-master.scala 161:86]
  wire  _GEN_11431 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11423 : _GEN_10527; // @[sequencer-master.scala 161:86]
  wire  _GEN_11432 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11424 : _GEN_10528; // @[sequencer-master.scala 161:86]
  wire  _GEN_11433 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_11425 : _GEN_10529; // @[sequencer-master.scala 161:86]
  wire  _GEN_11434 = _GEN_32729 | _GEN_10546; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11435 = _GEN_32730 | _GEN_10547; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11436 = _GEN_32731 | _GEN_10548; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11437 = _GEN_32732 | _GEN_10549; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11438 = _GEN_32733 | _GEN_10550; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11439 = _GEN_32734 | _GEN_10551; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11440 = _GEN_32735 | _GEN_10552; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11441 = _GEN_32736 | _GEN_10553; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11442 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11434 : _GEN_10546; // @[sequencer-master.scala 161:86]
  wire  _GEN_11443 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11435 : _GEN_10547; // @[sequencer-master.scala 161:86]
  wire  _GEN_11444 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11436 : _GEN_10548; // @[sequencer-master.scala 161:86]
  wire  _GEN_11445 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11437 : _GEN_10549; // @[sequencer-master.scala 161:86]
  wire  _GEN_11446 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11438 : _GEN_10550; // @[sequencer-master.scala 161:86]
  wire  _GEN_11447 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11439 : _GEN_10551; // @[sequencer-master.scala 161:86]
  wire  _GEN_11448 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11440 : _GEN_10552; // @[sequencer-master.scala 161:86]
  wire  _GEN_11449 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_11441 : _GEN_10553; // @[sequencer-master.scala 161:86]
  wire  _GEN_11450 = _GEN_32729 | _GEN_10386; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11451 = _GEN_32730 | _GEN_10387; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11452 = _GEN_32731 | _GEN_10388; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11453 = _GEN_32732 | _GEN_10389; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11454 = _GEN_32733 | _GEN_10390; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11455 = _GEN_32734 | _GEN_10391; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11456 = _GEN_32735 | _GEN_10392; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11457 = _GEN_32736 | _GEN_10393; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11458 = _T_1442 ? _GEN_11450 : _GEN_10386; // @[sequencer-master.scala 168:32]
  wire  _GEN_11459 = _T_1442 ? _GEN_11451 : _GEN_10387; // @[sequencer-master.scala 168:32]
  wire  _GEN_11460 = _T_1442 ? _GEN_11452 : _GEN_10388; // @[sequencer-master.scala 168:32]
  wire  _GEN_11461 = _T_1442 ? _GEN_11453 : _GEN_10389; // @[sequencer-master.scala 168:32]
  wire  _GEN_11462 = _T_1442 ? _GEN_11454 : _GEN_10390; // @[sequencer-master.scala 168:32]
  wire  _GEN_11463 = _T_1442 ? _GEN_11455 : _GEN_10391; // @[sequencer-master.scala 168:32]
  wire  _GEN_11464 = _T_1442 ? _GEN_11456 : _GEN_10392; // @[sequencer-master.scala 168:32]
  wire  _GEN_11465 = _T_1442 ? _GEN_11457 : _GEN_10393; // @[sequencer-master.scala 168:32]
  wire  _GEN_11466 = _GEN_32729 | _GEN_10410; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11467 = _GEN_32730 | _GEN_10411; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11468 = _GEN_32731 | _GEN_10412; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11469 = _GEN_32732 | _GEN_10413; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11470 = _GEN_32733 | _GEN_10414; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11471 = _GEN_32734 | _GEN_10415; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11472 = _GEN_32735 | _GEN_10416; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11473 = _GEN_32736 | _GEN_10417; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11474 = _T_1464 ? _GEN_11466 : _GEN_10410; // @[sequencer-master.scala 168:32]
  wire  _GEN_11475 = _T_1464 ? _GEN_11467 : _GEN_10411; // @[sequencer-master.scala 168:32]
  wire  _GEN_11476 = _T_1464 ? _GEN_11468 : _GEN_10412; // @[sequencer-master.scala 168:32]
  wire  _GEN_11477 = _T_1464 ? _GEN_11469 : _GEN_10413; // @[sequencer-master.scala 168:32]
  wire  _GEN_11478 = _T_1464 ? _GEN_11470 : _GEN_10414; // @[sequencer-master.scala 168:32]
  wire  _GEN_11479 = _T_1464 ? _GEN_11471 : _GEN_10415; // @[sequencer-master.scala 168:32]
  wire  _GEN_11480 = _T_1464 ? _GEN_11472 : _GEN_10416; // @[sequencer-master.scala 168:32]
  wire  _GEN_11481 = _T_1464 ? _GEN_11473 : _GEN_10417; // @[sequencer-master.scala 168:32]
  wire  _GEN_11482 = _GEN_32729 | _GEN_10434; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11483 = _GEN_32730 | _GEN_10435; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11484 = _GEN_32731 | _GEN_10436; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11485 = _GEN_32732 | _GEN_10437; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11486 = _GEN_32733 | _GEN_10438; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11487 = _GEN_32734 | _GEN_10439; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11488 = _GEN_32735 | _GEN_10440; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11489 = _GEN_32736 | _GEN_10441; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11490 = _T_1486 ? _GEN_11482 : _GEN_10434; // @[sequencer-master.scala 168:32]
  wire  _GEN_11491 = _T_1486 ? _GEN_11483 : _GEN_10435; // @[sequencer-master.scala 168:32]
  wire  _GEN_11492 = _T_1486 ? _GEN_11484 : _GEN_10436; // @[sequencer-master.scala 168:32]
  wire  _GEN_11493 = _T_1486 ? _GEN_11485 : _GEN_10437; // @[sequencer-master.scala 168:32]
  wire  _GEN_11494 = _T_1486 ? _GEN_11486 : _GEN_10438; // @[sequencer-master.scala 168:32]
  wire  _GEN_11495 = _T_1486 ? _GEN_11487 : _GEN_10439; // @[sequencer-master.scala 168:32]
  wire  _GEN_11496 = _T_1486 ? _GEN_11488 : _GEN_10440; // @[sequencer-master.scala 168:32]
  wire  _GEN_11497 = _T_1486 ? _GEN_11489 : _GEN_10441; // @[sequencer-master.scala 168:32]
  wire  _GEN_11498 = _GEN_32729 | _GEN_10458; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11499 = _GEN_32730 | _GEN_10459; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11500 = _GEN_32731 | _GEN_10460; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11501 = _GEN_32732 | _GEN_10461; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11502 = _GEN_32733 | _GEN_10462; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11503 = _GEN_32734 | _GEN_10463; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11504 = _GEN_32735 | _GEN_10464; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11505 = _GEN_32736 | _GEN_10465; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11506 = _T_1508 ? _GEN_11498 : _GEN_10458; // @[sequencer-master.scala 168:32]
  wire  _GEN_11507 = _T_1508 ? _GEN_11499 : _GEN_10459; // @[sequencer-master.scala 168:32]
  wire  _GEN_11508 = _T_1508 ? _GEN_11500 : _GEN_10460; // @[sequencer-master.scala 168:32]
  wire  _GEN_11509 = _T_1508 ? _GEN_11501 : _GEN_10461; // @[sequencer-master.scala 168:32]
  wire  _GEN_11510 = _T_1508 ? _GEN_11502 : _GEN_10462; // @[sequencer-master.scala 168:32]
  wire  _GEN_11511 = _T_1508 ? _GEN_11503 : _GEN_10463; // @[sequencer-master.scala 168:32]
  wire  _GEN_11512 = _T_1508 ? _GEN_11504 : _GEN_10464; // @[sequencer-master.scala 168:32]
  wire  _GEN_11513 = _T_1508 ? _GEN_11505 : _GEN_10465; // @[sequencer-master.scala 168:32]
  wire  _GEN_11514 = _GEN_32729 | _GEN_10482; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11515 = _GEN_32730 | _GEN_10483; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11516 = _GEN_32731 | _GEN_10484; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11517 = _GEN_32732 | _GEN_10485; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11518 = _GEN_32733 | _GEN_10486; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11519 = _GEN_32734 | _GEN_10487; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11520 = _GEN_32735 | _GEN_10488; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11521 = _GEN_32736 | _GEN_10489; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11522 = _T_1530 ? _GEN_11514 : _GEN_10482; // @[sequencer-master.scala 168:32]
  wire  _GEN_11523 = _T_1530 ? _GEN_11515 : _GEN_10483; // @[sequencer-master.scala 168:32]
  wire  _GEN_11524 = _T_1530 ? _GEN_11516 : _GEN_10484; // @[sequencer-master.scala 168:32]
  wire  _GEN_11525 = _T_1530 ? _GEN_11517 : _GEN_10485; // @[sequencer-master.scala 168:32]
  wire  _GEN_11526 = _T_1530 ? _GEN_11518 : _GEN_10486; // @[sequencer-master.scala 168:32]
  wire  _GEN_11527 = _T_1530 ? _GEN_11519 : _GEN_10487; // @[sequencer-master.scala 168:32]
  wire  _GEN_11528 = _T_1530 ? _GEN_11520 : _GEN_10488; // @[sequencer-master.scala 168:32]
  wire  _GEN_11529 = _T_1530 ? _GEN_11521 : _GEN_10489; // @[sequencer-master.scala 168:32]
  wire  _GEN_11530 = _GEN_32729 | _GEN_10506; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11531 = _GEN_32730 | _GEN_10507; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11532 = _GEN_32731 | _GEN_10508; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11533 = _GEN_32732 | _GEN_10509; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11534 = _GEN_32733 | _GEN_10510; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11535 = _GEN_32734 | _GEN_10511; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11536 = _GEN_32735 | _GEN_10512; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11537 = _GEN_32736 | _GEN_10513; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11538 = _T_1552 ? _GEN_11530 : _GEN_10506; // @[sequencer-master.scala 168:32]
  wire  _GEN_11539 = _T_1552 ? _GEN_11531 : _GEN_10507; // @[sequencer-master.scala 168:32]
  wire  _GEN_11540 = _T_1552 ? _GEN_11532 : _GEN_10508; // @[sequencer-master.scala 168:32]
  wire  _GEN_11541 = _T_1552 ? _GEN_11533 : _GEN_10509; // @[sequencer-master.scala 168:32]
  wire  _GEN_11542 = _T_1552 ? _GEN_11534 : _GEN_10510; // @[sequencer-master.scala 168:32]
  wire  _GEN_11543 = _T_1552 ? _GEN_11535 : _GEN_10511; // @[sequencer-master.scala 168:32]
  wire  _GEN_11544 = _T_1552 ? _GEN_11536 : _GEN_10512; // @[sequencer-master.scala 168:32]
  wire  _GEN_11545 = _T_1552 ? _GEN_11537 : _GEN_10513; // @[sequencer-master.scala 168:32]
  wire  _GEN_11546 = _GEN_32729 | _GEN_10530; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11547 = _GEN_32730 | _GEN_10531; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11548 = _GEN_32731 | _GEN_10532; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11549 = _GEN_32732 | _GEN_10533; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11550 = _GEN_32733 | _GEN_10534; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11551 = _GEN_32734 | _GEN_10535; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11552 = _GEN_32735 | _GEN_10536; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11553 = _GEN_32736 | _GEN_10537; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11554 = _T_1574 ? _GEN_11546 : _GEN_10530; // @[sequencer-master.scala 168:32]
  wire  _GEN_11555 = _T_1574 ? _GEN_11547 : _GEN_10531; // @[sequencer-master.scala 168:32]
  wire  _GEN_11556 = _T_1574 ? _GEN_11548 : _GEN_10532; // @[sequencer-master.scala 168:32]
  wire  _GEN_11557 = _T_1574 ? _GEN_11549 : _GEN_10533; // @[sequencer-master.scala 168:32]
  wire  _GEN_11558 = _T_1574 ? _GEN_11550 : _GEN_10534; // @[sequencer-master.scala 168:32]
  wire  _GEN_11559 = _T_1574 ? _GEN_11551 : _GEN_10535; // @[sequencer-master.scala 168:32]
  wire  _GEN_11560 = _T_1574 ? _GEN_11552 : _GEN_10536; // @[sequencer-master.scala 168:32]
  wire  _GEN_11561 = _T_1574 ? _GEN_11553 : _GEN_10537; // @[sequencer-master.scala 168:32]
  wire  _GEN_11562 = _GEN_32729 | _GEN_10554; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11563 = _GEN_32730 | _GEN_10555; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11564 = _GEN_32731 | _GEN_10556; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11565 = _GEN_32732 | _GEN_10557; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11566 = _GEN_32733 | _GEN_10558; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11567 = _GEN_32734 | _GEN_10559; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11568 = _GEN_32735 | _GEN_10560; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11569 = _GEN_32736 | _GEN_10561; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_11570 = _T_1596 ? _GEN_11562 : _GEN_10554; // @[sequencer-master.scala 168:32]
  wire  _GEN_11571 = _T_1596 ? _GEN_11563 : _GEN_10555; // @[sequencer-master.scala 168:32]
  wire  _GEN_11572 = _T_1596 ? _GEN_11564 : _GEN_10556; // @[sequencer-master.scala 168:32]
  wire  _GEN_11573 = _T_1596 ? _GEN_11565 : _GEN_10557; // @[sequencer-master.scala 168:32]
  wire  _GEN_11574 = _T_1596 ? _GEN_11566 : _GEN_10558; // @[sequencer-master.scala 168:32]
  wire  _GEN_11575 = _T_1596 ? _GEN_11567 : _GEN_10559; // @[sequencer-master.scala 168:32]
  wire  _GEN_11576 = _T_1596 ? _GEN_11568 : _GEN_10560; // @[sequencer-master.scala 168:32]
  wire  _GEN_11577 = _T_1596 ? _GEN_11569 : _GEN_10561; // @[sequencer-master.scala 168:32]
  wire  _GEN_11578 = 3'h0 == _T_1645 | (_GEN_32729 | _GEN_9776); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11579 = 3'h1 == _T_1645 | (_GEN_32730 | _GEN_9777); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11580 = 3'h2 == _T_1645 | (_GEN_32731 | _GEN_9778); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11581 = 3'h3 == _T_1645 | (_GEN_32732 | _GEN_9779); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11582 = 3'h4 == _T_1645 | (_GEN_32733 | _GEN_9780); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11583 = 3'h5 == _T_1645 | (_GEN_32734 | _GEN_9781); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11584 = 3'h6 == _T_1645 | (_GEN_32735 | _GEN_9782); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11585 = 3'h7 == _T_1645 | (_GEN_32736 | _GEN_9783); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_11594 = 3'h0 == _T_1645 ? 1'h0 : _GEN_10642; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11595 = 3'h1 == _T_1645 ? 1'h0 : _GEN_10643; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11596 = 3'h2 == _T_1645 ? 1'h0 : _GEN_10644; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11597 = 3'h3 == _T_1645 ? 1'h0 : _GEN_10645; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11598 = 3'h4 == _T_1645 ? 1'h0 : _GEN_10646; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11599 = 3'h5 == _T_1645 ? 1'h0 : _GEN_10647; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11600 = 3'h6 == _T_1645 ? 1'h0 : _GEN_10648; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11601 = 3'h7 == _T_1645 ? 1'h0 : _GEN_10649; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_11602 = 3'h0 == _T_1645 ? 1'h0 : _GEN_10874; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11603 = 3'h1 == _T_1645 ? 1'h0 : _GEN_10875; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11604 = 3'h2 == _T_1645 ? 1'h0 : _GEN_10876; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11605 = 3'h3 == _T_1645 ? 1'h0 : _GEN_10877; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11606 = 3'h4 == _T_1645 ? 1'h0 : _GEN_10878; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11607 = 3'h5 == _T_1645 ? 1'h0 : _GEN_10879; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11608 = 3'h6 == _T_1645 ? 1'h0 : _GEN_10880; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11609 = 3'h7 == _T_1645 ? 1'h0 : _GEN_10881; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_11610 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11122; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11611 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11123; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11612 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11124; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11613 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11125; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11614 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11126; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11615 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11127; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11616 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11128; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11617 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11129; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_11618 = 3'h0 == _T_1645 ? 1'h0 : _GEN_10346; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11619 = 3'h1 == _T_1645 ? 1'h0 : _GEN_10347; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11620 = 3'h2 == _T_1645 ? 1'h0 : _GEN_10348; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11621 = 3'h3 == _T_1645 ? 1'h0 : _GEN_10349; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11622 = 3'h4 == _T_1645 ? 1'h0 : _GEN_10350; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11623 = 3'h5 == _T_1645 ? 1'h0 : _GEN_10351; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11624 = 3'h6 == _T_1645 ? 1'h0 : _GEN_10352; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11625 = 3'h7 == _T_1645 ? 1'h0 : _GEN_10353; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_11626 = 3'h0 == _T_1645 ? 1'h0 : _GEN_10354; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11627 = 3'h1 == _T_1645 ? 1'h0 : _GEN_10355; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11628 = 3'h2 == _T_1645 ? 1'h0 : _GEN_10356; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11629 = 3'h3 == _T_1645 ? 1'h0 : _GEN_10357; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11630 = 3'h4 == _T_1645 ? 1'h0 : _GEN_10358; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11631 = 3'h5 == _T_1645 ? 1'h0 : _GEN_10359; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11632 = 3'h6 == _T_1645 ? 1'h0 : _GEN_10360; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11633 = 3'h7 == _T_1645 ? 1'h0 : _GEN_10361; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_11634 = _GEN_34121 | (_GEN_32729 | _GEN_9832); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11635 = _GEN_34122 | (_GEN_32730 | _GEN_9833); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11636 = _GEN_34123 | (_GEN_32731 | _GEN_9834); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11637 = _GEN_34124 | (_GEN_32732 | _GEN_9835); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11638 = _GEN_34125 | (_GEN_32733 | _GEN_9836); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11639 = _GEN_34126 | (_GEN_32734 | _GEN_9837); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11640 = _GEN_34127 | (_GEN_32735 | _GEN_9838); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11641 = _GEN_34128 | (_GEN_32736 | _GEN_9839); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_11642 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11178; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11643 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11179; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11644 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11180; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11645 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11181; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11646 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11182; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11647 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11183; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11648 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11184; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11649 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11185; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11650 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11330; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11651 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11331; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11652 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11332; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11653 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11333; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11654 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11334; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11655 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11335; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11656 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11336; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11657 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11337; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11658 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11458; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11659 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11459; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11660 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11460; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11661 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11461; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11662 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11462; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11663 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11463; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11664 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11464; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11665 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11465; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11666 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11194; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11667 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11195; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11668 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11196; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11669 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11197; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11670 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11198; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11671 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11199; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11672 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11200; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11673 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11201; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11674 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11346; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11675 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11347; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11676 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11348; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11677 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11349; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11678 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11350; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11679 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11351; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11680 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11352; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11681 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11353; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11682 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11474; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11683 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11475; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11684 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11476; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11685 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11477; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11686 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11478; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11687 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11479; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11688 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11480; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11689 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11481; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11690 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11210; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11691 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11211; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11692 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11212; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11693 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11213; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11694 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11214; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11695 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11215; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11696 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11216; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11697 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11217; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11698 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11362; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11699 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11363; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11700 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11364; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11701 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11365; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11702 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11366; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11703 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11367; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11704 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11368; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11705 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11369; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11706 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11490; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11707 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11491; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11708 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11492; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11709 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11493; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11710 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11494; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11711 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11495; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11712 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11496; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11713 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11497; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11714 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11226; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11715 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11227; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11716 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11228; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11717 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11229; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11718 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11230; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11719 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11231; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11720 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11232; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11721 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11233; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11722 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11378; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11723 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11379; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11724 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11380; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11725 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11381; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11726 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11382; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11727 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11383; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11728 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11384; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11729 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11385; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11730 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11506; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11731 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11507; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11732 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11508; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11733 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11509; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11734 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11510; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11735 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11511; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11736 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11512; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11737 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11513; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11738 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11242; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11739 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11243; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11740 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11244; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11741 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11245; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11742 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11246; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11743 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11247; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11744 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11248; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11745 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11249; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11746 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11394; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11747 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11395; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11748 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11396; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11749 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11397; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11750 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11398; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11751 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11399; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11752 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11400; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11753 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11401; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11754 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11522; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11755 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11523; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11756 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11524; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11757 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11525; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11758 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11526; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11759 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11527; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11760 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11528; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11761 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11529; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11762 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11258; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11763 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11259; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11764 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11260; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11765 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11261; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11766 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11262; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11767 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11263; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11768 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11264; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11769 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11265; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11770 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11410; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11771 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11411; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11772 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11412; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11773 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11413; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11774 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11414; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11775 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11415; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11776 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11416; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11777 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11417; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11778 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11538; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11779 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11539; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11780 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11540; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11781 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11541; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11782 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11542; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11783 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11543; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11784 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11544; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11785 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11545; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11786 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11274; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11787 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11275; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11788 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11276; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11789 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11277; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11790 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11278; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11791 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11279; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11792 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11280; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11793 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11281; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11794 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11426; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11795 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11427; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11796 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11428; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11797 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11429; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11798 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11430; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11799 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11431; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11800 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11432; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11801 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11433; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11802 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11554; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11803 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11555; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11804 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11556; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11805 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11557; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11806 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11558; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11807 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11559; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11808 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11560; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11809 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11561; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11810 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11290; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11811 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11291; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11812 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11292; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11813 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11293; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11814 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11294; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11815 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11295; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11816 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11296; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11817 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11297; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_11818 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11442; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11819 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11443; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11820 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11444; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11821 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11445; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11822 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11446; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11823 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11447; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11824 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11448; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11825 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11449; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_11826 = 3'h0 == _T_1645 ? 1'h0 : _GEN_11570; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11827 = 3'h1 == _T_1645 ? 1'h0 : _GEN_11571; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11828 = 3'h2 == _T_1645 ? 1'h0 : _GEN_11572; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11829 = 3'h3 == _T_1645 ? 1'h0 : _GEN_11573; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11830 = 3'h4 == _T_1645 ? 1'h0 : _GEN_11574; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11831 = 3'h5 == _T_1645 ? 1'h0 : _GEN_11575; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11832 = 3'h6 == _T_1645 ? 1'h0 : _GEN_11576; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11833 = 3'h7 == _T_1645 ? 1'h0 : _GEN_11577; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_11834 = 3'h0 == _T_1645 ? 1'h0 : _GEN_10562; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11835 = 3'h1 == _T_1645 ? 1'h0 : _GEN_10563; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11836 = 3'h2 == _T_1645 ? 1'h0 : _GEN_10564; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11837 = 3'h3 == _T_1645 ? 1'h0 : _GEN_10565; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11838 = 3'h4 == _T_1645 ? 1'h0 : _GEN_10566; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11839 = 3'h5 == _T_1645 ? 1'h0 : _GEN_10567; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11840 = 3'h6 == _T_1645 ? 1'h0 : _GEN_10568; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11841 = 3'h7 == _T_1645 ? 1'h0 : _GEN_10569; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_11850 = _GEN_34121 | e_0_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11851 = _GEN_34122 | e_1_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11852 = _GEN_34123 | e_2_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11853 = _GEN_34124 | e_3_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11854 = _GEN_34125 | e_4_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11855 = _GEN_34126 | e_5_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11856 = _GEN_34127 | e_6_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_11857 = _GEN_34128 | e_7_active_vfdu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_11858 = 3'h0 == _T_1645 ? io_op_bits_fn_union : _GEN_10586; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11859 = 3'h1 == _T_1645 ? io_op_bits_fn_union : _GEN_10587; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11860 = 3'h2 == _T_1645 ? io_op_bits_fn_union : _GEN_10588; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11861 = 3'h3 == _T_1645 ? io_op_bits_fn_union : _GEN_10589; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11862 = 3'h4 == _T_1645 ? io_op_bits_fn_union : _GEN_10590; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11863 = 3'h5 == _T_1645 ? io_op_bits_fn_union : _GEN_10591; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11864 = 3'h6 == _T_1645 ? io_op_bits_fn_union : _GEN_10592; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_11865 = 3'h7 == _T_1645 ? io_op_bits_fn_union : _GEN_10593; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [7:0] _GEN_11866 = 3'h0 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10240; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11867 = 3'h1 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10241; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11868 = 3'h2 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10242; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11869 = 3'h3 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10243; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11870 = 3'h4 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10244; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11871 = 3'h5 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10245; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11872 = 3'h6 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10246; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11873 = 3'h7 == _T_1645 ? io_op_bits_base_vd_id : _GEN_10247; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11874 = 3'h0 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11626; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11875 = 3'h1 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11627; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11876 = 3'h2 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11628; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11877 = 3'h3 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11629; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11878 = 3'h4 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11630; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11879 = 3'h5 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11631; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11880 = 3'h6 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11632; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11881 = 3'h7 == _T_1645 ? io_op_bits_base_vd_valid : _GEN_11633; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11882 = 3'h0 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10248; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11883 = 3'h1 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10249; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11884 = 3'h2 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10250; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11885 = 3'h3 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10251; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11886 = 3'h4 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10252; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11887 = 3'h5 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10253; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11888 = 3'h6 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10254; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11889 = 3'h7 == _T_1645 ? io_op_bits_base_vd_scalar : _GEN_10255; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11890 = 3'h0 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10256; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11891 = 3'h1 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10257; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11892 = 3'h2 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10258; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11893 = 3'h3 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10259; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11894 = 3'h4 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10260; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11895 = 3'h5 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10261; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11896 = 3'h6 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10262; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_11897 = 3'h7 == _T_1645 ? io_op_bits_base_vd_pred : _GEN_10263; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11898 = 3'h0 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10264; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11899 = 3'h1 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10265; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11900 = 3'h2 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10266; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11901 = 3'h3 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10267; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11902 = 3'h4 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10268; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11903 = 3'h5 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10269; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11904 = 3'h6 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10270; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_11905 = 3'h7 == _T_1645 ? io_op_bits_base_vd_prec : _GEN_10271; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_11906 = 3'h0 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10272; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11907 = 3'h1 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10273; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11908 = 3'h2 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10274; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11909 = 3'h3 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10275; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11910 = 3'h4 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10276; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11911 = 3'h5 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10277; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11912 = 3'h6 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10278; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11913 = 3'h7 == _T_1645 ? io_op_bits_reg_vd_id : _GEN_10279; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_11914 = io_op_bits_base_vd_valid ? _GEN_11866 : _GEN_10240; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11915 = io_op_bits_base_vd_valid ? _GEN_11867 : _GEN_10241; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11916 = io_op_bits_base_vd_valid ? _GEN_11868 : _GEN_10242; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11917 = io_op_bits_base_vd_valid ? _GEN_11869 : _GEN_10243; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11918 = io_op_bits_base_vd_valid ? _GEN_11870 : _GEN_10244; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11919 = io_op_bits_base_vd_valid ? _GEN_11871 : _GEN_10245; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11920 = io_op_bits_base_vd_valid ? _GEN_11872 : _GEN_10246; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11921 = io_op_bits_base_vd_valid ? _GEN_11873 : _GEN_10247; // @[sequencer-master.scala 362:41]
  wire  _GEN_11922 = io_op_bits_base_vd_valid ? _GEN_11874 : _GEN_11626; // @[sequencer-master.scala 362:41]
  wire  _GEN_11923 = io_op_bits_base_vd_valid ? _GEN_11875 : _GEN_11627; // @[sequencer-master.scala 362:41]
  wire  _GEN_11924 = io_op_bits_base_vd_valid ? _GEN_11876 : _GEN_11628; // @[sequencer-master.scala 362:41]
  wire  _GEN_11925 = io_op_bits_base_vd_valid ? _GEN_11877 : _GEN_11629; // @[sequencer-master.scala 362:41]
  wire  _GEN_11926 = io_op_bits_base_vd_valid ? _GEN_11878 : _GEN_11630; // @[sequencer-master.scala 362:41]
  wire  _GEN_11927 = io_op_bits_base_vd_valid ? _GEN_11879 : _GEN_11631; // @[sequencer-master.scala 362:41]
  wire  _GEN_11928 = io_op_bits_base_vd_valid ? _GEN_11880 : _GEN_11632; // @[sequencer-master.scala 362:41]
  wire  _GEN_11929 = io_op_bits_base_vd_valid ? _GEN_11881 : _GEN_11633; // @[sequencer-master.scala 362:41]
  wire  _GEN_11930 = io_op_bits_base_vd_valid ? _GEN_11882 : _GEN_10248; // @[sequencer-master.scala 362:41]
  wire  _GEN_11931 = io_op_bits_base_vd_valid ? _GEN_11883 : _GEN_10249; // @[sequencer-master.scala 362:41]
  wire  _GEN_11932 = io_op_bits_base_vd_valid ? _GEN_11884 : _GEN_10250; // @[sequencer-master.scala 362:41]
  wire  _GEN_11933 = io_op_bits_base_vd_valid ? _GEN_11885 : _GEN_10251; // @[sequencer-master.scala 362:41]
  wire  _GEN_11934 = io_op_bits_base_vd_valid ? _GEN_11886 : _GEN_10252; // @[sequencer-master.scala 362:41]
  wire  _GEN_11935 = io_op_bits_base_vd_valid ? _GEN_11887 : _GEN_10253; // @[sequencer-master.scala 362:41]
  wire  _GEN_11936 = io_op_bits_base_vd_valid ? _GEN_11888 : _GEN_10254; // @[sequencer-master.scala 362:41]
  wire  _GEN_11937 = io_op_bits_base_vd_valid ? _GEN_11889 : _GEN_10255; // @[sequencer-master.scala 362:41]
  wire  _GEN_11938 = io_op_bits_base_vd_valid ? _GEN_11890 : _GEN_10256; // @[sequencer-master.scala 362:41]
  wire  _GEN_11939 = io_op_bits_base_vd_valid ? _GEN_11891 : _GEN_10257; // @[sequencer-master.scala 362:41]
  wire  _GEN_11940 = io_op_bits_base_vd_valid ? _GEN_11892 : _GEN_10258; // @[sequencer-master.scala 362:41]
  wire  _GEN_11941 = io_op_bits_base_vd_valid ? _GEN_11893 : _GEN_10259; // @[sequencer-master.scala 362:41]
  wire  _GEN_11942 = io_op_bits_base_vd_valid ? _GEN_11894 : _GEN_10260; // @[sequencer-master.scala 362:41]
  wire  _GEN_11943 = io_op_bits_base_vd_valid ? _GEN_11895 : _GEN_10261; // @[sequencer-master.scala 362:41]
  wire  _GEN_11944 = io_op_bits_base_vd_valid ? _GEN_11896 : _GEN_10262; // @[sequencer-master.scala 362:41]
  wire  _GEN_11945 = io_op_bits_base_vd_valid ? _GEN_11897 : _GEN_10263; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11946 = io_op_bits_base_vd_valid ? _GEN_11898 : _GEN_10264; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11947 = io_op_bits_base_vd_valid ? _GEN_11899 : _GEN_10265; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11948 = io_op_bits_base_vd_valid ? _GEN_11900 : _GEN_10266; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11949 = io_op_bits_base_vd_valid ? _GEN_11901 : _GEN_10267; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11950 = io_op_bits_base_vd_valid ? _GEN_11902 : _GEN_10268; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11951 = io_op_bits_base_vd_valid ? _GEN_11903 : _GEN_10269; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11952 = io_op_bits_base_vd_valid ? _GEN_11904 : _GEN_10270; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_11953 = io_op_bits_base_vd_valid ? _GEN_11905 : _GEN_10271; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11954 = io_op_bits_base_vd_valid ? _GEN_11906 : _GEN_10272; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11955 = io_op_bits_base_vd_valid ? _GEN_11907 : _GEN_10273; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11956 = io_op_bits_base_vd_valid ? _GEN_11908 : _GEN_10274; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11957 = io_op_bits_base_vd_valid ? _GEN_11909 : _GEN_10275; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11958 = io_op_bits_base_vd_valid ? _GEN_11910 : _GEN_10276; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11959 = io_op_bits_base_vd_valid ? _GEN_11911 : _GEN_10277; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11960 = io_op_bits_base_vd_valid ? _GEN_11912 : _GEN_10278; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_11961 = io_op_bits_base_vd_valid ? _GEN_11913 : _GEN_10279; // @[sequencer-master.scala 362:41]
  wire  _GEN_11962 = _GEN_34121 | _GEN_11650; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11963 = _GEN_34122 | _GEN_11651; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11964 = _GEN_34123 | _GEN_11652; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11965 = _GEN_34124 | _GEN_11653; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11966 = _GEN_34125 | _GEN_11654; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11967 = _GEN_34126 | _GEN_11655; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11968 = _GEN_34127 | _GEN_11656; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11969 = _GEN_34128 | _GEN_11657; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11970 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11962 : _GEN_11650; // @[sequencer-master.scala 161:86]
  wire  _GEN_11971 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11963 : _GEN_11651; // @[sequencer-master.scala 161:86]
  wire  _GEN_11972 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11964 : _GEN_11652; // @[sequencer-master.scala 161:86]
  wire  _GEN_11973 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11965 : _GEN_11653; // @[sequencer-master.scala 161:86]
  wire  _GEN_11974 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11966 : _GEN_11654; // @[sequencer-master.scala 161:86]
  wire  _GEN_11975 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11967 : _GEN_11655; // @[sequencer-master.scala 161:86]
  wire  _GEN_11976 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11968 : _GEN_11656; // @[sequencer-master.scala 161:86]
  wire  _GEN_11977 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_11969 : _GEN_11657; // @[sequencer-master.scala 161:86]
  wire  _GEN_11978 = _GEN_34121 | _GEN_11674; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11979 = _GEN_34122 | _GEN_11675; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11980 = _GEN_34123 | _GEN_11676; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11981 = _GEN_34124 | _GEN_11677; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11982 = _GEN_34125 | _GEN_11678; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11983 = _GEN_34126 | _GEN_11679; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11984 = _GEN_34127 | _GEN_11680; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11985 = _GEN_34128 | _GEN_11681; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11986 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11978 : _GEN_11674; // @[sequencer-master.scala 161:86]
  wire  _GEN_11987 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11979 : _GEN_11675; // @[sequencer-master.scala 161:86]
  wire  _GEN_11988 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11980 : _GEN_11676; // @[sequencer-master.scala 161:86]
  wire  _GEN_11989 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11981 : _GEN_11677; // @[sequencer-master.scala 161:86]
  wire  _GEN_11990 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11982 : _GEN_11678; // @[sequencer-master.scala 161:86]
  wire  _GEN_11991 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11983 : _GEN_11679; // @[sequencer-master.scala 161:86]
  wire  _GEN_11992 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11984 : _GEN_11680; // @[sequencer-master.scala 161:86]
  wire  _GEN_11993 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_11985 : _GEN_11681; // @[sequencer-master.scala 161:86]
  wire  _GEN_11994 = _GEN_34121 | _GEN_11698; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11995 = _GEN_34122 | _GEN_11699; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11996 = _GEN_34123 | _GEN_11700; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11997 = _GEN_34124 | _GEN_11701; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11998 = _GEN_34125 | _GEN_11702; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_11999 = _GEN_34126 | _GEN_11703; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12000 = _GEN_34127 | _GEN_11704; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12001 = _GEN_34128 | _GEN_11705; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12002 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11994 : _GEN_11698; // @[sequencer-master.scala 161:86]
  wire  _GEN_12003 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11995 : _GEN_11699; // @[sequencer-master.scala 161:86]
  wire  _GEN_12004 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11996 : _GEN_11700; // @[sequencer-master.scala 161:86]
  wire  _GEN_12005 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11997 : _GEN_11701; // @[sequencer-master.scala 161:86]
  wire  _GEN_12006 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11998 : _GEN_11702; // @[sequencer-master.scala 161:86]
  wire  _GEN_12007 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_11999 : _GEN_11703; // @[sequencer-master.scala 161:86]
  wire  _GEN_12008 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_12000 : _GEN_11704; // @[sequencer-master.scala 161:86]
  wire  _GEN_12009 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_12001 : _GEN_11705; // @[sequencer-master.scala 161:86]
  wire  _GEN_12010 = _GEN_34121 | _GEN_11722; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12011 = _GEN_34122 | _GEN_11723; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12012 = _GEN_34123 | _GEN_11724; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12013 = _GEN_34124 | _GEN_11725; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12014 = _GEN_34125 | _GEN_11726; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12015 = _GEN_34126 | _GEN_11727; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12016 = _GEN_34127 | _GEN_11728; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12017 = _GEN_34128 | _GEN_11729; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12018 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12010 : _GEN_11722; // @[sequencer-master.scala 161:86]
  wire  _GEN_12019 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12011 : _GEN_11723; // @[sequencer-master.scala 161:86]
  wire  _GEN_12020 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12012 : _GEN_11724; // @[sequencer-master.scala 161:86]
  wire  _GEN_12021 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12013 : _GEN_11725; // @[sequencer-master.scala 161:86]
  wire  _GEN_12022 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12014 : _GEN_11726; // @[sequencer-master.scala 161:86]
  wire  _GEN_12023 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12015 : _GEN_11727; // @[sequencer-master.scala 161:86]
  wire  _GEN_12024 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12016 : _GEN_11728; // @[sequencer-master.scala 161:86]
  wire  _GEN_12025 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_12017 : _GEN_11729; // @[sequencer-master.scala 161:86]
  wire  _GEN_12026 = _GEN_34121 | _GEN_11746; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12027 = _GEN_34122 | _GEN_11747; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12028 = _GEN_34123 | _GEN_11748; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12029 = _GEN_34124 | _GEN_11749; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12030 = _GEN_34125 | _GEN_11750; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12031 = _GEN_34126 | _GEN_11751; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12032 = _GEN_34127 | _GEN_11752; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12033 = _GEN_34128 | _GEN_11753; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12034 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12026 : _GEN_11746; // @[sequencer-master.scala 161:86]
  wire  _GEN_12035 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12027 : _GEN_11747; // @[sequencer-master.scala 161:86]
  wire  _GEN_12036 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12028 : _GEN_11748; // @[sequencer-master.scala 161:86]
  wire  _GEN_12037 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12029 : _GEN_11749; // @[sequencer-master.scala 161:86]
  wire  _GEN_12038 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12030 : _GEN_11750; // @[sequencer-master.scala 161:86]
  wire  _GEN_12039 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12031 : _GEN_11751; // @[sequencer-master.scala 161:86]
  wire  _GEN_12040 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12032 : _GEN_11752; // @[sequencer-master.scala 161:86]
  wire  _GEN_12041 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_12033 : _GEN_11753; // @[sequencer-master.scala 161:86]
  wire  _GEN_12042 = _GEN_34121 | _GEN_11770; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12043 = _GEN_34122 | _GEN_11771; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12044 = _GEN_34123 | _GEN_11772; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12045 = _GEN_34124 | _GEN_11773; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12046 = _GEN_34125 | _GEN_11774; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12047 = _GEN_34126 | _GEN_11775; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12048 = _GEN_34127 | _GEN_11776; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12049 = _GEN_34128 | _GEN_11777; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12050 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12042 : _GEN_11770; // @[sequencer-master.scala 161:86]
  wire  _GEN_12051 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12043 : _GEN_11771; // @[sequencer-master.scala 161:86]
  wire  _GEN_12052 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12044 : _GEN_11772; // @[sequencer-master.scala 161:86]
  wire  _GEN_12053 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12045 : _GEN_11773; // @[sequencer-master.scala 161:86]
  wire  _GEN_12054 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12046 : _GEN_11774; // @[sequencer-master.scala 161:86]
  wire  _GEN_12055 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12047 : _GEN_11775; // @[sequencer-master.scala 161:86]
  wire  _GEN_12056 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12048 : _GEN_11776; // @[sequencer-master.scala 161:86]
  wire  _GEN_12057 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_12049 : _GEN_11777; // @[sequencer-master.scala 161:86]
  wire  _GEN_12058 = _GEN_34121 | _GEN_11794; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12059 = _GEN_34122 | _GEN_11795; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12060 = _GEN_34123 | _GEN_11796; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12061 = _GEN_34124 | _GEN_11797; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12062 = _GEN_34125 | _GEN_11798; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12063 = _GEN_34126 | _GEN_11799; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12064 = _GEN_34127 | _GEN_11800; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12065 = _GEN_34128 | _GEN_11801; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12066 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12058 : _GEN_11794; // @[sequencer-master.scala 161:86]
  wire  _GEN_12067 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12059 : _GEN_11795; // @[sequencer-master.scala 161:86]
  wire  _GEN_12068 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12060 : _GEN_11796; // @[sequencer-master.scala 161:86]
  wire  _GEN_12069 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12061 : _GEN_11797; // @[sequencer-master.scala 161:86]
  wire  _GEN_12070 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12062 : _GEN_11798; // @[sequencer-master.scala 161:86]
  wire  _GEN_12071 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12063 : _GEN_11799; // @[sequencer-master.scala 161:86]
  wire  _GEN_12072 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12064 : _GEN_11800; // @[sequencer-master.scala 161:86]
  wire  _GEN_12073 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_12065 : _GEN_11801; // @[sequencer-master.scala 161:86]
  wire  _GEN_12074 = _GEN_34121 | _GEN_11818; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12075 = _GEN_34122 | _GEN_11819; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12076 = _GEN_34123 | _GEN_11820; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12077 = _GEN_34124 | _GEN_11821; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12078 = _GEN_34125 | _GEN_11822; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12079 = _GEN_34126 | _GEN_11823; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12080 = _GEN_34127 | _GEN_11824; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12081 = _GEN_34128 | _GEN_11825; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_12082 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12074 : _GEN_11818; // @[sequencer-master.scala 161:86]
  wire  _GEN_12083 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12075 : _GEN_11819; // @[sequencer-master.scala 161:86]
  wire  _GEN_12084 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12076 : _GEN_11820; // @[sequencer-master.scala 161:86]
  wire  _GEN_12085 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12077 : _GEN_11821; // @[sequencer-master.scala 161:86]
  wire  _GEN_12086 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12078 : _GEN_11822; // @[sequencer-master.scala 161:86]
  wire  _GEN_12087 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12079 : _GEN_11823; // @[sequencer-master.scala 161:86]
  wire  _GEN_12088 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12080 : _GEN_11824; // @[sequencer-master.scala 161:86]
  wire  _GEN_12089 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_12081 : _GEN_11825; // @[sequencer-master.scala 161:86]
  wire  _GEN_12090 = _GEN_34121 | _GEN_11658; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12091 = _GEN_34122 | _GEN_11659; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12092 = _GEN_34123 | _GEN_11660; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12093 = _GEN_34124 | _GEN_11661; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12094 = _GEN_34125 | _GEN_11662; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12095 = _GEN_34126 | _GEN_11663; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12096 = _GEN_34127 | _GEN_11664; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12097 = _GEN_34128 | _GEN_11665; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12098 = _T_1442 ? _GEN_12090 : _GEN_11658; // @[sequencer-master.scala 168:32]
  wire  _GEN_12099 = _T_1442 ? _GEN_12091 : _GEN_11659; // @[sequencer-master.scala 168:32]
  wire  _GEN_12100 = _T_1442 ? _GEN_12092 : _GEN_11660; // @[sequencer-master.scala 168:32]
  wire  _GEN_12101 = _T_1442 ? _GEN_12093 : _GEN_11661; // @[sequencer-master.scala 168:32]
  wire  _GEN_12102 = _T_1442 ? _GEN_12094 : _GEN_11662; // @[sequencer-master.scala 168:32]
  wire  _GEN_12103 = _T_1442 ? _GEN_12095 : _GEN_11663; // @[sequencer-master.scala 168:32]
  wire  _GEN_12104 = _T_1442 ? _GEN_12096 : _GEN_11664; // @[sequencer-master.scala 168:32]
  wire  _GEN_12105 = _T_1442 ? _GEN_12097 : _GEN_11665; // @[sequencer-master.scala 168:32]
  wire  _GEN_12106 = _GEN_34121 | _GEN_11682; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12107 = _GEN_34122 | _GEN_11683; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12108 = _GEN_34123 | _GEN_11684; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12109 = _GEN_34124 | _GEN_11685; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12110 = _GEN_34125 | _GEN_11686; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12111 = _GEN_34126 | _GEN_11687; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12112 = _GEN_34127 | _GEN_11688; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12113 = _GEN_34128 | _GEN_11689; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12114 = _T_1464 ? _GEN_12106 : _GEN_11682; // @[sequencer-master.scala 168:32]
  wire  _GEN_12115 = _T_1464 ? _GEN_12107 : _GEN_11683; // @[sequencer-master.scala 168:32]
  wire  _GEN_12116 = _T_1464 ? _GEN_12108 : _GEN_11684; // @[sequencer-master.scala 168:32]
  wire  _GEN_12117 = _T_1464 ? _GEN_12109 : _GEN_11685; // @[sequencer-master.scala 168:32]
  wire  _GEN_12118 = _T_1464 ? _GEN_12110 : _GEN_11686; // @[sequencer-master.scala 168:32]
  wire  _GEN_12119 = _T_1464 ? _GEN_12111 : _GEN_11687; // @[sequencer-master.scala 168:32]
  wire  _GEN_12120 = _T_1464 ? _GEN_12112 : _GEN_11688; // @[sequencer-master.scala 168:32]
  wire  _GEN_12121 = _T_1464 ? _GEN_12113 : _GEN_11689; // @[sequencer-master.scala 168:32]
  wire  _GEN_12122 = _GEN_34121 | _GEN_11706; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12123 = _GEN_34122 | _GEN_11707; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12124 = _GEN_34123 | _GEN_11708; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12125 = _GEN_34124 | _GEN_11709; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12126 = _GEN_34125 | _GEN_11710; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12127 = _GEN_34126 | _GEN_11711; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12128 = _GEN_34127 | _GEN_11712; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12129 = _GEN_34128 | _GEN_11713; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12130 = _T_1486 ? _GEN_12122 : _GEN_11706; // @[sequencer-master.scala 168:32]
  wire  _GEN_12131 = _T_1486 ? _GEN_12123 : _GEN_11707; // @[sequencer-master.scala 168:32]
  wire  _GEN_12132 = _T_1486 ? _GEN_12124 : _GEN_11708; // @[sequencer-master.scala 168:32]
  wire  _GEN_12133 = _T_1486 ? _GEN_12125 : _GEN_11709; // @[sequencer-master.scala 168:32]
  wire  _GEN_12134 = _T_1486 ? _GEN_12126 : _GEN_11710; // @[sequencer-master.scala 168:32]
  wire  _GEN_12135 = _T_1486 ? _GEN_12127 : _GEN_11711; // @[sequencer-master.scala 168:32]
  wire  _GEN_12136 = _T_1486 ? _GEN_12128 : _GEN_11712; // @[sequencer-master.scala 168:32]
  wire  _GEN_12137 = _T_1486 ? _GEN_12129 : _GEN_11713; // @[sequencer-master.scala 168:32]
  wire  _GEN_12138 = _GEN_34121 | _GEN_11730; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12139 = _GEN_34122 | _GEN_11731; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12140 = _GEN_34123 | _GEN_11732; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12141 = _GEN_34124 | _GEN_11733; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12142 = _GEN_34125 | _GEN_11734; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12143 = _GEN_34126 | _GEN_11735; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12144 = _GEN_34127 | _GEN_11736; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12145 = _GEN_34128 | _GEN_11737; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12146 = _T_1508 ? _GEN_12138 : _GEN_11730; // @[sequencer-master.scala 168:32]
  wire  _GEN_12147 = _T_1508 ? _GEN_12139 : _GEN_11731; // @[sequencer-master.scala 168:32]
  wire  _GEN_12148 = _T_1508 ? _GEN_12140 : _GEN_11732; // @[sequencer-master.scala 168:32]
  wire  _GEN_12149 = _T_1508 ? _GEN_12141 : _GEN_11733; // @[sequencer-master.scala 168:32]
  wire  _GEN_12150 = _T_1508 ? _GEN_12142 : _GEN_11734; // @[sequencer-master.scala 168:32]
  wire  _GEN_12151 = _T_1508 ? _GEN_12143 : _GEN_11735; // @[sequencer-master.scala 168:32]
  wire  _GEN_12152 = _T_1508 ? _GEN_12144 : _GEN_11736; // @[sequencer-master.scala 168:32]
  wire  _GEN_12153 = _T_1508 ? _GEN_12145 : _GEN_11737; // @[sequencer-master.scala 168:32]
  wire  _GEN_12154 = _GEN_34121 | _GEN_11754; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12155 = _GEN_34122 | _GEN_11755; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12156 = _GEN_34123 | _GEN_11756; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12157 = _GEN_34124 | _GEN_11757; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12158 = _GEN_34125 | _GEN_11758; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12159 = _GEN_34126 | _GEN_11759; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12160 = _GEN_34127 | _GEN_11760; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12161 = _GEN_34128 | _GEN_11761; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12162 = _T_1530 ? _GEN_12154 : _GEN_11754; // @[sequencer-master.scala 168:32]
  wire  _GEN_12163 = _T_1530 ? _GEN_12155 : _GEN_11755; // @[sequencer-master.scala 168:32]
  wire  _GEN_12164 = _T_1530 ? _GEN_12156 : _GEN_11756; // @[sequencer-master.scala 168:32]
  wire  _GEN_12165 = _T_1530 ? _GEN_12157 : _GEN_11757; // @[sequencer-master.scala 168:32]
  wire  _GEN_12166 = _T_1530 ? _GEN_12158 : _GEN_11758; // @[sequencer-master.scala 168:32]
  wire  _GEN_12167 = _T_1530 ? _GEN_12159 : _GEN_11759; // @[sequencer-master.scala 168:32]
  wire  _GEN_12168 = _T_1530 ? _GEN_12160 : _GEN_11760; // @[sequencer-master.scala 168:32]
  wire  _GEN_12169 = _T_1530 ? _GEN_12161 : _GEN_11761; // @[sequencer-master.scala 168:32]
  wire  _GEN_12170 = _GEN_34121 | _GEN_11778; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12171 = _GEN_34122 | _GEN_11779; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12172 = _GEN_34123 | _GEN_11780; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12173 = _GEN_34124 | _GEN_11781; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12174 = _GEN_34125 | _GEN_11782; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12175 = _GEN_34126 | _GEN_11783; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12176 = _GEN_34127 | _GEN_11784; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12177 = _GEN_34128 | _GEN_11785; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12178 = _T_1552 ? _GEN_12170 : _GEN_11778; // @[sequencer-master.scala 168:32]
  wire  _GEN_12179 = _T_1552 ? _GEN_12171 : _GEN_11779; // @[sequencer-master.scala 168:32]
  wire  _GEN_12180 = _T_1552 ? _GEN_12172 : _GEN_11780; // @[sequencer-master.scala 168:32]
  wire  _GEN_12181 = _T_1552 ? _GEN_12173 : _GEN_11781; // @[sequencer-master.scala 168:32]
  wire  _GEN_12182 = _T_1552 ? _GEN_12174 : _GEN_11782; // @[sequencer-master.scala 168:32]
  wire  _GEN_12183 = _T_1552 ? _GEN_12175 : _GEN_11783; // @[sequencer-master.scala 168:32]
  wire  _GEN_12184 = _T_1552 ? _GEN_12176 : _GEN_11784; // @[sequencer-master.scala 168:32]
  wire  _GEN_12185 = _T_1552 ? _GEN_12177 : _GEN_11785; // @[sequencer-master.scala 168:32]
  wire  _GEN_12186 = _GEN_34121 | _GEN_11802; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12187 = _GEN_34122 | _GEN_11803; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12188 = _GEN_34123 | _GEN_11804; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12189 = _GEN_34124 | _GEN_11805; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12190 = _GEN_34125 | _GEN_11806; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12191 = _GEN_34126 | _GEN_11807; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12192 = _GEN_34127 | _GEN_11808; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12193 = _GEN_34128 | _GEN_11809; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12194 = _T_1574 ? _GEN_12186 : _GEN_11802; // @[sequencer-master.scala 168:32]
  wire  _GEN_12195 = _T_1574 ? _GEN_12187 : _GEN_11803; // @[sequencer-master.scala 168:32]
  wire  _GEN_12196 = _T_1574 ? _GEN_12188 : _GEN_11804; // @[sequencer-master.scala 168:32]
  wire  _GEN_12197 = _T_1574 ? _GEN_12189 : _GEN_11805; // @[sequencer-master.scala 168:32]
  wire  _GEN_12198 = _T_1574 ? _GEN_12190 : _GEN_11806; // @[sequencer-master.scala 168:32]
  wire  _GEN_12199 = _T_1574 ? _GEN_12191 : _GEN_11807; // @[sequencer-master.scala 168:32]
  wire  _GEN_12200 = _T_1574 ? _GEN_12192 : _GEN_11808; // @[sequencer-master.scala 168:32]
  wire  _GEN_12201 = _T_1574 ? _GEN_12193 : _GEN_11809; // @[sequencer-master.scala 168:32]
  wire  _GEN_12202 = _GEN_34121 | _GEN_11826; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12203 = _GEN_34122 | _GEN_11827; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12204 = _GEN_34123 | _GEN_11828; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12205 = _GEN_34124 | _GEN_11829; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12206 = _GEN_34125 | _GEN_11830; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12207 = _GEN_34126 | _GEN_11831; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12208 = _GEN_34127 | _GEN_11832; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12209 = _GEN_34128 | _GEN_11833; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_12210 = _T_1596 ? _GEN_12202 : _GEN_11826; // @[sequencer-master.scala 168:32]
  wire  _GEN_12211 = _T_1596 ? _GEN_12203 : _GEN_11827; // @[sequencer-master.scala 168:32]
  wire  _GEN_12212 = _T_1596 ? _GEN_12204 : _GEN_11828; // @[sequencer-master.scala 168:32]
  wire  _GEN_12213 = _T_1596 ? _GEN_12205 : _GEN_11829; // @[sequencer-master.scala 168:32]
  wire  _GEN_12214 = _T_1596 ? _GEN_12206 : _GEN_11830; // @[sequencer-master.scala 168:32]
  wire  _GEN_12215 = _T_1596 ? _GEN_12207 : _GEN_11831; // @[sequencer-master.scala 168:32]
  wire  _GEN_12216 = _T_1596 ? _GEN_12208 : _GEN_11832; // @[sequencer-master.scala 168:32]
  wire  _GEN_12217 = _T_1596 ? _GEN_12209 : _GEN_11833; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_12218 = 3'h0 == _T_1645 ? 2'h0 : _GEN_11298; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12219 = 3'h1 == _T_1645 ? 2'h0 : _GEN_11299; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12220 = 3'h2 == _T_1645 ? 2'h0 : _GEN_11300; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12221 = 3'h3 == _T_1645 ? 2'h0 : _GEN_11301; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12222 = 3'h4 == _T_1645 ? 2'h0 : _GEN_11302; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12223 = 3'h5 == _T_1645 ? 2'h0 : _GEN_11303; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12224 = 3'h6 == _T_1645 ? 2'h0 : _GEN_11304; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_12225 = 3'h7 == _T_1645 ? 2'h0 : _GEN_11305; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_12226 = 3'h0 == _T_1645 ? 4'h0 : _GEN_11306; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12227 = 3'h1 == _T_1645 ? 4'h0 : _GEN_11307; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12228 = 3'h2 == _T_1645 ? 4'h0 : _GEN_11308; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12229 = 3'h3 == _T_1645 ? 4'h0 : _GEN_11309; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12230 = 3'h4 == _T_1645 ? 4'h0 : _GEN_11310; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12231 = 3'h5 == _T_1645 ? 4'h0 : _GEN_11311; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12232 = 3'h6 == _T_1645 ? 4'h0 : _GEN_11312; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_12233 = 3'h7 == _T_1645 ? 4'h0 : _GEN_11313; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_12234 = 3'h0 == _T_1645 ? 3'h0 : _GEN_11314; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12235 = 3'h1 == _T_1645 ? 3'h0 : _GEN_11315; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12236 = 3'h2 == _T_1645 ? 3'h0 : _GEN_11316; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12237 = 3'h3 == _T_1645 ? 3'h0 : _GEN_11317; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12238 = 3'h4 == _T_1645 ? 3'h0 : _GEN_11318; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12239 = 3'h5 == _T_1645 ? 3'h0 : _GEN_11319; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12240 = 3'h6 == _T_1645 ? 3'h0 : _GEN_11320; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_12241 = 3'h7 == _T_1645 ? 3'h0 : _GEN_11321; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_12242 = io_op_bits_active_vfdiv ? _GEN_11578 : _GEN_9776; // @[sequencer-master.scala 645:40]
  wire  _GEN_12243 = io_op_bits_active_vfdiv ? _GEN_11579 : _GEN_9777; // @[sequencer-master.scala 645:40]
  wire  _GEN_12244 = io_op_bits_active_vfdiv ? _GEN_11580 : _GEN_9778; // @[sequencer-master.scala 645:40]
  wire  _GEN_12245 = io_op_bits_active_vfdiv ? _GEN_11581 : _GEN_9779; // @[sequencer-master.scala 645:40]
  wire  _GEN_12246 = io_op_bits_active_vfdiv ? _GEN_11582 : _GEN_9780; // @[sequencer-master.scala 645:40]
  wire  _GEN_12247 = io_op_bits_active_vfdiv ? _GEN_11583 : _GEN_9781; // @[sequencer-master.scala 645:40]
  wire  _GEN_12248 = io_op_bits_active_vfdiv ? _GEN_11584 : _GEN_9782; // @[sequencer-master.scala 645:40]
  wire  _GEN_12249 = io_op_bits_active_vfdiv ? _GEN_11585 : _GEN_9783; // @[sequencer-master.scala 645:40]
  wire  _GEN_12258 = io_op_bits_active_vfdiv ? _GEN_11594 : _GEN_9792; // @[sequencer-master.scala 645:40]
  wire  _GEN_12259 = io_op_bits_active_vfdiv ? _GEN_11595 : _GEN_9793; // @[sequencer-master.scala 645:40]
  wire  _GEN_12260 = io_op_bits_active_vfdiv ? _GEN_11596 : _GEN_9794; // @[sequencer-master.scala 645:40]
  wire  _GEN_12261 = io_op_bits_active_vfdiv ? _GEN_11597 : _GEN_9795; // @[sequencer-master.scala 645:40]
  wire  _GEN_12262 = io_op_bits_active_vfdiv ? _GEN_11598 : _GEN_9796; // @[sequencer-master.scala 645:40]
  wire  _GEN_12263 = io_op_bits_active_vfdiv ? _GEN_11599 : _GEN_9797; // @[sequencer-master.scala 645:40]
  wire  _GEN_12264 = io_op_bits_active_vfdiv ? _GEN_11600 : _GEN_9798; // @[sequencer-master.scala 645:40]
  wire  _GEN_12265 = io_op_bits_active_vfdiv ? _GEN_11601 : _GEN_9799; // @[sequencer-master.scala 645:40]
  wire  _GEN_12266 = io_op_bits_active_vfdiv ? _GEN_11602 : _GEN_9800; // @[sequencer-master.scala 645:40]
  wire  _GEN_12267 = io_op_bits_active_vfdiv ? _GEN_11603 : _GEN_9801; // @[sequencer-master.scala 645:40]
  wire  _GEN_12268 = io_op_bits_active_vfdiv ? _GEN_11604 : _GEN_9802; // @[sequencer-master.scala 645:40]
  wire  _GEN_12269 = io_op_bits_active_vfdiv ? _GEN_11605 : _GEN_9803; // @[sequencer-master.scala 645:40]
  wire  _GEN_12270 = io_op_bits_active_vfdiv ? _GEN_11606 : _GEN_9804; // @[sequencer-master.scala 645:40]
  wire  _GEN_12271 = io_op_bits_active_vfdiv ? _GEN_11607 : _GEN_9805; // @[sequencer-master.scala 645:40]
  wire  _GEN_12272 = io_op_bits_active_vfdiv ? _GEN_11608 : _GEN_9806; // @[sequencer-master.scala 645:40]
  wire  _GEN_12273 = io_op_bits_active_vfdiv ? _GEN_11609 : _GEN_9807; // @[sequencer-master.scala 645:40]
  wire  _GEN_12274 = io_op_bits_active_vfdiv ? _GEN_11610 : _GEN_9808; // @[sequencer-master.scala 645:40]
  wire  _GEN_12275 = io_op_bits_active_vfdiv ? _GEN_11611 : _GEN_9809; // @[sequencer-master.scala 645:40]
  wire  _GEN_12276 = io_op_bits_active_vfdiv ? _GEN_11612 : _GEN_9810; // @[sequencer-master.scala 645:40]
  wire  _GEN_12277 = io_op_bits_active_vfdiv ? _GEN_11613 : _GEN_9811; // @[sequencer-master.scala 645:40]
  wire  _GEN_12278 = io_op_bits_active_vfdiv ? _GEN_11614 : _GEN_9812; // @[sequencer-master.scala 645:40]
  wire  _GEN_12279 = io_op_bits_active_vfdiv ? _GEN_11615 : _GEN_9813; // @[sequencer-master.scala 645:40]
  wire  _GEN_12280 = io_op_bits_active_vfdiv ? _GEN_11616 : _GEN_9814; // @[sequencer-master.scala 645:40]
  wire  _GEN_12281 = io_op_bits_active_vfdiv ? _GEN_11617 : _GEN_9815; // @[sequencer-master.scala 645:40]
  wire  _GEN_12282 = io_op_bits_active_vfdiv ? _GEN_11618 : _GEN_9816; // @[sequencer-master.scala 645:40]
  wire  _GEN_12283 = io_op_bits_active_vfdiv ? _GEN_11619 : _GEN_9817; // @[sequencer-master.scala 645:40]
  wire  _GEN_12284 = io_op_bits_active_vfdiv ? _GEN_11620 : _GEN_9818; // @[sequencer-master.scala 645:40]
  wire  _GEN_12285 = io_op_bits_active_vfdiv ? _GEN_11621 : _GEN_9819; // @[sequencer-master.scala 645:40]
  wire  _GEN_12286 = io_op_bits_active_vfdiv ? _GEN_11622 : _GEN_9820; // @[sequencer-master.scala 645:40]
  wire  _GEN_12287 = io_op_bits_active_vfdiv ? _GEN_11623 : _GEN_9821; // @[sequencer-master.scala 645:40]
  wire  _GEN_12288 = io_op_bits_active_vfdiv ? _GEN_11624 : _GEN_9822; // @[sequencer-master.scala 645:40]
  wire  _GEN_12289 = io_op_bits_active_vfdiv ? _GEN_11625 : _GEN_9823; // @[sequencer-master.scala 645:40]
  wire  _GEN_12290 = io_op_bits_active_vfdiv ? _GEN_11922 : _GEN_9824; // @[sequencer-master.scala 645:40]
  wire  _GEN_12291 = io_op_bits_active_vfdiv ? _GEN_11923 : _GEN_9825; // @[sequencer-master.scala 645:40]
  wire  _GEN_12292 = io_op_bits_active_vfdiv ? _GEN_11924 : _GEN_9826; // @[sequencer-master.scala 645:40]
  wire  _GEN_12293 = io_op_bits_active_vfdiv ? _GEN_11925 : _GEN_9827; // @[sequencer-master.scala 645:40]
  wire  _GEN_12294 = io_op_bits_active_vfdiv ? _GEN_11926 : _GEN_9828; // @[sequencer-master.scala 645:40]
  wire  _GEN_12295 = io_op_bits_active_vfdiv ? _GEN_11927 : _GEN_9829; // @[sequencer-master.scala 645:40]
  wire  _GEN_12296 = io_op_bits_active_vfdiv ? _GEN_11928 : _GEN_9830; // @[sequencer-master.scala 645:40]
  wire  _GEN_12297 = io_op_bits_active_vfdiv ? _GEN_11929 : _GEN_9831; // @[sequencer-master.scala 645:40]
  wire  _GEN_12298 = io_op_bits_active_vfdiv ? _GEN_11634 : _GEN_9832; // @[sequencer-master.scala 645:40]
  wire  _GEN_12299 = io_op_bits_active_vfdiv ? _GEN_11635 : _GEN_9833; // @[sequencer-master.scala 645:40]
  wire  _GEN_12300 = io_op_bits_active_vfdiv ? _GEN_11636 : _GEN_9834; // @[sequencer-master.scala 645:40]
  wire  _GEN_12301 = io_op_bits_active_vfdiv ? _GEN_11637 : _GEN_9835; // @[sequencer-master.scala 645:40]
  wire  _GEN_12302 = io_op_bits_active_vfdiv ? _GEN_11638 : _GEN_9836; // @[sequencer-master.scala 645:40]
  wire  _GEN_12303 = io_op_bits_active_vfdiv ? _GEN_11639 : _GEN_9837; // @[sequencer-master.scala 645:40]
  wire  _GEN_12304 = io_op_bits_active_vfdiv ? _GEN_11640 : _GEN_9838; // @[sequencer-master.scala 645:40]
  wire  _GEN_12305 = io_op_bits_active_vfdiv ? _GEN_11641 : _GEN_9839; // @[sequencer-master.scala 645:40]
  wire  _GEN_12306 = io_op_bits_active_vfdiv ? _GEN_11642 : _GEN_9840; // @[sequencer-master.scala 645:40]
  wire  _GEN_12307 = io_op_bits_active_vfdiv ? _GEN_11643 : _GEN_9841; // @[sequencer-master.scala 645:40]
  wire  _GEN_12308 = io_op_bits_active_vfdiv ? _GEN_11644 : _GEN_9842; // @[sequencer-master.scala 645:40]
  wire  _GEN_12309 = io_op_bits_active_vfdiv ? _GEN_11645 : _GEN_9843; // @[sequencer-master.scala 645:40]
  wire  _GEN_12310 = io_op_bits_active_vfdiv ? _GEN_11646 : _GEN_9844; // @[sequencer-master.scala 645:40]
  wire  _GEN_12311 = io_op_bits_active_vfdiv ? _GEN_11647 : _GEN_9845; // @[sequencer-master.scala 645:40]
  wire  _GEN_12312 = io_op_bits_active_vfdiv ? _GEN_11648 : _GEN_9846; // @[sequencer-master.scala 645:40]
  wire  _GEN_12313 = io_op_bits_active_vfdiv ? _GEN_11649 : _GEN_9847; // @[sequencer-master.scala 645:40]
  wire  _GEN_12314 = io_op_bits_active_vfdiv ? _GEN_11970 : _GEN_9848; // @[sequencer-master.scala 645:40]
  wire  _GEN_12315 = io_op_bits_active_vfdiv ? _GEN_11971 : _GEN_9849; // @[sequencer-master.scala 645:40]
  wire  _GEN_12316 = io_op_bits_active_vfdiv ? _GEN_11972 : _GEN_9850; // @[sequencer-master.scala 645:40]
  wire  _GEN_12317 = io_op_bits_active_vfdiv ? _GEN_11973 : _GEN_9851; // @[sequencer-master.scala 645:40]
  wire  _GEN_12318 = io_op_bits_active_vfdiv ? _GEN_11974 : _GEN_9852; // @[sequencer-master.scala 645:40]
  wire  _GEN_12319 = io_op_bits_active_vfdiv ? _GEN_11975 : _GEN_9853; // @[sequencer-master.scala 645:40]
  wire  _GEN_12320 = io_op_bits_active_vfdiv ? _GEN_11976 : _GEN_9854; // @[sequencer-master.scala 645:40]
  wire  _GEN_12321 = io_op_bits_active_vfdiv ? _GEN_11977 : _GEN_9855; // @[sequencer-master.scala 645:40]
  wire  _GEN_12322 = io_op_bits_active_vfdiv ? _GEN_12098 : _GEN_9856; // @[sequencer-master.scala 645:40]
  wire  _GEN_12323 = io_op_bits_active_vfdiv ? _GEN_12099 : _GEN_9857; // @[sequencer-master.scala 645:40]
  wire  _GEN_12324 = io_op_bits_active_vfdiv ? _GEN_12100 : _GEN_9858; // @[sequencer-master.scala 645:40]
  wire  _GEN_12325 = io_op_bits_active_vfdiv ? _GEN_12101 : _GEN_9859; // @[sequencer-master.scala 645:40]
  wire  _GEN_12326 = io_op_bits_active_vfdiv ? _GEN_12102 : _GEN_9860; // @[sequencer-master.scala 645:40]
  wire  _GEN_12327 = io_op_bits_active_vfdiv ? _GEN_12103 : _GEN_9861; // @[sequencer-master.scala 645:40]
  wire  _GEN_12328 = io_op_bits_active_vfdiv ? _GEN_12104 : _GEN_9862; // @[sequencer-master.scala 645:40]
  wire  _GEN_12329 = io_op_bits_active_vfdiv ? _GEN_12105 : _GEN_9863; // @[sequencer-master.scala 645:40]
  wire  _GEN_12330 = io_op_bits_active_vfdiv ? _GEN_11666 : _GEN_9864; // @[sequencer-master.scala 645:40]
  wire  _GEN_12331 = io_op_bits_active_vfdiv ? _GEN_11667 : _GEN_9865; // @[sequencer-master.scala 645:40]
  wire  _GEN_12332 = io_op_bits_active_vfdiv ? _GEN_11668 : _GEN_9866; // @[sequencer-master.scala 645:40]
  wire  _GEN_12333 = io_op_bits_active_vfdiv ? _GEN_11669 : _GEN_9867; // @[sequencer-master.scala 645:40]
  wire  _GEN_12334 = io_op_bits_active_vfdiv ? _GEN_11670 : _GEN_9868; // @[sequencer-master.scala 645:40]
  wire  _GEN_12335 = io_op_bits_active_vfdiv ? _GEN_11671 : _GEN_9869; // @[sequencer-master.scala 645:40]
  wire  _GEN_12336 = io_op_bits_active_vfdiv ? _GEN_11672 : _GEN_9870; // @[sequencer-master.scala 645:40]
  wire  _GEN_12337 = io_op_bits_active_vfdiv ? _GEN_11673 : _GEN_9871; // @[sequencer-master.scala 645:40]
  wire  _GEN_12338 = io_op_bits_active_vfdiv ? _GEN_11986 : _GEN_9872; // @[sequencer-master.scala 645:40]
  wire  _GEN_12339 = io_op_bits_active_vfdiv ? _GEN_11987 : _GEN_9873; // @[sequencer-master.scala 645:40]
  wire  _GEN_12340 = io_op_bits_active_vfdiv ? _GEN_11988 : _GEN_9874; // @[sequencer-master.scala 645:40]
  wire  _GEN_12341 = io_op_bits_active_vfdiv ? _GEN_11989 : _GEN_9875; // @[sequencer-master.scala 645:40]
  wire  _GEN_12342 = io_op_bits_active_vfdiv ? _GEN_11990 : _GEN_9876; // @[sequencer-master.scala 645:40]
  wire  _GEN_12343 = io_op_bits_active_vfdiv ? _GEN_11991 : _GEN_9877; // @[sequencer-master.scala 645:40]
  wire  _GEN_12344 = io_op_bits_active_vfdiv ? _GEN_11992 : _GEN_9878; // @[sequencer-master.scala 645:40]
  wire  _GEN_12345 = io_op_bits_active_vfdiv ? _GEN_11993 : _GEN_9879; // @[sequencer-master.scala 645:40]
  wire  _GEN_12346 = io_op_bits_active_vfdiv ? _GEN_12114 : _GEN_9880; // @[sequencer-master.scala 645:40]
  wire  _GEN_12347 = io_op_bits_active_vfdiv ? _GEN_12115 : _GEN_9881; // @[sequencer-master.scala 645:40]
  wire  _GEN_12348 = io_op_bits_active_vfdiv ? _GEN_12116 : _GEN_9882; // @[sequencer-master.scala 645:40]
  wire  _GEN_12349 = io_op_bits_active_vfdiv ? _GEN_12117 : _GEN_9883; // @[sequencer-master.scala 645:40]
  wire  _GEN_12350 = io_op_bits_active_vfdiv ? _GEN_12118 : _GEN_9884; // @[sequencer-master.scala 645:40]
  wire  _GEN_12351 = io_op_bits_active_vfdiv ? _GEN_12119 : _GEN_9885; // @[sequencer-master.scala 645:40]
  wire  _GEN_12352 = io_op_bits_active_vfdiv ? _GEN_12120 : _GEN_9886; // @[sequencer-master.scala 645:40]
  wire  _GEN_12353 = io_op_bits_active_vfdiv ? _GEN_12121 : _GEN_9887; // @[sequencer-master.scala 645:40]
  wire  _GEN_12354 = io_op_bits_active_vfdiv ? _GEN_11690 : _GEN_9888; // @[sequencer-master.scala 645:40]
  wire  _GEN_12355 = io_op_bits_active_vfdiv ? _GEN_11691 : _GEN_9889; // @[sequencer-master.scala 645:40]
  wire  _GEN_12356 = io_op_bits_active_vfdiv ? _GEN_11692 : _GEN_9890; // @[sequencer-master.scala 645:40]
  wire  _GEN_12357 = io_op_bits_active_vfdiv ? _GEN_11693 : _GEN_9891; // @[sequencer-master.scala 645:40]
  wire  _GEN_12358 = io_op_bits_active_vfdiv ? _GEN_11694 : _GEN_9892; // @[sequencer-master.scala 645:40]
  wire  _GEN_12359 = io_op_bits_active_vfdiv ? _GEN_11695 : _GEN_9893; // @[sequencer-master.scala 645:40]
  wire  _GEN_12360 = io_op_bits_active_vfdiv ? _GEN_11696 : _GEN_9894; // @[sequencer-master.scala 645:40]
  wire  _GEN_12361 = io_op_bits_active_vfdiv ? _GEN_11697 : _GEN_9895; // @[sequencer-master.scala 645:40]
  wire  _GEN_12362 = io_op_bits_active_vfdiv ? _GEN_12002 : _GEN_9896; // @[sequencer-master.scala 645:40]
  wire  _GEN_12363 = io_op_bits_active_vfdiv ? _GEN_12003 : _GEN_9897; // @[sequencer-master.scala 645:40]
  wire  _GEN_12364 = io_op_bits_active_vfdiv ? _GEN_12004 : _GEN_9898; // @[sequencer-master.scala 645:40]
  wire  _GEN_12365 = io_op_bits_active_vfdiv ? _GEN_12005 : _GEN_9899; // @[sequencer-master.scala 645:40]
  wire  _GEN_12366 = io_op_bits_active_vfdiv ? _GEN_12006 : _GEN_9900; // @[sequencer-master.scala 645:40]
  wire  _GEN_12367 = io_op_bits_active_vfdiv ? _GEN_12007 : _GEN_9901; // @[sequencer-master.scala 645:40]
  wire  _GEN_12368 = io_op_bits_active_vfdiv ? _GEN_12008 : _GEN_9902; // @[sequencer-master.scala 645:40]
  wire  _GEN_12369 = io_op_bits_active_vfdiv ? _GEN_12009 : _GEN_9903; // @[sequencer-master.scala 645:40]
  wire  _GEN_12370 = io_op_bits_active_vfdiv ? _GEN_12130 : _GEN_9904; // @[sequencer-master.scala 645:40]
  wire  _GEN_12371 = io_op_bits_active_vfdiv ? _GEN_12131 : _GEN_9905; // @[sequencer-master.scala 645:40]
  wire  _GEN_12372 = io_op_bits_active_vfdiv ? _GEN_12132 : _GEN_9906; // @[sequencer-master.scala 645:40]
  wire  _GEN_12373 = io_op_bits_active_vfdiv ? _GEN_12133 : _GEN_9907; // @[sequencer-master.scala 645:40]
  wire  _GEN_12374 = io_op_bits_active_vfdiv ? _GEN_12134 : _GEN_9908; // @[sequencer-master.scala 645:40]
  wire  _GEN_12375 = io_op_bits_active_vfdiv ? _GEN_12135 : _GEN_9909; // @[sequencer-master.scala 645:40]
  wire  _GEN_12376 = io_op_bits_active_vfdiv ? _GEN_12136 : _GEN_9910; // @[sequencer-master.scala 645:40]
  wire  _GEN_12377 = io_op_bits_active_vfdiv ? _GEN_12137 : _GEN_9911; // @[sequencer-master.scala 645:40]
  wire  _GEN_12378 = io_op_bits_active_vfdiv ? _GEN_11714 : _GEN_9912; // @[sequencer-master.scala 645:40]
  wire  _GEN_12379 = io_op_bits_active_vfdiv ? _GEN_11715 : _GEN_9913; // @[sequencer-master.scala 645:40]
  wire  _GEN_12380 = io_op_bits_active_vfdiv ? _GEN_11716 : _GEN_9914; // @[sequencer-master.scala 645:40]
  wire  _GEN_12381 = io_op_bits_active_vfdiv ? _GEN_11717 : _GEN_9915; // @[sequencer-master.scala 645:40]
  wire  _GEN_12382 = io_op_bits_active_vfdiv ? _GEN_11718 : _GEN_9916; // @[sequencer-master.scala 645:40]
  wire  _GEN_12383 = io_op_bits_active_vfdiv ? _GEN_11719 : _GEN_9917; // @[sequencer-master.scala 645:40]
  wire  _GEN_12384 = io_op_bits_active_vfdiv ? _GEN_11720 : _GEN_9918; // @[sequencer-master.scala 645:40]
  wire  _GEN_12385 = io_op_bits_active_vfdiv ? _GEN_11721 : _GEN_9919; // @[sequencer-master.scala 645:40]
  wire  _GEN_12386 = io_op_bits_active_vfdiv ? _GEN_12018 : _GEN_9920; // @[sequencer-master.scala 645:40]
  wire  _GEN_12387 = io_op_bits_active_vfdiv ? _GEN_12019 : _GEN_9921; // @[sequencer-master.scala 645:40]
  wire  _GEN_12388 = io_op_bits_active_vfdiv ? _GEN_12020 : _GEN_9922; // @[sequencer-master.scala 645:40]
  wire  _GEN_12389 = io_op_bits_active_vfdiv ? _GEN_12021 : _GEN_9923; // @[sequencer-master.scala 645:40]
  wire  _GEN_12390 = io_op_bits_active_vfdiv ? _GEN_12022 : _GEN_9924; // @[sequencer-master.scala 645:40]
  wire  _GEN_12391 = io_op_bits_active_vfdiv ? _GEN_12023 : _GEN_9925; // @[sequencer-master.scala 645:40]
  wire  _GEN_12392 = io_op_bits_active_vfdiv ? _GEN_12024 : _GEN_9926; // @[sequencer-master.scala 645:40]
  wire  _GEN_12393 = io_op_bits_active_vfdiv ? _GEN_12025 : _GEN_9927; // @[sequencer-master.scala 645:40]
  wire  _GEN_12394 = io_op_bits_active_vfdiv ? _GEN_12146 : _GEN_9928; // @[sequencer-master.scala 645:40]
  wire  _GEN_12395 = io_op_bits_active_vfdiv ? _GEN_12147 : _GEN_9929; // @[sequencer-master.scala 645:40]
  wire  _GEN_12396 = io_op_bits_active_vfdiv ? _GEN_12148 : _GEN_9930; // @[sequencer-master.scala 645:40]
  wire  _GEN_12397 = io_op_bits_active_vfdiv ? _GEN_12149 : _GEN_9931; // @[sequencer-master.scala 645:40]
  wire  _GEN_12398 = io_op_bits_active_vfdiv ? _GEN_12150 : _GEN_9932; // @[sequencer-master.scala 645:40]
  wire  _GEN_12399 = io_op_bits_active_vfdiv ? _GEN_12151 : _GEN_9933; // @[sequencer-master.scala 645:40]
  wire  _GEN_12400 = io_op_bits_active_vfdiv ? _GEN_12152 : _GEN_9934; // @[sequencer-master.scala 645:40]
  wire  _GEN_12401 = io_op_bits_active_vfdiv ? _GEN_12153 : _GEN_9935; // @[sequencer-master.scala 645:40]
  wire  _GEN_12402 = io_op_bits_active_vfdiv ? _GEN_11738 : _GEN_9936; // @[sequencer-master.scala 645:40]
  wire  _GEN_12403 = io_op_bits_active_vfdiv ? _GEN_11739 : _GEN_9937; // @[sequencer-master.scala 645:40]
  wire  _GEN_12404 = io_op_bits_active_vfdiv ? _GEN_11740 : _GEN_9938; // @[sequencer-master.scala 645:40]
  wire  _GEN_12405 = io_op_bits_active_vfdiv ? _GEN_11741 : _GEN_9939; // @[sequencer-master.scala 645:40]
  wire  _GEN_12406 = io_op_bits_active_vfdiv ? _GEN_11742 : _GEN_9940; // @[sequencer-master.scala 645:40]
  wire  _GEN_12407 = io_op_bits_active_vfdiv ? _GEN_11743 : _GEN_9941; // @[sequencer-master.scala 645:40]
  wire  _GEN_12408 = io_op_bits_active_vfdiv ? _GEN_11744 : _GEN_9942; // @[sequencer-master.scala 645:40]
  wire  _GEN_12409 = io_op_bits_active_vfdiv ? _GEN_11745 : _GEN_9943; // @[sequencer-master.scala 645:40]
  wire  _GEN_12410 = io_op_bits_active_vfdiv ? _GEN_12034 : _GEN_9944; // @[sequencer-master.scala 645:40]
  wire  _GEN_12411 = io_op_bits_active_vfdiv ? _GEN_12035 : _GEN_9945; // @[sequencer-master.scala 645:40]
  wire  _GEN_12412 = io_op_bits_active_vfdiv ? _GEN_12036 : _GEN_9946; // @[sequencer-master.scala 645:40]
  wire  _GEN_12413 = io_op_bits_active_vfdiv ? _GEN_12037 : _GEN_9947; // @[sequencer-master.scala 645:40]
  wire  _GEN_12414 = io_op_bits_active_vfdiv ? _GEN_12038 : _GEN_9948; // @[sequencer-master.scala 645:40]
  wire  _GEN_12415 = io_op_bits_active_vfdiv ? _GEN_12039 : _GEN_9949; // @[sequencer-master.scala 645:40]
  wire  _GEN_12416 = io_op_bits_active_vfdiv ? _GEN_12040 : _GEN_9950; // @[sequencer-master.scala 645:40]
  wire  _GEN_12417 = io_op_bits_active_vfdiv ? _GEN_12041 : _GEN_9951; // @[sequencer-master.scala 645:40]
  wire  _GEN_12418 = io_op_bits_active_vfdiv ? _GEN_12162 : _GEN_9952; // @[sequencer-master.scala 645:40]
  wire  _GEN_12419 = io_op_bits_active_vfdiv ? _GEN_12163 : _GEN_9953; // @[sequencer-master.scala 645:40]
  wire  _GEN_12420 = io_op_bits_active_vfdiv ? _GEN_12164 : _GEN_9954; // @[sequencer-master.scala 645:40]
  wire  _GEN_12421 = io_op_bits_active_vfdiv ? _GEN_12165 : _GEN_9955; // @[sequencer-master.scala 645:40]
  wire  _GEN_12422 = io_op_bits_active_vfdiv ? _GEN_12166 : _GEN_9956; // @[sequencer-master.scala 645:40]
  wire  _GEN_12423 = io_op_bits_active_vfdiv ? _GEN_12167 : _GEN_9957; // @[sequencer-master.scala 645:40]
  wire  _GEN_12424 = io_op_bits_active_vfdiv ? _GEN_12168 : _GEN_9958; // @[sequencer-master.scala 645:40]
  wire  _GEN_12425 = io_op_bits_active_vfdiv ? _GEN_12169 : _GEN_9959; // @[sequencer-master.scala 645:40]
  wire  _GEN_12426 = io_op_bits_active_vfdiv ? _GEN_11762 : _GEN_9960; // @[sequencer-master.scala 645:40]
  wire  _GEN_12427 = io_op_bits_active_vfdiv ? _GEN_11763 : _GEN_9961; // @[sequencer-master.scala 645:40]
  wire  _GEN_12428 = io_op_bits_active_vfdiv ? _GEN_11764 : _GEN_9962; // @[sequencer-master.scala 645:40]
  wire  _GEN_12429 = io_op_bits_active_vfdiv ? _GEN_11765 : _GEN_9963; // @[sequencer-master.scala 645:40]
  wire  _GEN_12430 = io_op_bits_active_vfdiv ? _GEN_11766 : _GEN_9964; // @[sequencer-master.scala 645:40]
  wire  _GEN_12431 = io_op_bits_active_vfdiv ? _GEN_11767 : _GEN_9965; // @[sequencer-master.scala 645:40]
  wire  _GEN_12432 = io_op_bits_active_vfdiv ? _GEN_11768 : _GEN_9966; // @[sequencer-master.scala 645:40]
  wire  _GEN_12433 = io_op_bits_active_vfdiv ? _GEN_11769 : _GEN_9967; // @[sequencer-master.scala 645:40]
  wire  _GEN_12434 = io_op_bits_active_vfdiv ? _GEN_12050 : _GEN_9968; // @[sequencer-master.scala 645:40]
  wire  _GEN_12435 = io_op_bits_active_vfdiv ? _GEN_12051 : _GEN_9969; // @[sequencer-master.scala 645:40]
  wire  _GEN_12436 = io_op_bits_active_vfdiv ? _GEN_12052 : _GEN_9970; // @[sequencer-master.scala 645:40]
  wire  _GEN_12437 = io_op_bits_active_vfdiv ? _GEN_12053 : _GEN_9971; // @[sequencer-master.scala 645:40]
  wire  _GEN_12438 = io_op_bits_active_vfdiv ? _GEN_12054 : _GEN_9972; // @[sequencer-master.scala 645:40]
  wire  _GEN_12439 = io_op_bits_active_vfdiv ? _GEN_12055 : _GEN_9973; // @[sequencer-master.scala 645:40]
  wire  _GEN_12440 = io_op_bits_active_vfdiv ? _GEN_12056 : _GEN_9974; // @[sequencer-master.scala 645:40]
  wire  _GEN_12441 = io_op_bits_active_vfdiv ? _GEN_12057 : _GEN_9975; // @[sequencer-master.scala 645:40]
  wire  _GEN_12442 = io_op_bits_active_vfdiv ? _GEN_12178 : _GEN_9976; // @[sequencer-master.scala 645:40]
  wire  _GEN_12443 = io_op_bits_active_vfdiv ? _GEN_12179 : _GEN_9977; // @[sequencer-master.scala 645:40]
  wire  _GEN_12444 = io_op_bits_active_vfdiv ? _GEN_12180 : _GEN_9978; // @[sequencer-master.scala 645:40]
  wire  _GEN_12445 = io_op_bits_active_vfdiv ? _GEN_12181 : _GEN_9979; // @[sequencer-master.scala 645:40]
  wire  _GEN_12446 = io_op_bits_active_vfdiv ? _GEN_12182 : _GEN_9980; // @[sequencer-master.scala 645:40]
  wire  _GEN_12447 = io_op_bits_active_vfdiv ? _GEN_12183 : _GEN_9981; // @[sequencer-master.scala 645:40]
  wire  _GEN_12448 = io_op_bits_active_vfdiv ? _GEN_12184 : _GEN_9982; // @[sequencer-master.scala 645:40]
  wire  _GEN_12449 = io_op_bits_active_vfdiv ? _GEN_12185 : _GEN_9983; // @[sequencer-master.scala 645:40]
  wire  _GEN_12450 = io_op_bits_active_vfdiv ? _GEN_11786 : _GEN_9984; // @[sequencer-master.scala 645:40]
  wire  _GEN_12451 = io_op_bits_active_vfdiv ? _GEN_11787 : _GEN_9985; // @[sequencer-master.scala 645:40]
  wire  _GEN_12452 = io_op_bits_active_vfdiv ? _GEN_11788 : _GEN_9986; // @[sequencer-master.scala 645:40]
  wire  _GEN_12453 = io_op_bits_active_vfdiv ? _GEN_11789 : _GEN_9987; // @[sequencer-master.scala 645:40]
  wire  _GEN_12454 = io_op_bits_active_vfdiv ? _GEN_11790 : _GEN_9988; // @[sequencer-master.scala 645:40]
  wire  _GEN_12455 = io_op_bits_active_vfdiv ? _GEN_11791 : _GEN_9989; // @[sequencer-master.scala 645:40]
  wire  _GEN_12456 = io_op_bits_active_vfdiv ? _GEN_11792 : _GEN_9990; // @[sequencer-master.scala 645:40]
  wire  _GEN_12457 = io_op_bits_active_vfdiv ? _GEN_11793 : _GEN_9991; // @[sequencer-master.scala 645:40]
  wire  _GEN_12458 = io_op_bits_active_vfdiv ? _GEN_12066 : _GEN_9992; // @[sequencer-master.scala 645:40]
  wire  _GEN_12459 = io_op_bits_active_vfdiv ? _GEN_12067 : _GEN_9993; // @[sequencer-master.scala 645:40]
  wire  _GEN_12460 = io_op_bits_active_vfdiv ? _GEN_12068 : _GEN_9994; // @[sequencer-master.scala 645:40]
  wire  _GEN_12461 = io_op_bits_active_vfdiv ? _GEN_12069 : _GEN_9995; // @[sequencer-master.scala 645:40]
  wire  _GEN_12462 = io_op_bits_active_vfdiv ? _GEN_12070 : _GEN_9996; // @[sequencer-master.scala 645:40]
  wire  _GEN_12463 = io_op_bits_active_vfdiv ? _GEN_12071 : _GEN_9997; // @[sequencer-master.scala 645:40]
  wire  _GEN_12464 = io_op_bits_active_vfdiv ? _GEN_12072 : _GEN_9998; // @[sequencer-master.scala 645:40]
  wire  _GEN_12465 = io_op_bits_active_vfdiv ? _GEN_12073 : _GEN_9999; // @[sequencer-master.scala 645:40]
  wire  _GEN_12466 = io_op_bits_active_vfdiv ? _GEN_12194 : _GEN_10000; // @[sequencer-master.scala 645:40]
  wire  _GEN_12467 = io_op_bits_active_vfdiv ? _GEN_12195 : _GEN_10001; // @[sequencer-master.scala 645:40]
  wire  _GEN_12468 = io_op_bits_active_vfdiv ? _GEN_12196 : _GEN_10002; // @[sequencer-master.scala 645:40]
  wire  _GEN_12469 = io_op_bits_active_vfdiv ? _GEN_12197 : _GEN_10003; // @[sequencer-master.scala 645:40]
  wire  _GEN_12470 = io_op_bits_active_vfdiv ? _GEN_12198 : _GEN_10004; // @[sequencer-master.scala 645:40]
  wire  _GEN_12471 = io_op_bits_active_vfdiv ? _GEN_12199 : _GEN_10005; // @[sequencer-master.scala 645:40]
  wire  _GEN_12472 = io_op_bits_active_vfdiv ? _GEN_12200 : _GEN_10006; // @[sequencer-master.scala 645:40]
  wire  _GEN_12473 = io_op_bits_active_vfdiv ? _GEN_12201 : _GEN_10007; // @[sequencer-master.scala 645:40]
  wire  _GEN_12474 = io_op_bits_active_vfdiv ? _GEN_11810 : _GEN_10008; // @[sequencer-master.scala 645:40]
  wire  _GEN_12475 = io_op_bits_active_vfdiv ? _GEN_11811 : _GEN_10009; // @[sequencer-master.scala 645:40]
  wire  _GEN_12476 = io_op_bits_active_vfdiv ? _GEN_11812 : _GEN_10010; // @[sequencer-master.scala 645:40]
  wire  _GEN_12477 = io_op_bits_active_vfdiv ? _GEN_11813 : _GEN_10011; // @[sequencer-master.scala 645:40]
  wire  _GEN_12478 = io_op_bits_active_vfdiv ? _GEN_11814 : _GEN_10012; // @[sequencer-master.scala 645:40]
  wire  _GEN_12479 = io_op_bits_active_vfdiv ? _GEN_11815 : _GEN_10013; // @[sequencer-master.scala 645:40]
  wire  _GEN_12480 = io_op_bits_active_vfdiv ? _GEN_11816 : _GEN_10014; // @[sequencer-master.scala 645:40]
  wire  _GEN_12481 = io_op_bits_active_vfdiv ? _GEN_11817 : _GEN_10015; // @[sequencer-master.scala 645:40]
  wire  _GEN_12482 = io_op_bits_active_vfdiv ? _GEN_12082 : _GEN_10016; // @[sequencer-master.scala 645:40]
  wire  _GEN_12483 = io_op_bits_active_vfdiv ? _GEN_12083 : _GEN_10017; // @[sequencer-master.scala 645:40]
  wire  _GEN_12484 = io_op_bits_active_vfdiv ? _GEN_12084 : _GEN_10018; // @[sequencer-master.scala 645:40]
  wire  _GEN_12485 = io_op_bits_active_vfdiv ? _GEN_12085 : _GEN_10019; // @[sequencer-master.scala 645:40]
  wire  _GEN_12486 = io_op_bits_active_vfdiv ? _GEN_12086 : _GEN_10020; // @[sequencer-master.scala 645:40]
  wire  _GEN_12487 = io_op_bits_active_vfdiv ? _GEN_12087 : _GEN_10021; // @[sequencer-master.scala 645:40]
  wire  _GEN_12488 = io_op_bits_active_vfdiv ? _GEN_12088 : _GEN_10022; // @[sequencer-master.scala 645:40]
  wire  _GEN_12489 = io_op_bits_active_vfdiv ? _GEN_12089 : _GEN_10023; // @[sequencer-master.scala 645:40]
  wire  _GEN_12490 = io_op_bits_active_vfdiv ? _GEN_12210 : _GEN_10024; // @[sequencer-master.scala 645:40]
  wire  _GEN_12491 = io_op_bits_active_vfdiv ? _GEN_12211 : _GEN_10025; // @[sequencer-master.scala 645:40]
  wire  _GEN_12492 = io_op_bits_active_vfdiv ? _GEN_12212 : _GEN_10026; // @[sequencer-master.scala 645:40]
  wire  _GEN_12493 = io_op_bits_active_vfdiv ? _GEN_12213 : _GEN_10027; // @[sequencer-master.scala 645:40]
  wire  _GEN_12494 = io_op_bits_active_vfdiv ? _GEN_12214 : _GEN_10028; // @[sequencer-master.scala 645:40]
  wire  _GEN_12495 = io_op_bits_active_vfdiv ? _GEN_12215 : _GEN_10029; // @[sequencer-master.scala 645:40]
  wire  _GEN_12496 = io_op_bits_active_vfdiv ? _GEN_12216 : _GEN_10030; // @[sequencer-master.scala 645:40]
  wire  _GEN_12497 = io_op_bits_active_vfdiv ? _GEN_12217 : _GEN_10031; // @[sequencer-master.scala 645:40]
  wire  _GEN_12498 = io_op_bits_active_vfdiv ? _GEN_11834 : _GEN_10032; // @[sequencer-master.scala 645:40]
  wire  _GEN_12499 = io_op_bits_active_vfdiv ? _GEN_11835 : _GEN_10033; // @[sequencer-master.scala 645:40]
  wire  _GEN_12500 = io_op_bits_active_vfdiv ? _GEN_11836 : _GEN_10034; // @[sequencer-master.scala 645:40]
  wire  _GEN_12501 = io_op_bits_active_vfdiv ? _GEN_11837 : _GEN_10035; // @[sequencer-master.scala 645:40]
  wire  _GEN_12502 = io_op_bits_active_vfdiv ? _GEN_11838 : _GEN_10036; // @[sequencer-master.scala 645:40]
  wire  _GEN_12503 = io_op_bits_active_vfdiv ? _GEN_11839 : _GEN_10037; // @[sequencer-master.scala 645:40]
  wire  _GEN_12504 = io_op_bits_active_vfdiv ? _GEN_11840 : _GEN_10038; // @[sequencer-master.scala 645:40]
  wire  _GEN_12505 = io_op_bits_active_vfdiv ? _GEN_11841 : _GEN_10039; // @[sequencer-master.scala 645:40]
  wire  _GEN_12514 = io_op_bits_active_vfdiv ? _GEN_10578 : _GEN_7910; // @[sequencer-master.scala 645:40]
  wire  _GEN_12515 = io_op_bits_active_vfdiv ? _GEN_10579 : _GEN_7911; // @[sequencer-master.scala 645:40]
  wire  _GEN_12516 = io_op_bits_active_vfdiv ? _GEN_10580 : _GEN_7912; // @[sequencer-master.scala 645:40]
  wire  _GEN_12517 = io_op_bits_active_vfdiv ? _GEN_10581 : _GEN_7913; // @[sequencer-master.scala 645:40]
  wire  _GEN_12518 = io_op_bits_active_vfdiv ? _GEN_10582 : _GEN_7914; // @[sequencer-master.scala 645:40]
  wire  _GEN_12519 = io_op_bits_active_vfdiv ? _GEN_10583 : _GEN_7915; // @[sequencer-master.scala 645:40]
  wire  _GEN_12520 = io_op_bits_active_vfdiv ? _GEN_10584 : _GEN_7916; // @[sequencer-master.scala 645:40]
  wire  _GEN_12521 = io_op_bits_active_vfdiv ? _GEN_10585 : _GEN_7917; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12522 = io_op_bits_active_vfdiv ? _GEN_11858 : _GEN_10056; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12523 = io_op_bits_active_vfdiv ? _GEN_11859 : _GEN_10057; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12524 = io_op_bits_active_vfdiv ? _GEN_11860 : _GEN_10058; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12525 = io_op_bits_active_vfdiv ? _GEN_11861 : _GEN_10059; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12526 = io_op_bits_active_vfdiv ? _GEN_11862 : _GEN_10060; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12527 = io_op_bits_active_vfdiv ? _GEN_11863 : _GEN_10061; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12528 = io_op_bits_active_vfdiv ? _GEN_11864 : _GEN_10062; // @[sequencer-master.scala 645:40]
  wire [9:0] _GEN_12529 = io_op_bits_active_vfdiv ? _GEN_11865 : _GEN_10063; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12530 = io_op_bits_active_vfdiv ? _GEN_10634 : _GEN_10064; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12531 = io_op_bits_active_vfdiv ? _GEN_10635 : _GEN_10065; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12532 = io_op_bits_active_vfdiv ? _GEN_10636 : _GEN_10066; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12533 = io_op_bits_active_vfdiv ? _GEN_10637 : _GEN_10067; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12534 = io_op_bits_active_vfdiv ? _GEN_10638 : _GEN_10068; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12535 = io_op_bits_active_vfdiv ? _GEN_10639 : _GEN_10069; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12536 = io_op_bits_active_vfdiv ? _GEN_10640 : _GEN_10070; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12537 = io_op_bits_active_vfdiv ? _GEN_10641 : _GEN_10071; // @[sequencer-master.scala 645:40]
  wire  _GEN_12538 = io_op_bits_active_vfdiv ? _GEN_10650 : _GEN_10072; // @[sequencer-master.scala 645:40]
  wire  _GEN_12539 = io_op_bits_active_vfdiv ? _GEN_10651 : _GEN_10073; // @[sequencer-master.scala 645:40]
  wire  _GEN_12540 = io_op_bits_active_vfdiv ? _GEN_10652 : _GEN_10074; // @[sequencer-master.scala 645:40]
  wire  _GEN_12541 = io_op_bits_active_vfdiv ? _GEN_10653 : _GEN_10075; // @[sequencer-master.scala 645:40]
  wire  _GEN_12542 = io_op_bits_active_vfdiv ? _GEN_10654 : _GEN_10076; // @[sequencer-master.scala 645:40]
  wire  _GEN_12543 = io_op_bits_active_vfdiv ? _GEN_10655 : _GEN_10077; // @[sequencer-master.scala 645:40]
  wire  _GEN_12544 = io_op_bits_active_vfdiv ? _GEN_10656 : _GEN_10078; // @[sequencer-master.scala 645:40]
  wire  _GEN_12545 = io_op_bits_active_vfdiv ? _GEN_10657 : _GEN_10079; // @[sequencer-master.scala 645:40]
  wire  _GEN_12546 = io_op_bits_active_vfdiv ? _GEN_10658 : _GEN_10080; // @[sequencer-master.scala 645:40]
  wire  _GEN_12547 = io_op_bits_active_vfdiv ? _GEN_10659 : _GEN_10081; // @[sequencer-master.scala 645:40]
  wire  _GEN_12548 = io_op_bits_active_vfdiv ? _GEN_10660 : _GEN_10082; // @[sequencer-master.scala 645:40]
  wire  _GEN_12549 = io_op_bits_active_vfdiv ? _GEN_10661 : _GEN_10083; // @[sequencer-master.scala 645:40]
  wire  _GEN_12550 = io_op_bits_active_vfdiv ? _GEN_10662 : _GEN_10084; // @[sequencer-master.scala 645:40]
  wire  _GEN_12551 = io_op_bits_active_vfdiv ? _GEN_10663 : _GEN_10085; // @[sequencer-master.scala 645:40]
  wire  _GEN_12552 = io_op_bits_active_vfdiv ? _GEN_10664 : _GEN_10086; // @[sequencer-master.scala 645:40]
  wire  _GEN_12553 = io_op_bits_active_vfdiv ? _GEN_10665 : _GEN_10087; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12554 = io_op_bits_active_vfdiv ? _GEN_10666 : _GEN_10088; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12555 = io_op_bits_active_vfdiv ? _GEN_10667 : _GEN_10089; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12556 = io_op_bits_active_vfdiv ? _GEN_10668 : _GEN_10090; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12557 = io_op_bits_active_vfdiv ? _GEN_10669 : _GEN_10091; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12558 = io_op_bits_active_vfdiv ? _GEN_10670 : _GEN_10092; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12559 = io_op_bits_active_vfdiv ? _GEN_10671 : _GEN_10093; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12560 = io_op_bits_active_vfdiv ? _GEN_10672 : _GEN_10094; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12561 = io_op_bits_active_vfdiv ? _GEN_10673 : _GEN_10095; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12562 = io_op_bits_active_vfdiv ? _GEN_10866 : _GEN_10096; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12563 = io_op_bits_active_vfdiv ? _GEN_10867 : _GEN_10097; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12564 = io_op_bits_active_vfdiv ? _GEN_10868 : _GEN_10098; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12565 = io_op_bits_active_vfdiv ? _GEN_10869 : _GEN_10099; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12566 = io_op_bits_active_vfdiv ? _GEN_10870 : _GEN_10100; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12567 = io_op_bits_active_vfdiv ? _GEN_10871 : _GEN_10101; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12568 = io_op_bits_active_vfdiv ? _GEN_10872 : _GEN_10102; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12569 = io_op_bits_active_vfdiv ? _GEN_10873 : _GEN_10103; // @[sequencer-master.scala 645:40]
  wire  _GEN_12570 = io_op_bits_active_vfdiv ? _GEN_10882 : _GEN_10104; // @[sequencer-master.scala 645:40]
  wire  _GEN_12571 = io_op_bits_active_vfdiv ? _GEN_10883 : _GEN_10105; // @[sequencer-master.scala 645:40]
  wire  _GEN_12572 = io_op_bits_active_vfdiv ? _GEN_10884 : _GEN_10106; // @[sequencer-master.scala 645:40]
  wire  _GEN_12573 = io_op_bits_active_vfdiv ? _GEN_10885 : _GEN_10107; // @[sequencer-master.scala 645:40]
  wire  _GEN_12574 = io_op_bits_active_vfdiv ? _GEN_10886 : _GEN_10108; // @[sequencer-master.scala 645:40]
  wire  _GEN_12575 = io_op_bits_active_vfdiv ? _GEN_10887 : _GEN_10109; // @[sequencer-master.scala 645:40]
  wire  _GEN_12576 = io_op_bits_active_vfdiv ? _GEN_10888 : _GEN_10110; // @[sequencer-master.scala 645:40]
  wire  _GEN_12577 = io_op_bits_active_vfdiv ? _GEN_10889 : _GEN_10111; // @[sequencer-master.scala 645:40]
  wire  _GEN_12578 = io_op_bits_active_vfdiv ? _GEN_10890 : _GEN_10112; // @[sequencer-master.scala 645:40]
  wire  _GEN_12579 = io_op_bits_active_vfdiv ? _GEN_10891 : _GEN_10113; // @[sequencer-master.scala 645:40]
  wire  _GEN_12580 = io_op_bits_active_vfdiv ? _GEN_10892 : _GEN_10114; // @[sequencer-master.scala 645:40]
  wire  _GEN_12581 = io_op_bits_active_vfdiv ? _GEN_10893 : _GEN_10115; // @[sequencer-master.scala 645:40]
  wire  _GEN_12582 = io_op_bits_active_vfdiv ? _GEN_10894 : _GEN_10116; // @[sequencer-master.scala 645:40]
  wire  _GEN_12583 = io_op_bits_active_vfdiv ? _GEN_10895 : _GEN_10117; // @[sequencer-master.scala 645:40]
  wire  _GEN_12584 = io_op_bits_active_vfdiv ? _GEN_10896 : _GEN_10118; // @[sequencer-master.scala 645:40]
  wire  _GEN_12585 = io_op_bits_active_vfdiv ? _GEN_10897 : _GEN_10119; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12586 = io_op_bits_active_vfdiv ? _GEN_10898 : _GEN_10120; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12587 = io_op_bits_active_vfdiv ? _GEN_10899 : _GEN_10121; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12588 = io_op_bits_active_vfdiv ? _GEN_10900 : _GEN_10122; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12589 = io_op_bits_active_vfdiv ? _GEN_10901 : _GEN_10123; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12590 = io_op_bits_active_vfdiv ? _GEN_10902 : _GEN_10124; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12591 = io_op_bits_active_vfdiv ? _GEN_10903 : _GEN_10125; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12592 = io_op_bits_active_vfdiv ? _GEN_10904 : _GEN_10126; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12593 = io_op_bits_active_vfdiv ? _GEN_10905 : _GEN_10127; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12594 = io_op_bits_active_vfdiv ? _GEN_10906 : _GEN_10128; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12595 = io_op_bits_active_vfdiv ? _GEN_10907 : _GEN_10129; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12596 = io_op_bits_active_vfdiv ? _GEN_10908 : _GEN_10130; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12597 = io_op_bits_active_vfdiv ? _GEN_10909 : _GEN_10131; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12598 = io_op_bits_active_vfdiv ? _GEN_10910 : _GEN_10132; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12599 = io_op_bits_active_vfdiv ? _GEN_10911 : _GEN_10133; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12600 = io_op_bits_active_vfdiv ? _GEN_10912 : _GEN_10134; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12601 = io_op_bits_active_vfdiv ? _GEN_10913 : _GEN_10135; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12602 = io_op_bits_active_vfdiv ? _GEN_10914 : _GEN_10136; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12603 = io_op_bits_active_vfdiv ? _GEN_10915 : _GEN_10137; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12604 = io_op_bits_active_vfdiv ? _GEN_10916 : _GEN_10138; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12605 = io_op_bits_active_vfdiv ? _GEN_10917 : _GEN_10139; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12606 = io_op_bits_active_vfdiv ? _GEN_10918 : _GEN_10140; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12607 = io_op_bits_active_vfdiv ? _GEN_10919 : _GEN_10141; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12608 = io_op_bits_active_vfdiv ? _GEN_10920 : _GEN_10142; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12609 = io_op_bits_active_vfdiv ? _GEN_10921 : _GEN_10143; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12610 = io_op_bits_active_vfdiv ? _GEN_11114 : _GEN_10144; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12611 = io_op_bits_active_vfdiv ? _GEN_11115 : _GEN_10145; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12612 = io_op_bits_active_vfdiv ? _GEN_11116 : _GEN_10146; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12613 = io_op_bits_active_vfdiv ? _GEN_11117 : _GEN_10147; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12614 = io_op_bits_active_vfdiv ? _GEN_11118 : _GEN_10148; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12615 = io_op_bits_active_vfdiv ? _GEN_11119 : _GEN_10149; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12616 = io_op_bits_active_vfdiv ? _GEN_11120 : _GEN_10150; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12617 = io_op_bits_active_vfdiv ? _GEN_11121 : _GEN_10151; // @[sequencer-master.scala 645:40]
  wire  _GEN_12618 = io_op_bits_active_vfdiv ? _GEN_11130 : _GEN_10152; // @[sequencer-master.scala 645:40]
  wire  _GEN_12619 = io_op_bits_active_vfdiv ? _GEN_11131 : _GEN_10153; // @[sequencer-master.scala 645:40]
  wire  _GEN_12620 = io_op_bits_active_vfdiv ? _GEN_11132 : _GEN_10154; // @[sequencer-master.scala 645:40]
  wire  _GEN_12621 = io_op_bits_active_vfdiv ? _GEN_11133 : _GEN_10155; // @[sequencer-master.scala 645:40]
  wire  _GEN_12622 = io_op_bits_active_vfdiv ? _GEN_11134 : _GEN_10156; // @[sequencer-master.scala 645:40]
  wire  _GEN_12623 = io_op_bits_active_vfdiv ? _GEN_11135 : _GEN_10157; // @[sequencer-master.scala 645:40]
  wire  _GEN_12624 = io_op_bits_active_vfdiv ? _GEN_11136 : _GEN_10158; // @[sequencer-master.scala 645:40]
  wire  _GEN_12625 = io_op_bits_active_vfdiv ? _GEN_11137 : _GEN_10159; // @[sequencer-master.scala 645:40]
  wire  _GEN_12626 = io_op_bits_active_vfdiv ? _GEN_11138 : _GEN_10160; // @[sequencer-master.scala 645:40]
  wire  _GEN_12627 = io_op_bits_active_vfdiv ? _GEN_11139 : _GEN_10161; // @[sequencer-master.scala 645:40]
  wire  _GEN_12628 = io_op_bits_active_vfdiv ? _GEN_11140 : _GEN_10162; // @[sequencer-master.scala 645:40]
  wire  _GEN_12629 = io_op_bits_active_vfdiv ? _GEN_11141 : _GEN_10163; // @[sequencer-master.scala 645:40]
  wire  _GEN_12630 = io_op_bits_active_vfdiv ? _GEN_11142 : _GEN_10164; // @[sequencer-master.scala 645:40]
  wire  _GEN_12631 = io_op_bits_active_vfdiv ? _GEN_11143 : _GEN_10165; // @[sequencer-master.scala 645:40]
  wire  _GEN_12632 = io_op_bits_active_vfdiv ? _GEN_11144 : _GEN_10166; // @[sequencer-master.scala 645:40]
  wire  _GEN_12633 = io_op_bits_active_vfdiv ? _GEN_11145 : _GEN_10167; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12634 = io_op_bits_active_vfdiv ? _GEN_11146 : _GEN_10168; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12635 = io_op_bits_active_vfdiv ? _GEN_11147 : _GEN_10169; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12636 = io_op_bits_active_vfdiv ? _GEN_11148 : _GEN_10170; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12637 = io_op_bits_active_vfdiv ? _GEN_11149 : _GEN_10171; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12638 = io_op_bits_active_vfdiv ? _GEN_11150 : _GEN_10172; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12639 = io_op_bits_active_vfdiv ? _GEN_11151 : _GEN_10173; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12640 = io_op_bits_active_vfdiv ? _GEN_11152 : _GEN_10174; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12641 = io_op_bits_active_vfdiv ? _GEN_11153 : _GEN_10175; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12642 = io_op_bits_active_vfdiv ? _GEN_11154 : _GEN_10176; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12643 = io_op_bits_active_vfdiv ? _GEN_11155 : _GEN_10177; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12644 = io_op_bits_active_vfdiv ? _GEN_11156 : _GEN_10178; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12645 = io_op_bits_active_vfdiv ? _GEN_11157 : _GEN_10179; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12646 = io_op_bits_active_vfdiv ? _GEN_11158 : _GEN_10180; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12647 = io_op_bits_active_vfdiv ? _GEN_11159 : _GEN_10181; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12648 = io_op_bits_active_vfdiv ? _GEN_11160 : _GEN_10182; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12649 = io_op_bits_active_vfdiv ? _GEN_11161 : _GEN_10183; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12650 = io_op_bits_active_vfdiv ? _GEN_11162 : _GEN_10184; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12651 = io_op_bits_active_vfdiv ? _GEN_11163 : _GEN_10185; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12652 = io_op_bits_active_vfdiv ? _GEN_11164 : _GEN_10186; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12653 = io_op_bits_active_vfdiv ? _GEN_11165 : _GEN_10187; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12654 = io_op_bits_active_vfdiv ? _GEN_11166 : _GEN_10188; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12655 = io_op_bits_active_vfdiv ? _GEN_11167 : _GEN_10189; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12656 = io_op_bits_active_vfdiv ? _GEN_11168 : _GEN_10190; // @[sequencer-master.scala 645:40]
  wire [63:0] _GEN_12657 = io_op_bits_active_vfdiv ? _GEN_11169 : _GEN_10191; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12658 = io_op_bits_active_vfdiv ? _GEN_12218 : _GEN_10280; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12659 = io_op_bits_active_vfdiv ? _GEN_12219 : _GEN_10281; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12660 = io_op_bits_active_vfdiv ? _GEN_12220 : _GEN_10282; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12661 = io_op_bits_active_vfdiv ? _GEN_12221 : _GEN_10283; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12662 = io_op_bits_active_vfdiv ? _GEN_12222 : _GEN_10284; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12663 = io_op_bits_active_vfdiv ? _GEN_12223 : _GEN_10285; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12664 = io_op_bits_active_vfdiv ? _GEN_12224 : _GEN_10286; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12665 = io_op_bits_active_vfdiv ? _GEN_12225 : _GEN_10287; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12666 = io_op_bits_active_vfdiv ? _GEN_12226 : _GEN_10288; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12667 = io_op_bits_active_vfdiv ? _GEN_12227 : _GEN_10289; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12668 = io_op_bits_active_vfdiv ? _GEN_12228 : _GEN_10290; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12669 = io_op_bits_active_vfdiv ? _GEN_12229 : _GEN_10291; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12670 = io_op_bits_active_vfdiv ? _GEN_12230 : _GEN_10292; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12671 = io_op_bits_active_vfdiv ? _GEN_12231 : _GEN_10293; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12672 = io_op_bits_active_vfdiv ? _GEN_12232 : _GEN_10294; // @[sequencer-master.scala 645:40]
  wire [3:0] _GEN_12673 = io_op_bits_active_vfdiv ? _GEN_12233 : _GEN_10295; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12674 = io_op_bits_active_vfdiv ? _GEN_12234 : _GEN_10296; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12675 = io_op_bits_active_vfdiv ? _GEN_12235 : _GEN_10297; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12676 = io_op_bits_active_vfdiv ? _GEN_12236 : _GEN_10298; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12677 = io_op_bits_active_vfdiv ? _GEN_12237 : _GEN_10299; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12678 = io_op_bits_active_vfdiv ? _GEN_12238 : _GEN_10300; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12679 = io_op_bits_active_vfdiv ? _GEN_12239 : _GEN_10301; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12680 = io_op_bits_active_vfdiv ? _GEN_12240 : _GEN_10302; // @[sequencer-master.scala 645:40]
  wire [2:0] _GEN_12681 = io_op_bits_active_vfdiv ? _GEN_12241 : _GEN_10303; // @[sequencer-master.scala 645:40]
  wire  _GEN_12682 = io_op_bits_active_vfdiv ? _GEN_11850 : e_0_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12683 = io_op_bits_active_vfdiv ? _GEN_11851 : e_1_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12684 = io_op_bits_active_vfdiv ? _GEN_11852 : e_2_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12685 = io_op_bits_active_vfdiv ? _GEN_11853 : e_3_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12686 = io_op_bits_active_vfdiv ? _GEN_11854 : e_4_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12687 = io_op_bits_active_vfdiv ? _GEN_11855 : e_5_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12688 = io_op_bits_active_vfdiv ? _GEN_11856 : e_6_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire  _GEN_12689 = io_op_bits_active_vfdiv ? _GEN_11857 : e_7_active_vfdu; // @[sequencer-master.scala 645:40 sequencer-master.scala 109:14]
  wire [7:0] _GEN_12690 = io_op_bits_active_vfdiv ? _GEN_11914 : _GEN_10240; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12691 = io_op_bits_active_vfdiv ? _GEN_11915 : _GEN_10241; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12692 = io_op_bits_active_vfdiv ? _GEN_11916 : _GEN_10242; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12693 = io_op_bits_active_vfdiv ? _GEN_11917 : _GEN_10243; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12694 = io_op_bits_active_vfdiv ? _GEN_11918 : _GEN_10244; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12695 = io_op_bits_active_vfdiv ? _GEN_11919 : _GEN_10245; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12696 = io_op_bits_active_vfdiv ? _GEN_11920 : _GEN_10246; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12697 = io_op_bits_active_vfdiv ? _GEN_11921 : _GEN_10247; // @[sequencer-master.scala 645:40]
  wire  _GEN_12698 = io_op_bits_active_vfdiv ? _GEN_11930 : _GEN_10248; // @[sequencer-master.scala 645:40]
  wire  _GEN_12699 = io_op_bits_active_vfdiv ? _GEN_11931 : _GEN_10249; // @[sequencer-master.scala 645:40]
  wire  _GEN_12700 = io_op_bits_active_vfdiv ? _GEN_11932 : _GEN_10250; // @[sequencer-master.scala 645:40]
  wire  _GEN_12701 = io_op_bits_active_vfdiv ? _GEN_11933 : _GEN_10251; // @[sequencer-master.scala 645:40]
  wire  _GEN_12702 = io_op_bits_active_vfdiv ? _GEN_11934 : _GEN_10252; // @[sequencer-master.scala 645:40]
  wire  _GEN_12703 = io_op_bits_active_vfdiv ? _GEN_11935 : _GEN_10253; // @[sequencer-master.scala 645:40]
  wire  _GEN_12704 = io_op_bits_active_vfdiv ? _GEN_11936 : _GEN_10254; // @[sequencer-master.scala 645:40]
  wire  _GEN_12705 = io_op_bits_active_vfdiv ? _GEN_11937 : _GEN_10255; // @[sequencer-master.scala 645:40]
  wire  _GEN_12706 = io_op_bits_active_vfdiv ? _GEN_11938 : _GEN_10256; // @[sequencer-master.scala 645:40]
  wire  _GEN_12707 = io_op_bits_active_vfdiv ? _GEN_11939 : _GEN_10257; // @[sequencer-master.scala 645:40]
  wire  _GEN_12708 = io_op_bits_active_vfdiv ? _GEN_11940 : _GEN_10258; // @[sequencer-master.scala 645:40]
  wire  _GEN_12709 = io_op_bits_active_vfdiv ? _GEN_11941 : _GEN_10259; // @[sequencer-master.scala 645:40]
  wire  _GEN_12710 = io_op_bits_active_vfdiv ? _GEN_11942 : _GEN_10260; // @[sequencer-master.scala 645:40]
  wire  _GEN_12711 = io_op_bits_active_vfdiv ? _GEN_11943 : _GEN_10261; // @[sequencer-master.scala 645:40]
  wire  _GEN_12712 = io_op_bits_active_vfdiv ? _GEN_11944 : _GEN_10262; // @[sequencer-master.scala 645:40]
  wire  _GEN_12713 = io_op_bits_active_vfdiv ? _GEN_11945 : _GEN_10263; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12714 = io_op_bits_active_vfdiv ? _GEN_11946 : _GEN_10264; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12715 = io_op_bits_active_vfdiv ? _GEN_11947 : _GEN_10265; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12716 = io_op_bits_active_vfdiv ? _GEN_11948 : _GEN_10266; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12717 = io_op_bits_active_vfdiv ? _GEN_11949 : _GEN_10267; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12718 = io_op_bits_active_vfdiv ? _GEN_11950 : _GEN_10268; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12719 = io_op_bits_active_vfdiv ? _GEN_11951 : _GEN_10269; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12720 = io_op_bits_active_vfdiv ? _GEN_11952 : _GEN_10270; // @[sequencer-master.scala 645:40]
  wire [1:0] _GEN_12721 = io_op_bits_active_vfdiv ? _GEN_11953 : _GEN_10271; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12722 = io_op_bits_active_vfdiv ? _GEN_11954 : _GEN_10272; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12723 = io_op_bits_active_vfdiv ? _GEN_11955 : _GEN_10273; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12724 = io_op_bits_active_vfdiv ? _GEN_11956 : _GEN_10274; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12725 = io_op_bits_active_vfdiv ? _GEN_11957 : _GEN_10275; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12726 = io_op_bits_active_vfdiv ? _GEN_11958 : _GEN_10276; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12727 = io_op_bits_active_vfdiv ? _GEN_11959 : _GEN_10277; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12728 = io_op_bits_active_vfdiv ? _GEN_11960 : _GEN_10278; // @[sequencer-master.scala 645:40]
  wire [7:0] _GEN_12729 = io_op_bits_active_vfdiv ? _GEN_11961 : _GEN_10279; // @[sequencer-master.scala 645:40]
  wire  _GEN_12730 = io_op_bits_active_vfdiv | _GEN_10304; // @[sequencer-master.scala 645:40 sequencer-master.scala 265:41]
  wire [2:0] _GEN_12731 = io_op_bits_active_vfdiv ? _T_1647 : _GEN_10305; // @[sequencer-master.scala 645:40 sequencer-master.scala 265:66]
  wire  _GEN_12732 = _GEN_32729 | _GEN_12242; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12733 = _GEN_32730 | _GEN_12243; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12734 = _GEN_32731 | _GEN_12244; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12735 = _GEN_32732 | _GEN_12245; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12736 = _GEN_32733 | _GEN_12246; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12737 = _GEN_32734 | _GEN_12247; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12738 = _GEN_32735 | _GEN_12248; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12739 = _GEN_32736 | _GEN_12249; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_12748 = 3'h0 == tail ? 1'h0 : _GEN_12258; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12749 = 3'h1 == tail ? 1'h0 : _GEN_12259; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12750 = 3'h2 == tail ? 1'h0 : _GEN_12260; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12751 = 3'h3 == tail ? 1'h0 : _GEN_12261; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12752 = 3'h4 == tail ? 1'h0 : _GEN_12262; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12753 = 3'h5 == tail ? 1'h0 : _GEN_12263; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12754 = 3'h6 == tail ? 1'h0 : _GEN_12264; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12755 = 3'h7 == tail ? 1'h0 : _GEN_12265; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_12756 = 3'h0 == tail ? 1'h0 : _GEN_12266; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12757 = 3'h1 == tail ? 1'h0 : _GEN_12267; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12758 = 3'h2 == tail ? 1'h0 : _GEN_12268; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12759 = 3'h3 == tail ? 1'h0 : _GEN_12269; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12760 = 3'h4 == tail ? 1'h0 : _GEN_12270; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12761 = 3'h5 == tail ? 1'h0 : _GEN_12271; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12762 = 3'h6 == tail ? 1'h0 : _GEN_12272; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12763 = 3'h7 == tail ? 1'h0 : _GEN_12273; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_12764 = 3'h0 == tail ? 1'h0 : _GEN_12274; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12765 = 3'h1 == tail ? 1'h0 : _GEN_12275; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12766 = 3'h2 == tail ? 1'h0 : _GEN_12276; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12767 = 3'h3 == tail ? 1'h0 : _GEN_12277; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12768 = 3'h4 == tail ? 1'h0 : _GEN_12278; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12769 = 3'h5 == tail ? 1'h0 : _GEN_12279; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12770 = 3'h6 == tail ? 1'h0 : _GEN_12280; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12771 = 3'h7 == tail ? 1'h0 : _GEN_12281; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_12772 = 3'h0 == tail ? 1'h0 : _GEN_12282; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12773 = 3'h1 == tail ? 1'h0 : _GEN_12283; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12774 = 3'h2 == tail ? 1'h0 : _GEN_12284; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12775 = 3'h3 == tail ? 1'h0 : _GEN_12285; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12776 = 3'h4 == tail ? 1'h0 : _GEN_12286; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12777 = 3'h5 == tail ? 1'h0 : _GEN_12287; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12778 = 3'h6 == tail ? 1'h0 : _GEN_12288; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12779 = 3'h7 == tail ? 1'h0 : _GEN_12289; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_12780 = 3'h0 == tail ? 1'h0 : _GEN_12290; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12781 = 3'h1 == tail ? 1'h0 : _GEN_12291; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12782 = 3'h2 == tail ? 1'h0 : _GEN_12292; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12783 = 3'h3 == tail ? 1'h0 : _GEN_12293; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12784 = 3'h4 == tail ? 1'h0 : _GEN_12294; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12785 = 3'h5 == tail ? 1'h0 : _GEN_12295; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12786 = 3'h6 == tail ? 1'h0 : _GEN_12296; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12787 = 3'h7 == tail ? 1'h0 : _GEN_12297; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_12788 = _GEN_32729 | _GEN_12298; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12789 = _GEN_32730 | _GEN_12299; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12790 = _GEN_32731 | _GEN_12300; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12791 = _GEN_32732 | _GEN_12301; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12792 = _GEN_32733 | _GEN_12302; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12793 = _GEN_32734 | _GEN_12303; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12794 = _GEN_32735 | _GEN_12304; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12795 = _GEN_32736 | _GEN_12305; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_12796 = 3'h0 == tail ? 1'h0 : _GEN_12306; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12797 = 3'h1 == tail ? 1'h0 : _GEN_12307; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12798 = 3'h2 == tail ? 1'h0 : _GEN_12308; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12799 = 3'h3 == tail ? 1'h0 : _GEN_12309; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12800 = 3'h4 == tail ? 1'h0 : _GEN_12310; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12801 = 3'h5 == tail ? 1'h0 : _GEN_12311; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12802 = 3'h6 == tail ? 1'h0 : _GEN_12312; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12803 = 3'h7 == tail ? 1'h0 : _GEN_12313; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12804 = 3'h0 == tail ? 1'h0 : _GEN_12314; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12805 = 3'h1 == tail ? 1'h0 : _GEN_12315; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12806 = 3'h2 == tail ? 1'h0 : _GEN_12316; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12807 = 3'h3 == tail ? 1'h0 : _GEN_12317; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12808 = 3'h4 == tail ? 1'h0 : _GEN_12318; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12809 = 3'h5 == tail ? 1'h0 : _GEN_12319; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12810 = 3'h6 == tail ? 1'h0 : _GEN_12320; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12811 = 3'h7 == tail ? 1'h0 : _GEN_12321; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12812 = 3'h0 == tail ? 1'h0 : _GEN_12322; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12813 = 3'h1 == tail ? 1'h0 : _GEN_12323; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12814 = 3'h2 == tail ? 1'h0 : _GEN_12324; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12815 = 3'h3 == tail ? 1'h0 : _GEN_12325; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12816 = 3'h4 == tail ? 1'h0 : _GEN_12326; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12817 = 3'h5 == tail ? 1'h0 : _GEN_12327; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12818 = 3'h6 == tail ? 1'h0 : _GEN_12328; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12819 = 3'h7 == tail ? 1'h0 : _GEN_12329; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12820 = 3'h0 == tail ? 1'h0 : _GEN_12330; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12821 = 3'h1 == tail ? 1'h0 : _GEN_12331; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12822 = 3'h2 == tail ? 1'h0 : _GEN_12332; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12823 = 3'h3 == tail ? 1'h0 : _GEN_12333; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12824 = 3'h4 == tail ? 1'h0 : _GEN_12334; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12825 = 3'h5 == tail ? 1'h0 : _GEN_12335; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12826 = 3'h6 == tail ? 1'h0 : _GEN_12336; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12827 = 3'h7 == tail ? 1'h0 : _GEN_12337; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12828 = 3'h0 == tail ? 1'h0 : _GEN_12338; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12829 = 3'h1 == tail ? 1'h0 : _GEN_12339; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12830 = 3'h2 == tail ? 1'h0 : _GEN_12340; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12831 = 3'h3 == tail ? 1'h0 : _GEN_12341; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12832 = 3'h4 == tail ? 1'h0 : _GEN_12342; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12833 = 3'h5 == tail ? 1'h0 : _GEN_12343; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12834 = 3'h6 == tail ? 1'h0 : _GEN_12344; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12835 = 3'h7 == tail ? 1'h0 : _GEN_12345; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12836 = 3'h0 == tail ? 1'h0 : _GEN_12346; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12837 = 3'h1 == tail ? 1'h0 : _GEN_12347; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12838 = 3'h2 == tail ? 1'h0 : _GEN_12348; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12839 = 3'h3 == tail ? 1'h0 : _GEN_12349; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12840 = 3'h4 == tail ? 1'h0 : _GEN_12350; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12841 = 3'h5 == tail ? 1'h0 : _GEN_12351; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12842 = 3'h6 == tail ? 1'h0 : _GEN_12352; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12843 = 3'h7 == tail ? 1'h0 : _GEN_12353; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12844 = 3'h0 == tail ? 1'h0 : _GEN_12354; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12845 = 3'h1 == tail ? 1'h0 : _GEN_12355; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12846 = 3'h2 == tail ? 1'h0 : _GEN_12356; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12847 = 3'h3 == tail ? 1'h0 : _GEN_12357; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12848 = 3'h4 == tail ? 1'h0 : _GEN_12358; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12849 = 3'h5 == tail ? 1'h0 : _GEN_12359; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12850 = 3'h6 == tail ? 1'h0 : _GEN_12360; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12851 = 3'h7 == tail ? 1'h0 : _GEN_12361; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12852 = 3'h0 == tail ? 1'h0 : _GEN_12362; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12853 = 3'h1 == tail ? 1'h0 : _GEN_12363; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12854 = 3'h2 == tail ? 1'h0 : _GEN_12364; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12855 = 3'h3 == tail ? 1'h0 : _GEN_12365; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12856 = 3'h4 == tail ? 1'h0 : _GEN_12366; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12857 = 3'h5 == tail ? 1'h0 : _GEN_12367; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12858 = 3'h6 == tail ? 1'h0 : _GEN_12368; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12859 = 3'h7 == tail ? 1'h0 : _GEN_12369; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12860 = 3'h0 == tail ? 1'h0 : _GEN_12370; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12861 = 3'h1 == tail ? 1'h0 : _GEN_12371; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12862 = 3'h2 == tail ? 1'h0 : _GEN_12372; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12863 = 3'h3 == tail ? 1'h0 : _GEN_12373; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12864 = 3'h4 == tail ? 1'h0 : _GEN_12374; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12865 = 3'h5 == tail ? 1'h0 : _GEN_12375; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12866 = 3'h6 == tail ? 1'h0 : _GEN_12376; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12867 = 3'h7 == tail ? 1'h0 : _GEN_12377; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12868 = 3'h0 == tail ? 1'h0 : _GEN_12378; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12869 = 3'h1 == tail ? 1'h0 : _GEN_12379; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12870 = 3'h2 == tail ? 1'h0 : _GEN_12380; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12871 = 3'h3 == tail ? 1'h0 : _GEN_12381; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12872 = 3'h4 == tail ? 1'h0 : _GEN_12382; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12873 = 3'h5 == tail ? 1'h0 : _GEN_12383; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12874 = 3'h6 == tail ? 1'h0 : _GEN_12384; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12875 = 3'h7 == tail ? 1'h0 : _GEN_12385; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12876 = 3'h0 == tail ? 1'h0 : _GEN_12386; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12877 = 3'h1 == tail ? 1'h0 : _GEN_12387; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12878 = 3'h2 == tail ? 1'h0 : _GEN_12388; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12879 = 3'h3 == tail ? 1'h0 : _GEN_12389; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12880 = 3'h4 == tail ? 1'h0 : _GEN_12390; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12881 = 3'h5 == tail ? 1'h0 : _GEN_12391; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12882 = 3'h6 == tail ? 1'h0 : _GEN_12392; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12883 = 3'h7 == tail ? 1'h0 : _GEN_12393; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12884 = 3'h0 == tail ? 1'h0 : _GEN_12394; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12885 = 3'h1 == tail ? 1'h0 : _GEN_12395; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12886 = 3'h2 == tail ? 1'h0 : _GEN_12396; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12887 = 3'h3 == tail ? 1'h0 : _GEN_12397; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12888 = 3'h4 == tail ? 1'h0 : _GEN_12398; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12889 = 3'h5 == tail ? 1'h0 : _GEN_12399; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12890 = 3'h6 == tail ? 1'h0 : _GEN_12400; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12891 = 3'h7 == tail ? 1'h0 : _GEN_12401; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12892 = 3'h0 == tail ? 1'h0 : _GEN_12402; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12893 = 3'h1 == tail ? 1'h0 : _GEN_12403; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12894 = 3'h2 == tail ? 1'h0 : _GEN_12404; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12895 = 3'h3 == tail ? 1'h0 : _GEN_12405; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12896 = 3'h4 == tail ? 1'h0 : _GEN_12406; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12897 = 3'h5 == tail ? 1'h0 : _GEN_12407; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12898 = 3'h6 == tail ? 1'h0 : _GEN_12408; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12899 = 3'h7 == tail ? 1'h0 : _GEN_12409; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12900 = 3'h0 == tail ? 1'h0 : _GEN_12410; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12901 = 3'h1 == tail ? 1'h0 : _GEN_12411; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12902 = 3'h2 == tail ? 1'h0 : _GEN_12412; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12903 = 3'h3 == tail ? 1'h0 : _GEN_12413; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12904 = 3'h4 == tail ? 1'h0 : _GEN_12414; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12905 = 3'h5 == tail ? 1'h0 : _GEN_12415; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12906 = 3'h6 == tail ? 1'h0 : _GEN_12416; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12907 = 3'h7 == tail ? 1'h0 : _GEN_12417; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12908 = 3'h0 == tail ? 1'h0 : _GEN_12418; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12909 = 3'h1 == tail ? 1'h0 : _GEN_12419; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12910 = 3'h2 == tail ? 1'h0 : _GEN_12420; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12911 = 3'h3 == tail ? 1'h0 : _GEN_12421; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12912 = 3'h4 == tail ? 1'h0 : _GEN_12422; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12913 = 3'h5 == tail ? 1'h0 : _GEN_12423; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12914 = 3'h6 == tail ? 1'h0 : _GEN_12424; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12915 = 3'h7 == tail ? 1'h0 : _GEN_12425; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12916 = 3'h0 == tail ? 1'h0 : _GEN_12426; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12917 = 3'h1 == tail ? 1'h0 : _GEN_12427; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12918 = 3'h2 == tail ? 1'h0 : _GEN_12428; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12919 = 3'h3 == tail ? 1'h0 : _GEN_12429; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12920 = 3'h4 == tail ? 1'h0 : _GEN_12430; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12921 = 3'h5 == tail ? 1'h0 : _GEN_12431; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12922 = 3'h6 == tail ? 1'h0 : _GEN_12432; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12923 = 3'h7 == tail ? 1'h0 : _GEN_12433; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12924 = 3'h0 == tail ? 1'h0 : _GEN_12434; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12925 = 3'h1 == tail ? 1'h0 : _GEN_12435; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12926 = 3'h2 == tail ? 1'h0 : _GEN_12436; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12927 = 3'h3 == tail ? 1'h0 : _GEN_12437; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12928 = 3'h4 == tail ? 1'h0 : _GEN_12438; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12929 = 3'h5 == tail ? 1'h0 : _GEN_12439; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12930 = 3'h6 == tail ? 1'h0 : _GEN_12440; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12931 = 3'h7 == tail ? 1'h0 : _GEN_12441; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12932 = 3'h0 == tail ? 1'h0 : _GEN_12442; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12933 = 3'h1 == tail ? 1'h0 : _GEN_12443; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12934 = 3'h2 == tail ? 1'h0 : _GEN_12444; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12935 = 3'h3 == tail ? 1'h0 : _GEN_12445; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12936 = 3'h4 == tail ? 1'h0 : _GEN_12446; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12937 = 3'h5 == tail ? 1'h0 : _GEN_12447; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12938 = 3'h6 == tail ? 1'h0 : _GEN_12448; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12939 = 3'h7 == tail ? 1'h0 : _GEN_12449; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12940 = 3'h0 == tail ? 1'h0 : _GEN_12450; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12941 = 3'h1 == tail ? 1'h0 : _GEN_12451; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12942 = 3'h2 == tail ? 1'h0 : _GEN_12452; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12943 = 3'h3 == tail ? 1'h0 : _GEN_12453; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12944 = 3'h4 == tail ? 1'h0 : _GEN_12454; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12945 = 3'h5 == tail ? 1'h0 : _GEN_12455; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12946 = 3'h6 == tail ? 1'h0 : _GEN_12456; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12947 = 3'h7 == tail ? 1'h0 : _GEN_12457; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12948 = 3'h0 == tail ? 1'h0 : _GEN_12458; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12949 = 3'h1 == tail ? 1'h0 : _GEN_12459; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12950 = 3'h2 == tail ? 1'h0 : _GEN_12460; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12951 = 3'h3 == tail ? 1'h0 : _GEN_12461; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12952 = 3'h4 == tail ? 1'h0 : _GEN_12462; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12953 = 3'h5 == tail ? 1'h0 : _GEN_12463; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12954 = 3'h6 == tail ? 1'h0 : _GEN_12464; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12955 = 3'h7 == tail ? 1'h0 : _GEN_12465; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12956 = 3'h0 == tail ? 1'h0 : _GEN_12466; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12957 = 3'h1 == tail ? 1'h0 : _GEN_12467; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12958 = 3'h2 == tail ? 1'h0 : _GEN_12468; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12959 = 3'h3 == tail ? 1'h0 : _GEN_12469; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12960 = 3'h4 == tail ? 1'h0 : _GEN_12470; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12961 = 3'h5 == tail ? 1'h0 : _GEN_12471; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12962 = 3'h6 == tail ? 1'h0 : _GEN_12472; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12963 = 3'h7 == tail ? 1'h0 : _GEN_12473; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12964 = 3'h0 == tail ? 1'h0 : _GEN_12474; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12965 = 3'h1 == tail ? 1'h0 : _GEN_12475; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12966 = 3'h2 == tail ? 1'h0 : _GEN_12476; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12967 = 3'h3 == tail ? 1'h0 : _GEN_12477; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12968 = 3'h4 == tail ? 1'h0 : _GEN_12478; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12969 = 3'h5 == tail ? 1'h0 : _GEN_12479; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12970 = 3'h6 == tail ? 1'h0 : _GEN_12480; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12971 = 3'h7 == tail ? 1'h0 : _GEN_12481; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_12972 = 3'h0 == tail ? 1'h0 : _GEN_12482; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12973 = 3'h1 == tail ? 1'h0 : _GEN_12483; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12974 = 3'h2 == tail ? 1'h0 : _GEN_12484; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12975 = 3'h3 == tail ? 1'h0 : _GEN_12485; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12976 = 3'h4 == tail ? 1'h0 : _GEN_12486; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12977 = 3'h5 == tail ? 1'h0 : _GEN_12487; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12978 = 3'h6 == tail ? 1'h0 : _GEN_12488; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12979 = 3'h7 == tail ? 1'h0 : _GEN_12489; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_12980 = 3'h0 == tail ? 1'h0 : _GEN_12490; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12981 = 3'h1 == tail ? 1'h0 : _GEN_12491; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12982 = 3'h2 == tail ? 1'h0 : _GEN_12492; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12983 = 3'h3 == tail ? 1'h0 : _GEN_12493; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12984 = 3'h4 == tail ? 1'h0 : _GEN_12494; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12985 = 3'h5 == tail ? 1'h0 : _GEN_12495; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12986 = 3'h6 == tail ? 1'h0 : _GEN_12496; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12987 = 3'h7 == tail ? 1'h0 : _GEN_12497; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_12988 = 3'h0 == tail ? 1'h0 : _GEN_12498; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12989 = 3'h1 == tail ? 1'h0 : _GEN_12499; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12990 = 3'h2 == tail ? 1'h0 : _GEN_12500; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12991 = 3'h3 == tail ? 1'h0 : _GEN_12501; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12992 = 3'h4 == tail ? 1'h0 : _GEN_12502; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12993 = 3'h5 == tail ? 1'h0 : _GEN_12503; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12994 = 3'h6 == tail ? 1'h0 : _GEN_12504; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_12995 = 3'h7 == tail ? 1'h0 : _GEN_12505; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_13004 = _GEN_32729 | e_0_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13005 = _GEN_32730 | e_1_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13006 = _GEN_32731 | e_2_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13007 = _GEN_32732 | e_3_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13008 = _GEN_32733 | e_4_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13009 = _GEN_32734 | e_5_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13010 = _GEN_32735 | e_6_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_13011 = _GEN_32736 | e_7_active_vfcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_13012 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_12522; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13013 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_12523; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13014 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_12524; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13015 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_12525; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13016 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_12526; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13017 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_12527; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13018 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_12528; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_13019 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_12529; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_13020 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_12530; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13021 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_12531; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13022 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_12532; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13023 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_12533; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13024 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_12534; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13025 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_12535; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13026 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_12536; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_13027 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_12537; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13028 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_12748; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13029 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_12749; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13030 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_12750; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13031 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_12751; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13032 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_12752; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13033 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_12753; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13034 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_12754; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13035 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_12755; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13036 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_12538; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13037 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_12539; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13038 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_12540; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13039 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_12541; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13040 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_12542; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13041 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_12543; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13042 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_12544; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13043 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_12545; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13044 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_12546; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13045 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_12547; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13046 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_12548; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13047 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_12549; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13048 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_12550; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13049 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_12551; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13050 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_12552; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_13051 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_12553; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_13052 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_12554; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13053 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_12555; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13054 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_12556; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13055 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_12557; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13056 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_12558; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13057 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_12559; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13058 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_12560; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_13059 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_12561; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_13060 = io_op_bits_base_vp_valid ? _GEN_13020 : _GEN_12530; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13061 = io_op_bits_base_vp_valid ? _GEN_13021 : _GEN_12531; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13062 = io_op_bits_base_vp_valid ? _GEN_13022 : _GEN_12532; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13063 = io_op_bits_base_vp_valid ? _GEN_13023 : _GEN_12533; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13064 = io_op_bits_base_vp_valid ? _GEN_13024 : _GEN_12534; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13065 = io_op_bits_base_vp_valid ? _GEN_13025 : _GEN_12535; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13066 = io_op_bits_base_vp_valid ? _GEN_13026 : _GEN_12536; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_13067 = io_op_bits_base_vp_valid ? _GEN_13027 : _GEN_12537; // @[sequencer-master.scala 320:41]
  wire  _GEN_13068 = io_op_bits_base_vp_valid ? _GEN_13028 : _GEN_12748; // @[sequencer-master.scala 320:41]
  wire  _GEN_13069 = io_op_bits_base_vp_valid ? _GEN_13029 : _GEN_12749; // @[sequencer-master.scala 320:41]
  wire  _GEN_13070 = io_op_bits_base_vp_valid ? _GEN_13030 : _GEN_12750; // @[sequencer-master.scala 320:41]
  wire  _GEN_13071 = io_op_bits_base_vp_valid ? _GEN_13031 : _GEN_12751; // @[sequencer-master.scala 320:41]
  wire  _GEN_13072 = io_op_bits_base_vp_valid ? _GEN_13032 : _GEN_12752; // @[sequencer-master.scala 320:41]
  wire  _GEN_13073 = io_op_bits_base_vp_valid ? _GEN_13033 : _GEN_12753; // @[sequencer-master.scala 320:41]
  wire  _GEN_13074 = io_op_bits_base_vp_valid ? _GEN_13034 : _GEN_12754; // @[sequencer-master.scala 320:41]
  wire  _GEN_13075 = io_op_bits_base_vp_valid ? _GEN_13035 : _GEN_12755; // @[sequencer-master.scala 320:41]
  wire  _GEN_13076 = io_op_bits_base_vp_valid ? _GEN_13036 : _GEN_12538; // @[sequencer-master.scala 320:41]
  wire  _GEN_13077 = io_op_bits_base_vp_valid ? _GEN_13037 : _GEN_12539; // @[sequencer-master.scala 320:41]
  wire  _GEN_13078 = io_op_bits_base_vp_valid ? _GEN_13038 : _GEN_12540; // @[sequencer-master.scala 320:41]
  wire  _GEN_13079 = io_op_bits_base_vp_valid ? _GEN_13039 : _GEN_12541; // @[sequencer-master.scala 320:41]
  wire  _GEN_13080 = io_op_bits_base_vp_valid ? _GEN_13040 : _GEN_12542; // @[sequencer-master.scala 320:41]
  wire  _GEN_13081 = io_op_bits_base_vp_valid ? _GEN_13041 : _GEN_12543; // @[sequencer-master.scala 320:41]
  wire  _GEN_13082 = io_op_bits_base_vp_valid ? _GEN_13042 : _GEN_12544; // @[sequencer-master.scala 320:41]
  wire  _GEN_13083 = io_op_bits_base_vp_valid ? _GEN_13043 : _GEN_12545; // @[sequencer-master.scala 320:41]
  wire  _GEN_13084 = io_op_bits_base_vp_valid ? _GEN_13044 : _GEN_12546; // @[sequencer-master.scala 320:41]
  wire  _GEN_13085 = io_op_bits_base_vp_valid ? _GEN_13045 : _GEN_12547; // @[sequencer-master.scala 320:41]
  wire  _GEN_13086 = io_op_bits_base_vp_valid ? _GEN_13046 : _GEN_12548; // @[sequencer-master.scala 320:41]
  wire  _GEN_13087 = io_op_bits_base_vp_valid ? _GEN_13047 : _GEN_12549; // @[sequencer-master.scala 320:41]
  wire  _GEN_13088 = io_op_bits_base_vp_valid ? _GEN_13048 : _GEN_12550; // @[sequencer-master.scala 320:41]
  wire  _GEN_13089 = io_op_bits_base_vp_valid ? _GEN_13049 : _GEN_12551; // @[sequencer-master.scala 320:41]
  wire  _GEN_13090 = io_op_bits_base_vp_valid ? _GEN_13050 : _GEN_12552; // @[sequencer-master.scala 320:41]
  wire  _GEN_13091 = io_op_bits_base_vp_valid ? _GEN_13051 : _GEN_12553; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13092 = io_op_bits_base_vp_valid ? _GEN_13052 : _GEN_12554; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13093 = io_op_bits_base_vp_valid ? _GEN_13053 : _GEN_12555; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13094 = io_op_bits_base_vp_valid ? _GEN_13054 : _GEN_12556; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13095 = io_op_bits_base_vp_valid ? _GEN_13055 : _GEN_12557; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13096 = io_op_bits_base_vp_valid ? _GEN_13056 : _GEN_12558; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13097 = io_op_bits_base_vp_valid ? _GEN_13057 : _GEN_12559; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13098 = io_op_bits_base_vp_valid ? _GEN_13058 : _GEN_12560; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_13099 = io_op_bits_base_vp_valid ? _GEN_13059 : _GEN_12561; // @[sequencer-master.scala 320:41]
  wire  _GEN_13100 = _GEN_32729 | _GEN_12796; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13101 = _GEN_32730 | _GEN_12797; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13102 = _GEN_32731 | _GEN_12798; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13103 = _GEN_32732 | _GEN_12799; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13104 = _GEN_32733 | _GEN_12800; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13105 = _GEN_32734 | _GEN_12801; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13106 = _GEN_32735 | _GEN_12802; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13107 = _GEN_32736 | _GEN_12803; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13108 = _T_26 ? _GEN_13100 : _GEN_12796; // @[sequencer-master.scala 154:24]
  wire  _GEN_13109 = _T_26 ? _GEN_13101 : _GEN_12797; // @[sequencer-master.scala 154:24]
  wire  _GEN_13110 = _T_26 ? _GEN_13102 : _GEN_12798; // @[sequencer-master.scala 154:24]
  wire  _GEN_13111 = _T_26 ? _GEN_13103 : _GEN_12799; // @[sequencer-master.scala 154:24]
  wire  _GEN_13112 = _T_26 ? _GEN_13104 : _GEN_12800; // @[sequencer-master.scala 154:24]
  wire  _GEN_13113 = _T_26 ? _GEN_13105 : _GEN_12801; // @[sequencer-master.scala 154:24]
  wire  _GEN_13114 = _T_26 ? _GEN_13106 : _GEN_12802; // @[sequencer-master.scala 154:24]
  wire  _GEN_13115 = _T_26 ? _GEN_13107 : _GEN_12803; // @[sequencer-master.scala 154:24]
  wire  _GEN_13116 = _GEN_32729 | _GEN_12820; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13117 = _GEN_32730 | _GEN_12821; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13118 = _GEN_32731 | _GEN_12822; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13119 = _GEN_32732 | _GEN_12823; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13120 = _GEN_32733 | _GEN_12824; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13121 = _GEN_32734 | _GEN_12825; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13122 = _GEN_32735 | _GEN_12826; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13123 = _GEN_32736 | _GEN_12827; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13124 = _T_48 ? _GEN_13116 : _GEN_12820; // @[sequencer-master.scala 154:24]
  wire  _GEN_13125 = _T_48 ? _GEN_13117 : _GEN_12821; // @[sequencer-master.scala 154:24]
  wire  _GEN_13126 = _T_48 ? _GEN_13118 : _GEN_12822; // @[sequencer-master.scala 154:24]
  wire  _GEN_13127 = _T_48 ? _GEN_13119 : _GEN_12823; // @[sequencer-master.scala 154:24]
  wire  _GEN_13128 = _T_48 ? _GEN_13120 : _GEN_12824; // @[sequencer-master.scala 154:24]
  wire  _GEN_13129 = _T_48 ? _GEN_13121 : _GEN_12825; // @[sequencer-master.scala 154:24]
  wire  _GEN_13130 = _T_48 ? _GEN_13122 : _GEN_12826; // @[sequencer-master.scala 154:24]
  wire  _GEN_13131 = _T_48 ? _GEN_13123 : _GEN_12827; // @[sequencer-master.scala 154:24]
  wire  _GEN_13132 = _GEN_32729 | _GEN_12844; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13133 = _GEN_32730 | _GEN_12845; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13134 = _GEN_32731 | _GEN_12846; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13135 = _GEN_32732 | _GEN_12847; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13136 = _GEN_32733 | _GEN_12848; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13137 = _GEN_32734 | _GEN_12849; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13138 = _GEN_32735 | _GEN_12850; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13139 = _GEN_32736 | _GEN_12851; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13140 = _T_70 ? _GEN_13132 : _GEN_12844; // @[sequencer-master.scala 154:24]
  wire  _GEN_13141 = _T_70 ? _GEN_13133 : _GEN_12845; // @[sequencer-master.scala 154:24]
  wire  _GEN_13142 = _T_70 ? _GEN_13134 : _GEN_12846; // @[sequencer-master.scala 154:24]
  wire  _GEN_13143 = _T_70 ? _GEN_13135 : _GEN_12847; // @[sequencer-master.scala 154:24]
  wire  _GEN_13144 = _T_70 ? _GEN_13136 : _GEN_12848; // @[sequencer-master.scala 154:24]
  wire  _GEN_13145 = _T_70 ? _GEN_13137 : _GEN_12849; // @[sequencer-master.scala 154:24]
  wire  _GEN_13146 = _T_70 ? _GEN_13138 : _GEN_12850; // @[sequencer-master.scala 154:24]
  wire  _GEN_13147 = _T_70 ? _GEN_13139 : _GEN_12851; // @[sequencer-master.scala 154:24]
  wire  _GEN_13148 = _GEN_32729 | _GEN_12868; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13149 = _GEN_32730 | _GEN_12869; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13150 = _GEN_32731 | _GEN_12870; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13151 = _GEN_32732 | _GEN_12871; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13152 = _GEN_32733 | _GEN_12872; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13153 = _GEN_32734 | _GEN_12873; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13154 = _GEN_32735 | _GEN_12874; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13155 = _GEN_32736 | _GEN_12875; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13156 = _T_92 ? _GEN_13148 : _GEN_12868; // @[sequencer-master.scala 154:24]
  wire  _GEN_13157 = _T_92 ? _GEN_13149 : _GEN_12869; // @[sequencer-master.scala 154:24]
  wire  _GEN_13158 = _T_92 ? _GEN_13150 : _GEN_12870; // @[sequencer-master.scala 154:24]
  wire  _GEN_13159 = _T_92 ? _GEN_13151 : _GEN_12871; // @[sequencer-master.scala 154:24]
  wire  _GEN_13160 = _T_92 ? _GEN_13152 : _GEN_12872; // @[sequencer-master.scala 154:24]
  wire  _GEN_13161 = _T_92 ? _GEN_13153 : _GEN_12873; // @[sequencer-master.scala 154:24]
  wire  _GEN_13162 = _T_92 ? _GEN_13154 : _GEN_12874; // @[sequencer-master.scala 154:24]
  wire  _GEN_13163 = _T_92 ? _GEN_13155 : _GEN_12875; // @[sequencer-master.scala 154:24]
  wire  _GEN_13164 = _GEN_32729 | _GEN_12892; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13165 = _GEN_32730 | _GEN_12893; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13166 = _GEN_32731 | _GEN_12894; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13167 = _GEN_32732 | _GEN_12895; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13168 = _GEN_32733 | _GEN_12896; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13169 = _GEN_32734 | _GEN_12897; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13170 = _GEN_32735 | _GEN_12898; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13171 = _GEN_32736 | _GEN_12899; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13172 = _T_114 ? _GEN_13164 : _GEN_12892; // @[sequencer-master.scala 154:24]
  wire  _GEN_13173 = _T_114 ? _GEN_13165 : _GEN_12893; // @[sequencer-master.scala 154:24]
  wire  _GEN_13174 = _T_114 ? _GEN_13166 : _GEN_12894; // @[sequencer-master.scala 154:24]
  wire  _GEN_13175 = _T_114 ? _GEN_13167 : _GEN_12895; // @[sequencer-master.scala 154:24]
  wire  _GEN_13176 = _T_114 ? _GEN_13168 : _GEN_12896; // @[sequencer-master.scala 154:24]
  wire  _GEN_13177 = _T_114 ? _GEN_13169 : _GEN_12897; // @[sequencer-master.scala 154:24]
  wire  _GEN_13178 = _T_114 ? _GEN_13170 : _GEN_12898; // @[sequencer-master.scala 154:24]
  wire  _GEN_13179 = _T_114 ? _GEN_13171 : _GEN_12899; // @[sequencer-master.scala 154:24]
  wire  _GEN_13180 = _GEN_32729 | _GEN_12916; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13181 = _GEN_32730 | _GEN_12917; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13182 = _GEN_32731 | _GEN_12918; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13183 = _GEN_32732 | _GEN_12919; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13184 = _GEN_32733 | _GEN_12920; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13185 = _GEN_32734 | _GEN_12921; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13186 = _GEN_32735 | _GEN_12922; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13187 = _GEN_32736 | _GEN_12923; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13188 = _T_136 ? _GEN_13180 : _GEN_12916; // @[sequencer-master.scala 154:24]
  wire  _GEN_13189 = _T_136 ? _GEN_13181 : _GEN_12917; // @[sequencer-master.scala 154:24]
  wire  _GEN_13190 = _T_136 ? _GEN_13182 : _GEN_12918; // @[sequencer-master.scala 154:24]
  wire  _GEN_13191 = _T_136 ? _GEN_13183 : _GEN_12919; // @[sequencer-master.scala 154:24]
  wire  _GEN_13192 = _T_136 ? _GEN_13184 : _GEN_12920; // @[sequencer-master.scala 154:24]
  wire  _GEN_13193 = _T_136 ? _GEN_13185 : _GEN_12921; // @[sequencer-master.scala 154:24]
  wire  _GEN_13194 = _T_136 ? _GEN_13186 : _GEN_12922; // @[sequencer-master.scala 154:24]
  wire  _GEN_13195 = _T_136 ? _GEN_13187 : _GEN_12923; // @[sequencer-master.scala 154:24]
  wire  _GEN_13196 = _GEN_32729 | _GEN_12940; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13197 = _GEN_32730 | _GEN_12941; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13198 = _GEN_32731 | _GEN_12942; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13199 = _GEN_32732 | _GEN_12943; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13200 = _GEN_32733 | _GEN_12944; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13201 = _GEN_32734 | _GEN_12945; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13202 = _GEN_32735 | _GEN_12946; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13203 = _GEN_32736 | _GEN_12947; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13204 = _T_158 ? _GEN_13196 : _GEN_12940; // @[sequencer-master.scala 154:24]
  wire  _GEN_13205 = _T_158 ? _GEN_13197 : _GEN_12941; // @[sequencer-master.scala 154:24]
  wire  _GEN_13206 = _T_158 ? _GEN_13198 : _GEN_12942; // @[sequencer-master.scala 154:24]
  wire  _GEN_13207 = _T_158 ? _GEN_13199 : _GEN_12943; // @[sequencer-master.scala 154:24]
  wire  _GEN_13208 = _T_158 ? _GEN_13200 : _GEN_12944; // @[sequencer-master.scala 154:24]
  wire  _GEN_13209 = _T_158 ? _GEN_13201 : _GEN_12945; // @[sequencer-master.scala 154:24]
  wire  _GEN_13210 = _T_158 ? _GEN_13202 : _GEN_12946; // @[sequencer-master.scala 154:24]
  wire  _GEN_13211 = _T_158 ? _GEN_13203 : _GEN_12947; // @[sequencer-master.scala 154:24]
  wire  _GEN_13212 = _GEN_32729 | _GEN_12964; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13213 = _GEN_32730 | _GEN_12965; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13214 = _GEN_32731 | _GEN_12966; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13215 = _GEN_32732 | _GEN_12967; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13216 = _GEN_32733 | _GEN_12968; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13217 = _GEN_32734 | _GEN_12969; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13218 = _GEN_32735 | _GEN_12970; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13219 = _GEN_32736 | _GEN_12971; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13220 = _T_180 ? _GEN_13212 : _GEN_12964; // @[sequencer-master.scala 154:24]
  wire  _GEN_13221 = _T_180 ? _GEN_13213 : _GEN_12965; // @[sequencer-master.scala 154:24]
  wire  _GEN_13222 = _T_180 ? _GEN_13214 : _GEN_12966; // @[sequencer-master.scala 154:24]
  wire  _GEN_13223 = _T_180 ? _GEN_13215 : _GEN_12967; // @[sequencer-master.scala 154:24]
  wire  _GEN_13224 = _T_180 ? _GEN_13216 : _GEN_12968; // @[sequencer-master.scala 154:24]
  wire  _GEN_13225 = _T_180 ? _GEN_13217 : _GEN_12969; // @[sequencer-master.scala 154:24]
  wire  _GEN_13226 = _T_180 ? _GEN_13218 : _GEN_12970; // @[sequencer-master.scala 154:24]
  wire  _GEN_13227 = _T_180 ? _GEN_13219 : _GEN_12971; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_13228 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_12562; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13229 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_12563; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13230 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_12564; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13231 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_12565; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13232 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_12566; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13233 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_12567; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13234 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_12568; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13235 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_12569; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13236 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_12756; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13237 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_12757; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13238 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_12758; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13239 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_12759; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13240 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_12760; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13241 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_12761; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13242 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_12762; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13243 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_12763; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13244 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_12570; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13245 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_12571; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13246 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_12572; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13247 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_12573; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13248 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_12574; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13249 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_12575; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13250 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_12576; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13251 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_12577; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13252 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_12578; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13253 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_12579; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13254 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_12580; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13255 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_12581; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13256 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_12582; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13257 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_12583; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13258 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_12584; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13259 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_12585; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13260 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_12586; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13261 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_12587; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13262 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_12588; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13263 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_12589; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13264 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_12590; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13265 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_12591; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13266 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_12592; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_13267 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_12593; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13268 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_12594; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13269 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_12595; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13270 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_12596; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13271 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_12597; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13272 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_12598; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13273 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_12599; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13274 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_12600; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13275 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_12601; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_13276 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_12602; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13277 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_12603; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13278 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_12604; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13279 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_12605; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13280 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_12606; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13281 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_12607; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13282 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_12608; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13283 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_12609; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13284 = _T_189 ? _GEN_13276 : _GEN_12602; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13285 = _T_189 ? _GEN_13277 : _GEN_12603; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13286 = _T_189 ? _GEN_13278 : _GEN_12604; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13287 = _T_189 ? _GEN_13279 : _GEN_12605; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13288 = _T_189 ? _GEN_13280 : _GEN_12606; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13289 = _T_189 ? _GEN_13281 : _GEN_12607; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13290 = _T_189 ? _GEN_13282 : _GEN_12608; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_13291 = _T_189 ? _GEN_13283 : _GEN_12609; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_13292 = io_op_bits_base_vs1_valid ? _GEN_13228 : _GEN_12562; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13293 = io_op_bits_base_vs1_valid ? _GEN_13229 : _GEN_12563; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13294 = io_op_bits_base_vs1_valid ? _GEN_13230 : _GEN_12564; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13295 = io_op_bits_base_vs1_valid ? _GEN_13231 : _GEN_12565; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13296 = io_op_bits_base_vs1_valid ? _GEN_13232 : _GEN_12566; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13297 = io_op_bits_base_vs1_valid ? _GEN_13233 : _GEN_12567; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13298 = io_op_bits_base_vs1_valid ? _GEN_13234 : _GEN_12568; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13299 = io_op_bits_base_vs1_valid ? _GEN_13235 : _GEN_12569; // @[sequencer-master.scala 328:47]
  wire  _GEN_13300 = io_op_bits_base_vs1_valid ? _GEN_13236 : _GEN_12756; // @[sequencer-master.scala 328:47]
  wire  _GEN_13301 = io_op_bits_base_vs1_valid ? _GEN_13237 : _GEN_12757; // @[sequencer-master.scala 328:47]
  wire  _GEN_13302 = io_op_bits_base_vs1_valid ? _GEN_13238 : _GEN_12758; // @[sequencer-master.scala 328:47]
  wire  _GEN_13303 = io_op_bits_base_vs1_valid ? _GEN_13239 : _GEN_12759; // @[sequencer-master.scala 328:47]
  wire  _GEN_13304 = io_op_bits_base_vs1_valid ? _GEN_13240 : _GEN_12760; // @[sequencer-master.scala 328:47]
  wire  _GEN_13305 = io_op_bits_base_vs1_valid ? _GEN_13241 : _GEN_12761; // @[sequencer-master.scala 328:47]
  wire  _GEN_13306 = io_op_bits_base_vs1_valid ? _GEN_13242 : _GEN_12762; // @[sequencer-master.scala 328:47]
  wire  _GEN_13307 = io_op_bits_base_vs1_valid ? _GEN_13243 : _GEN_12763; // @[sequencer-master.scala 328:47]
  wire  _GEN_13308 = io_op_bits_base_vs1_valid ? _GEN_13244 : _GEN_12570; // @[sequencer-master.scala 328:47]
  wire  _GEN_13309 = io_op_bits_base_vs1_valid ? _GEN_13245 : _GEN_12571; // @[sequencer-master.scala 328:47]
  wire  _GEN_13310 = io_op_bits_base_vs1_valid ? _GEN_13246 : _GEN_12572; // @[sequencer-master.scala 328:47]
  wire  _GEN_13311 = io_op_bits_base_vs1_valid ? _GEN_13247 : _GEN_12573; // @[sequencer-master.scala 328:47]
  wire  _GEN_13312 = io_op_bits_base_vs1_valid ? _GEN_13248 : _GEN_12574; // @[sequencer-master.scala 328:47]
  wire  _GEN_13313 = io_op_bits_base_vs1_valid ? _GEN_13249 : _GEN_12575; // @[sequencer-master.scala 328:47]
  wire  _GEN_13314 = io_op_bits_base_vs1_valid ? _GEN_13250 : _GEN_12576; // @[sequencer-master.scala 328:47]
  wire  _GEN_13315 = io_op_bits_base_vs1_valid ? _GEN_13251 : _GEN_12577; // @[sequencer-master.scala 328:47]
  wire  _GEN_13316 = io_op_bits_base_vs1_valid ? _GEN_13252 : _GEN_12578; // @[sequencer-master.scala 328:47]
  wire  _GEN_13317 = io_op_bits_base_vs1_valid ? _GEN_13253 : _GEN_12579; // @[sequencer-master.scala 328:47]
  wire  _GEN_13318 = io_op_bits_base_vs1_valid ? _GEN_13254 : _GEN_12580; // @[sequencer-master.scala 328:47]
  wire  _GEN_13319 = io_op_bits_base_vs1_valid ? _GEN_13255 : _GEN_12581; // @[sequencer-master.scala 328:47]
  wire  _GEN_13320 = io_op_bits_base_vs1_valid ? _GEN_13256 : _GEN_12582; // @[sequencer-master.scala 328:47]
  wire  _GEN_13321 = io_op_bits_base_vs1_valid ? _GEN_13257 : _GEN_12583; // @[sequencer-master.scala 328:47]
  wire  _GEN_13322 = io_op_bits_base_vs1_valid ? _GEN_13258 : _GEN_12584; // @[sequencer-master.scala 328:47]
  wire  _GEN_13323 = io_op_bits_base_vs1_valid ? _GEN_13259 : _GEN_12585; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13324 = io_op_bits_base_vs1_valid ? _GEN_13260 : _GEN_12586; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13325 = io_op_bits_base_vs1_valid ? _GEN_13261 : _GEN_12587; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13326 = io_op_bits_base_vs1_valid ? _GEN_13262 : _GEN_12588; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13327 = io_op_bits_base_vs1_valid ? _GEN_13263 : _GEN_12589; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13328 = io_op_bits_base_vs1_valid ? _GEN_13264 : _GEN_12590; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13329 = io_op_bits_base_vs1_valid ? _GEN_13265 : _GEN_12591; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13330 = io_op_bits_base_vs1_valid ? _GEN_13266 : _GEN_12592; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_13331 = io_op_bits_base_vs1_valid ? _GEN_13267 : _GEN_12593; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13332 = io_op_bits_base_vs1_valid ? _GEN_13268 : _GEN_12594; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13333 = io_op_bits_base_vs1_valid ? _GEN_13269 : _GEN_12595; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13334 = io_op_bits_base_vs1_valid ? _GEN_13270 : _GEN_12596; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13335 = io_op_bits_base_vs1_valid ? _GEN_13271 : _GEN_12597; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13336 = io_op_bits_base_vs1_valid ? _GEN_13272 : _GEN_12598; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13337 = io_op_bits_base_vs1_valid ? _GEN_13273 : _GEN_12599; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13338 = io_op_bits_base_vs1_valid ? _GEN_13274 : _GEN_12600; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13339 = io_op_bits_base_vs1_valid ? _GEN_13275 : _GEN_12601; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13340 = io_op_bits_base_vs1_valid ? _GEN_13284 : _GEN_12602; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13341 = io_op_bits_base_vs1_valid ? _GEN_13285 : _GEN_12603; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13342 = io_op_bits_base_vs1_valid ? _GEN_13286 : _GEN_12604; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13343 = io_op_bits_base_vs1_valid ? _GEN_13287 : _GEN_12605; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13344 = io_op_bits_base_vs1_valid ? _GEN_13288 : _GEN_12606; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13345 = io_op_bits_base_vs1_valid ? _GEN_13289 : _GEN_12607; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13346 = io_op_bits_base_vs1_valid ? _GEN_13290 : _GEN_12608; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_13347 = io_op_bits_base_vs1_valid ? _GEN_13291 : _GEN_12609; // @[sequencer-master.scala 328:47]
  wire  _GEN_13348 = _GEN_32729 | _GEN_13108; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13349 = _GEN_32730 | _GEN_13109; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13350 = _GEN_32731 | _GEN_13110; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13351 = _GEN_32732 | _GEN_13111; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13352 = _GEN_32733 | _GEN_13112; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13353 = _GEN_32734 | _GEN_13113; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13354 = _GEN_32735 | _GEN_13114; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13355 = _GEN_32736 | _GEN_13115; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13356 = _T_203 ? _GEN_13348 : _GEN_13108; // @[sequencer-master.scala 154:24]
  wire  _GEN_13357 = _T_203 ? _GEN_13349 : _GEN_13109; // @[sequencer-master.scala 154:24]
  wire  _GEN_13358 = _T_203 ? _GEN_13350 : _GEN_13110; // @[sequencer-master.scala 154:24]
  wire  _GEN_13359 = _T_203 ? _GEN_13351 : _GEN_13111; // @[sequencer-master.scala 154:24]
  wire  _GEN_13360 = _T_203 ? _GEN_13352 : _GEN_13112; // @[sequencer-master.scala 154:24]
  wire  _GEN_13361 = _T_203 ? _GEN_13353 : _GEN_13113; // @[sequencer-master.scala 154:24]
  wire  _GEN_13362 = _T_203 ? _GEN_13354 : _GEN_13114; // @[sequencer-master.scala 154:24]
  wire  _GEN_13363 = _T_203 ? _GEN_13355 : _GEN_13115; // @[sequencer-master.scala 154:24]
  wire  _GEN_13364 = _GEN_32729 | _GEN_13124; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13365 = _GEN_32730 | _GEN_13125; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13366 = _GEN_32731 | _GEN_13126; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13367 = _GEN_32732 | _GEN_13127; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13368 = _GEN_32733 | _GEN_13128; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13369 = _GEN_32734 | _GEN_13129; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13370 = _GEN_32735 | _GEN_13130; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13371 = _GEN_32736 | _GEN_13131; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13372 = _T_225 ? _GEN_13364 : _GEN_13124; // @[sequencer-master.scala 154:24]
  wire  _GEN_13373 = _T_225 ? _GEN_13365 : _GEN_13125; // @[sequencer-master.scala 154:24]
  wire  _GEN_13374 = _T_225 ? _GEN_13366 : _GEN_13126; // @[sequencer-master.scala 154:24]
  wire  _GEN_13375 = _T_225 ? _GEN_13367 : _GEN_13127; // @[sequencer-master.scala 154:24]
  wire  _GEN_13376 = _T_225 ? _GEN_13368 : _GEN_13128; // @[sequencer-master.scala 154:24]
  wire  _GEN_13377 = _T_225 ? _GEN_13369 : _GEN_13129; // @[sequencer-master.scala 154:24]
  wire  _GEN_13378 = _T_225 ? _GEN_13370 : _GEN_13130; // @[sequencer-master.scala 154:24]
  wire  _GEN_13379 = _T_225 ? _GEN_13371 : _GEN_13131; // @[sequencer-master.scala 154:24]
  wire  _GEN_13380 = _GEN_32729 | _GEN_13140; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13381 = _GEN_32730 | _GEN_13141; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13382 = _GEN_32731 | _GEN_13142; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13383 = _GEN_32732 | _GEN_13143; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13384 = _GEN_32733 | _GEN_13144; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13385 = _GEN_32734 | _GEN_13145; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13386 = _GEN_32735 | _GEN_13146; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13387 = _GEN_32736 | _GEN_13147; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13388 = _T_247 ? _GEN_13380 : _GEN_13140; // @[sequencer-master.scala 154:24]
  wire  _GEN_13389 = _T_247 ? _GEN_13381 : _GEN_13141; // @[sequencer-master.scala 154:24]
  wire  _GEN_13390 = _T_247 ? _GEN_13382 : _GEN_13142; // @[sequencer-master.scala 154:24]
  wire  _GEN_13391 = _T_247 ? _GEN_13383 : _GEN_13143; // @[sequencer-master.scala 154:24]
  wire  _GEN_13392 = _T_247 ? _GEN_13384 : _GEN_13144; // @[sequencer-master.scala 154:24]
  wire  _GEN_13393 = _T_247 ? _GEN_13385 : _GEN_13145; // @[sequencer-master.scala 154:24]
  wire  _GEN_13394 = _T_247 ? _GEN_13386 : _GEN_13146; // @[sequencer-master.scala 154:24]
  wire  _GEN_13395 = _T_247 ? _GEN_13387 : _GEN_13147; // @[sequencer-master.scala 154:24]
  wire  _GEN_13396 = _GEN_32729 | _GEN_13156; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13397 = _GEN_32730 | _GEN_13157; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13398 = _GEN_32731 | _GEN_13158; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13399 = _GEN_32732 | _GEN_13159; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13400 = _GEN_32733 | _GEN_13160; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13401 = _GEN_32734 | _GEN_13161; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13402 = _GEN_32735 | _GEN_13162; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13403 = _GEN_32736 | _GEN_13163; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13404 = _T_269 ? _GEN_13396 : _GEN_13156; // @[sequencer-master.scala 154:24]
  wire  _GEN_13405 = _T_269 ? _GEN_13397 : _GEN_13157; // @[sequencer-master.scala 154:24]
  wire  _GEN_13406 = _T_269 ? _GEN_13398 : _GEN_13158; // @[sequencer-master.scala 154:24]
  wire  _GEN_13407 = _T_269 ? _GEN_13399 : _GEN_13159; // @[sequencer-master.scala 154:24]
  wire  _GEN_13408 = _T_269 ? _GEN_13400 : _GEN_13160; // @[sequencer-master.scala 154:24]
  wire  _GEN_13409 = _T_269 ? _GEN_13401 : _GEN_13161; // @[sequencer-master.scala 154:24]
  wire  _GEN_13410 = _T_269 ? _GEN_13402 : _GEN_13162; // @[sequencer-master.scala 154:24]
  wire  _GEN_13411 = _T_269 ? _GEN_13403 : _GEN_13163; // @[sequencer-master.scala 154:24]
  wire  _GEN_13412 = _GEN_32729 | _GEN_13172; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13413 = _GEN_32730 | _GEN_13173; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13414 = _GEN_32731 | _GEN_13174; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13415 = _GEN_32732 | _GEN_13175; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13416 = _GEN_32733 | _GEN_13176; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13417 = _GEN_32734 | _GEN_13177; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13418 = _GEN_32735 | _GEN_13178; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13419 = _GEN_32736 | _GEN_13179; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13420 = _T_291 ? _GEN_13412 : _GEN_13172; // @[sequencer-master.scala 154:24]
  wire  _GEN_13421 = _T_291 ? _GEN_13413 : _GEN_13173; // @[sequencer-master.scala 154:24]
  wire  _GEN_13422 = _T_291 ? _GEN_13414 : _GEN_13174; // @[sequencer-master.scala 154:24]
  wire  _GEN_13423 = _T_291 ? _GEN_13415 : _GEN_13175; // @[sequencer-master.scala 154:24]
  wire  _GEN_13424 = _T_291 ? _GEN_13416 : _GEN_13176; // @[sequencer-master.scala 154:24]
  wire  _GEN_13425 = _T_291 ? _GEN_13417 : _GEN_13177; // @[sequencer-master.scala 154:24]
  wire  _GEN_13426 = _T_291 ? _GEN_13418 : _GEN_13178; // @[sequencer-master.scala 154:24]
  wire  _GEN_13427 = _T_291 ? _GEN_13419 : _GEN_13179; // @[sequencer-master.scala 154:24]
  wire  _GEN_13428 = _GEN_32729 | _GEN_13188; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13429 = _GEN_32730 | _GEN_13189; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13430 = _GEN_32731 | _GEN_13190; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13431 = _GEN_32732 | _GEN_13191; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13432 = _GEN_32733 | _GEN_13192; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13433 = _GEN_32734 | _GEN_13193; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13434 = _GEN_32735 | _GEN_13194; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13435 = _GEN_32736 | _GEN_13195; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13436 = _T_313 ? _GEN_13428 : _GEN_13188; // @[sequencer-master.scala 154:24]
  wire  _GEN_13437 = _T_313 ? _GEN_13429 : _GEN_13189; // @[sequencer-master.scala 154:24]
  wire  _GEN_13438 = _T_313 ? _GEN_13430 : _GEN_13190; // @[sequencer-master.scala 154:24]
  wire  _GEN_13439 = _T_313 ? _GEN_13431 : _GEN_13191; // @[sequencer-master.scala 154:24]
  wire  _GEN_13440 = _T_313 ? _GEN_13432 : _GEN_13192; // @[sequencer-master.scala 154:24]
  wire  _GEN_13441 = _T_313 ? _GEN_13433 : _GEN_13193; // @[sequencer-master.scala 154:24]
  wire  _GEN_13442 = _T_313 ? _GEN_13434 : _GEN_13194; // @[sequencer-master.scala 154:24]
  wire  _GEN_13443 = _T_313 ? _GEN_13435 : _GEN_13195; // @[sequencer-master.scala 154:24]
  wire  _GEN_13444 = _GEN_32729 | _GEN_13204; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13445 = _GEN_32730 | _GEN_13205; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13446 = _GEN_32731 | _GEN_13206; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13447 = _GEN_32732 | _GEN_13207; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13448 = _GEN_32733 | _GEN_13208; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13449 = _GEN_32734 | _GEN_13209; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13450 = _GEN_32735 | _GEN_13210; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13451 = _GEN_32736 | _GEN_13211; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13452 = _T_335 ? _GEN_13444 : _GEN_13204; // @[sequencer-master.scala 154:24]
  wire  _GEN_13453 = _T_335 ? _GEN_13445 : _GEN_13205; // @[sequencer-master.scala 154:24]
  wire  _GEN_13454 = _T_335 ? _GEN_13446 : _GEN_13206; // @[sequencer-master.scala 154:24]
  wire  _GEN_13455 = _T_335 ? _GEN_13447 : _GEN_13207; // @[sequencer-master.scala 154:24]
  wire  _GEN_13456 = _T_335 ? _GEN_13448 : _GEN_13208; // @[sequencer-master.scala 154:24]
  wire  _GEN_13457 = _T_335 ? _GEN_13449 : _GEN_13209; // @[sequencer-master.scala 154:24]
  wire  _GEN_13458 = _T_335 ? _GEN_13450 : _GEN_13210; // @[sequencer-master.scala 154:24]
  wire  _GEN_13459 = _T_335 ? _GEN_13451 : _GEN_13211; // @[sequencer-master.scala 154:24]
  wire  _GEN_13460 = _GEN_32729 | _GEN_13220; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13461 = _GEN_32730 | _GEN_13221; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13462 = _GEN_32731 | _GEN_13222; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13463 = _GEN_32732 | _GEN_13223; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13464 = _GEN_32733 | _GEN_13224; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13465 = _GEN_32734 | _GEN_13225; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13466 = _GEN_32735 | _GEN_13226; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13467 = _GEN_32736 | _GEN_13227; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13468 = _T_357 ? _GEN_13460 : _GEN_13220; // @[sequencer-master.scala 154:24]
  wire  _GEN_13469 = _T_357 ? _GEN_13461 : _GEN_13221; // @[sequencer-master.scala 154:24]
  wire  _GEN_13470 = _T_357 ? _GEN_13462 : _GEN_13222; // @[sequencer-master.scala 154:24]
  wire  _GEN_13471 = _T_357 ? _GEN_13463 : _GEN_13223; // @[sequencer-master.scala 154:24]
  wire  _GEN_13472 = _T_357 ? _GEN_13464 : _GEN_13224; // @[sequencer-master.scala 154:24]
  wire  _GEN_13473 = _T_357 ? _GEN_13465 : _GEN_13225; // @[sequencer-master.scala 154:24]
  wire  _GEN_13474 = _T_357 ? _GEN_13466 : _GEN_13226; // @[sequencer-master.scala 154:24]
  wire  _GEN_13475 = _T_357 ? _GEN_13467 : _GEN_13227; // @[sequencer-master.scala 154:24]
  wire  _GEN_13484 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_12764; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13485 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_12765; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13486 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_12766; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13487 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_12767; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13488 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_12768; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13489 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_12769; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13490 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_12770; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_13491 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_12771; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_13516 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_12642; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13517 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_12643; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13518 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_12644; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13519 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_12645; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13520 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_12646; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13521 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_12647; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13522 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_12648; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_13523 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_12649; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_13524 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_12650; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13525 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_12651; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13526 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_12652; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13527 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_12653; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13528 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_12654; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13529 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_12655; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13530 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_12656; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_13531 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_12657; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire  _GEN_13548 = io_op_bits_base_vs2_valid ? _GEN_13484 : _GEN_12764; // @[sequencer-master.scala 328:47]
  wire  _GEN_13549 = io_op_bits_base_vs2_valid ? _GEN_13485 : _GEN_12765; // @[sequencer-master.scala 328:47]
  wire  _GEN_13550 = io_op_bits_base_vs2_valid ? _GEN_13486 : _GEN_12766; // @[sequencer-master.scala 328:47]
  wire  _GEN_13551 = io_op_bits_base_vs2_valid ? _GEN_13487 : _GEN_12767; // @[sequencer-master.scala 328:47]
  wire  _GEN_13552 = io_op_bits_base_vs2_valid ? _GEN_13488 : _GEN_12768; // @[sequencer-master.scala 328:47]
  wire  _GEN_13553 = io_op_bits_base_vs2_valid ? _GEN_13489 : _GEN_12769; // @[sequencer-master.scala 328:47]
  wire  _GEN_13554 = io_op_bits_base_vs2_valid ? _GEN_13490 : _GEN_12770; // @[sequencer-master.scala 328:47]
  wire  _GEN_13555 = io_op_bits_base_vs2_valid ? _GEN_13491 : _GEN_12771; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13580 = io_op_bits_base_vs2_valid ? _GEN_13516 : _GEN_12642; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13581 = io_op_bits_base_vs2_valid ? _GEN_13517 : _GEN_12643; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13582 = io_op_bits_base_vs2_valid ? _GEN_13518 : _GEN_12644; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13583 = io_op_bits_base_vs2_valid ? _GEN_13519 : _GEN_12645; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13584 = io_op_bits_base_vs2_valid ? _GEN_13520 : _GEN_12646; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13585 = io_op_bits_base_vs2_valid ? _GEN_13521 : _GEN_12647; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13586 = io_op_bits_base_vs2_valid ? _GEN_13522 : _GEN_12648; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_13587 = io_op_bits_base_vs2_valid ? _GEN_13523 : _GEN_12649; // @[sequencer-master.scala 328:47]
  wire  _GEN_13596 = _GEN_32729 | _GEN_13356; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13597 = _GEN_32730 | _GEN_13357; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13598 = _GEN_32731 | _GEN_13358; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13599 = _GEN_32732 | _GEN_13359; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13600 = _GEN_32733 | _GEN_13360; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13601 = _GEN_32734 | _GEN_13361; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13602 = _GEN_32735 | _GEN_13362; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13603 = _GEN_32736 | _GEN_13363; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13604 = _T_380 ? _GEN_13596 : _GEN_13356; // @[sequencer-master.scala 154:24]
  wire  _GEN_13605 = _T_380 ? _GEN_13597 : _GEN_13357; // @[sequencer-master.scala 154:24]
  wire  _GEN_13606 = _T_380 ? _GEN_13598 : _GEN_13358; // @[sequencer-master.scala 154:24]
  wire  _GEN_13607 = _T_380 ? _GEN_13599 : _GEN_13359; // @[sequencer-master.scala 154:24]
  wire  _GEN_13608 = _T_380 ? _GEN_13600 : _GEN_13360; // @[sequencer-master.scala 154:24]
  wire  _GEN_13609 = _T_380 ? _GEN_13601 : _GEN_13361; // @[sequencer-master.scala 154:24]
  wire  _GEN_13610 = _T_380 ? _GEN_13602 : _GEN_13362; // @[sequencer-master.scala 154:24]
  wire  _GEN_13611 = _T_380 ? _GEN_13603 : _GEN_13363; // @[sequencer-master.scala 154:24]
  wire  _GEN_13612 = _GEN_32729 | _GEN_13372; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13613 = _GEN_32730 | _GEN_13373; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13614 = _GEN_32731 | _GEN_13374; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13615 = _GEN_32732 | _GEN_13375; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13616 = _GEN_32733 | _GEN_13376; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13617 = _GEN_32734 | _GEN_13377; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13618 = _GEN_32735 | _GEN_13378; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13619 = _GEN_32736 | _GEN_13379; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13620 = _T_402 ? _GEN_13612 : _GEN_13372; // @[sequencer-master.scala 154:24]
  wire  _GEN_13621 = _T_402 ? _GEN_13613 : _GEN_13373; // @[sequencer-master.scala 154:24]
  wire  _GEN_13622 = _T_402 ? _GEN_13614 : _GEN_13374; // @[sequencer-master.scala 154:24]
  wire  _GEN_13623 = _T_402 ? _GEN_13615 : _GEN_13375; // @[sequencer-master.scala 154:24]
  wire  _GEN_13624 = _T_402 ? _GEN_13616 : _GEN_13376; // @[sequencer-master.scala 154:24]
  wire  _GEN_13625 = _T_402 ? _GEN_13617 : _GEN_13377; // @[sequencer-master.scala 154:24]
  wire  _GEN_13626 = _T_402 ? _GEN_13618 : _GEN_13378; // @[sequencer-master.scala 154:24]
  wire  _GEN_13627 = _T_402 ? _GEN_13619 : _GEN_13379; // @[sequencer-master.scala 154:24]
  wire  _GEN_13628 = _GEN_32729 | _GEN_13388; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13629 = _GEN_32730 | _GEN_13389; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13630 = _GEN_32731 | _GEN_13390; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13631 = _GEN_32732 | _GEN_13391; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13632 = _GEN_32733 | _GEN_13392; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13633 = _GEN_32734 | _GEN_13393; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13634 = _GEN_32735 | _GEN_13394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13635 = _GEN_32736 | _GEN_13395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13636 = _T_424 ? _GEN_13628 : _GEN_13388; // @[sequencer-master.scala 154:24]
  wire  _GEN_13637 = _T_424 ? _GEN_13629 : _GEN_13389; // @[sequencer-master.scala 154:24]
  wire  _GEN_13638 = _T_424 ? _GEN_13630 : _GEN_13390; // @[sequencer-master.scala 154:24]
  wire  _GEN_13639 = _T_424 ? _GEN_13631 : _GEN_13391; // @[sequencer-master.scala 154:24]
  wire  _GEN_13640 = _T_424 ? _GEN_13632 : _GEN_13392; // @[sequencer-master.scala 154:24]
  wire  _GEN_13641 = _T_424 ? _GEN_13633 : _GEN_13393; // @[sequencer-master.scala 154:24]
  wire  _GEN_13642 = _T_424 ? _GEN_13634 : _GEN_13394; // @[sequencer-master.scala 154:24]
  wire  _GEN_13643 = _T_424 ? _GEN_13635 : _GEN_13395; // @[sequencer-master.scala 154:24]
  wire  _GEN_13644 = _GEN_32729 | _GEN_13404; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13645 = _GEN_32730 | _GEN_13405; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13646 = _GEN_32731 | _GEN_13406; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13647 = _GEN_32732 | _GEN_13407; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13648 = _GEN_32733 | _GEN_13408; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13649 = _GEN_32734 | _GEN_13409; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13650 = _GEN_32735 | _GEN_13410; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13651 = _GEN_32736 | _GEN_13411; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13652 = _T_446 ? _GEN_13644 : _GEN_13404; // @[sequencer-master.scala 154:24]
  wire  _GEN_13653 = _T_446 ? _GEN_13645 : _GEN_13405; // @[sequencer-master.scala 154:24]
  wire  _GEN_13654 = _T_446 ? _GEN_13646 : _GEN_13406; // @[sequencer-master.scala 154:24]
  wire  _GEN_13655 = _T_446 ? _GEN_13647 : _GEN_13407; // @[sequencer-master.scala 154:24]
  wire  _GEN_13656 = _T_446 ? _GEN_13648 : _GEN_13408; // @[sequencer-master.scala 154:24]
  wire  _GEN_13657 = _T_446 ? _GEN_13649 : _GEN_13409; // @[sequencer-master.scala 154:24]
  wire  _GEN_13658 = _T_446 ? _GEN_13650 : _GEN_13410; // @[sequencer-master.scala 154:24]
  wire  _GEN_13659 = _T_446 ? _GEN_13651 : _GEN_13411; // @[sequencer-master.scala 154:24]
  wire  _GEN_13660 = _GEN_32729 | _GEN_13420; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13661 = _GEN_32730 | _GEN_13421; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13662 = _GEN_32731 | _GEN_13422; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13663 = _GEN_32732 | _GEN_13423; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13664 = _GEN_32733 | _GEN_13424; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13665 = _GEN_32734 | _GEN_13425; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13666 = _GEN_32735 | _GEN_13426; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13667 = _GEN_32736 | _GEN_13427; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13668 = _T_468 ? _GEN_13660 : _GEN_13420; // @[sequencer-master.scala 154:24]
  wire  _GEN_13669 = _T_468 ? _GEN_13661 : _GEN_13421; // @[sequencer-master.scala 154:24]
  wire  _GEN_13670 = _T_468 ? _GEN_13662 : _GEN_13422; // @[sequencer-master.scala 154:24]
  wire  _GEN_13671 = _T_468 ? _GEN_13663 : _GEN_13423; // @[sequencer-master.scala 154:24]
  wire  _GEN_13672 = _T_468 ? _GEN_13664 : _GEN_13424; // @[sequencer-master.scala 154:24]
  wire  _GEN_13673 = _T_468 ? _GEN_13665 : _GEN_13425; // @[sequencer-master.scala 154:24]
  wire  _GEN_13674 = _T_468 ? _GEN_13666 : _GEN_13426; // @[sequencer-master.scala 154:24]
  wire  _GEN_13675 = _T_468 ? _GEN_13667 : _GEN_13427; // @[sequencer-master.scala 154:24]
  wire  _GEN_13676 = _GEN_32729 | _GEN_13436; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13677 = _GEN_32730 | _GEN_13437; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13678 = _GEN_32731 | _GEN_13438; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13679 = _GEN_32732 | _GEN_13439; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13680 = _GEN_32733 | _GEN_13440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13681 = _GEN_32734 | _GEN_13441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13682 = _GEN_32735 | _GEN_13442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13683 = _GEN_32736 | _GEN_13443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13684 = _T_490 ? _GEN_13676 : _GEN_13436; // @[sequencer-master.scala 154:24]
  wire  _GEN_13685 = _T_490 ? _GEN_13677 : _GEN_13437; // @[sequencer-master.scala 154:24]
  wire  _GEN_13686 = _T_490 ? _GEN_13678 : _GEN_13438; // @[sequencer-master.scala 154:24]
  wire  _GEN_13687 = _T_490 ? _GEN_13679 : _GEN_13439; // @[sequencer-master.scala 154:24]
  wire  _GEN_13688 = _T_490 ? _GEN_13680 : _GEN_13440; // @[sequencer-master.scala 154:24]
  wire  _GEN_13689 = _T_490 ? _GEN_13681 : _GEN_13441; // @[sequencer-master.scala 154:24]
  wire  _GEN_13690 = _T_490 ? _GEN_13682 : _GEN_13442; // @[sequencer-master.scala 154:24]
  wire  _GEN_13691 = _T_490 ? _GEN_13683 : _GEN_13443; // @[sequencer-master.scala 154:24]
  wire  _GEN_13692 = _GEN_32729 | _GEN_13452; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13693 = _GEN_32730 | _GEN_13453; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13694 = _GEN_32731 | _GEN_13454; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13695 = _GEN_32732 | _GEN_13455; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13696 = _GEN_32733 | _GEN_13456; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13697 = _GEN_32734 | _GEN_13457; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13698 = _GEN_32735 | _GEN_13458; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13699 = _GEN_32736 | _GEN_13459; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13700 = _T_512 ? _GEN_13692 : _GEN_13452; // @[sequencer-master.scala 154:24]
  wire  _GEN_13701 = _T_512 ? _GEN_13693 : _GEN_13453; // @[sequencer-master.scala 154:24]
  wire  _GEN_13702 = _T_512 ? _GEN_13694 : _GEN_13454; // @[sequencer-master.scala 154:24]
  wire  _GEN_13703 = _T_512 ? _GEN_13695 : _GEN_13455; // @[sequencer-master.scala 154:24]
  wire  _GEN_13704 = _T_512 ? _GEN_13696 : _GEN_13456; // @[sequencer-master.scala 154:24]
  wire  _GEN_13705 = _T_512 ? _GEN_13697 : _GEN_13457; // @[sequencer-master.scala 154:24]
  wire  _GEN_13706 = _T_512 ? _GEN_13698 : _GEN_13458; // @[sequencer-master.scala 154:24]
  wire  _GEN_13707 = _T_512 ? _GEN_13699 : _GEN_13459; // @[sequencer-master.scala 154:24]
  wire  _GEN_13708 = _GEN_32729 | _GEN_13468; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13709 = _GEN_32730 | _GEN_13469; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13710 = _GEN_32731 | _GEN_13470; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13711 = _GEN_32732 | _GEN_13471; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13712 = _GEN_32733 | _GEN_13472; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13713 = _GEN_32734 | _GEN_13473; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13714 = _GEN_32735 | _GEN_13474; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13715 = _GEN_32736 | _GEN_13475; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_13716 = _T_534 ? _GEN_13708 : _GEN_13468; // @[sequencer-master.scala 154:24]
  wire  _GEN_13717 = _T_534 ? _GEN_13709 : _GEN_13469; // @[sequencer-master.scala 154:24]
  wire  _GEN_13718 = _T_534 ? _GEN_13710 : _GEN_13470; // @[sequencer-master.scala 154:24]
  wire  _GEN_13719 = _T_534 ? _GEN_13711 : _GEN_13471; // @[sequencer-master.scala 154:24]
  wire  _GEN_13720 = _T_534 ? _GEN_13712 : _GEN_13472; // @[sequencer-master.scala 154:24]
  wire  _GEN_13721 = _T_534 ? _GEN_13713 : _GEN_13473; // @[sequencer-master.scala 154:24]
  wire  _GEN_13722 = _T_534 ? _GEN_13714 : _GEN_13474; // @[sequencer-master.scala 154:24]
  wire  _GEN_13723 = _T_534 ? _GEN_13715 : _GEN_13475; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_13724 = 3'h0 == tail ? io_op_bits_base_vd_id : _GEN_12690; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13725 = 3'h1 == tail ? io_op_bits_base_vd_id : _GEN_12691; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13726 = 3'h2 == tail ? io_op_bits_base_vd_id : _GEN_12692; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13727 = 3'h3 == tail ? io_op_bits_base_vd_id : _GEN_12693; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13728 = 3'h4 == tail ? io_op_bits_base_vd_id : _GEN_12694; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13729 = 3'h5 == tail ? io_op_bits_base_vd_id : _GEN_12695; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13730 = 3'h6 == tail ? io_op_bits_base_vd_id : _GEN_12696; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13731 = 3'h7 == tail ? io_op_bits_base_vd_id : _GEN_12697; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13732 = 3'h0 == tail ? io_op_bits_base_vd_valid : _GEN_12780; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13733 = 3'h1 == tail ? io_op_bits_base_vd_valid : _GEN_12781; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13734 = 3'h2 == tail ? io_op_bits_base_vd_valid : _GEN_12782; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13735 = 3'h3 == tail ? io_op_bits_base_vd_valid : _GEN_12783; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13736 = 3'h4 == tail ? io_op_bits_base_vd_valid : _GEN_12784; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13737 = 3'h5 == tail ? io_op_bits_base_vd_valid : _GEN_12785; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13738 = 3'h6 == tail ? io_op_bits_base_vd_valid : _GEN_12786; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13739 = 3'h7 == tail ? io_op_bits_base_vd_valid : _GEN_12787; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13740 = 3'h0 == tail ? io_op_bits_base_vd_scalar : _GEN_12698; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13741 = 3'h1 == tail ? io_op_bits_base_vd_scalar : _GEN_12699; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13742 = 3'h2 == tail ? io_op_bits_base_vd_scalar : _GEN_12700; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13743 = 3'h3 == tail ? io_op_bits_base_vd_scalar : _GEN_12701; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13744 = 3'h4 == tail ? io_op_bits_base_vd_scalar : _GEN_12702; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13745 = 3'h5 == tail ? io_op_bits_base_vd_scalar : _GEN_12703; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13746 = 3'h6 == tail ? io_op_bits_base_vd_scalar : _GEN_12704; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13747 = 3'h7 == tail ? io_op_bits_base_vd_scalar : _GEN_12705; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13748 = 3'h0 == tail ? io_op_bits_base_vd_pred : _GEN_12706; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13749 = 3'h1 == tail ? io_op_bits_base_vd_pred : _GEN_12707; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13750 = 3'h2 == tail ? io_op_bits_base_vd_pred : _GEN_12708; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13751 = 3'h3 == tail ? io_op_bits_base_vd_pred : _GEN_12709; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13752 = 3'h4 == tail ? io_op_bits_base_vd_pred : _GEN_12710; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13753 = 3'h5 == tail ? io_op_bits_base_vd_pred : _GEN_12711; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13754 = 3'h6 == tail ? io_op_bits_base_vd_pred : _GEN_12712; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_13755 = 3'h7 == tail ? io_op_bits_base_vd_pred : _GEN_12713; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13756 = 3'h0 == tail ? io_op_bits_base_vd_prec : _GEN_12714; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13757 = 3'h1 == tail ? io_op_bits_base_vd_prec : _GEN_12715; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13758 = 3'h2 == tail ? io_op_bits_base_vd_prec : _GEN_12716; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13759 = 3'h3 == tail ? io_op_bits_base_vd_prec : _GEN_12717; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13760 = 3'h4 == tail ? io_op_bits_base_vd_prec : _GEN_12718; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13761 = 3'h5 == tail ? io_op_bits_base_vd_prec : _GEN_12719; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13762 = 3'h6 == tail ? io_op_bits_base_vd_prec : _GEN_12720; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_13763 = 3'h7 == tail ? io_op_bits_base_vd_prec : _GEN_12721; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_13764 = 3'h0 == tail ? io_op_bits_reg_vd_id : _GEN_12722; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13765 = 3'h1 == tail ? io_op_bits_reg_vd_id : _GEN_12723; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13766 = 3'h2 == tail ? io_op_bits_reg_vd_id : _GEN_12724; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13767 = 3'h3 == tail ? io_op_bits_reg_vd_id : _GEN_12725; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13768 = 3'h4 == tail ? io_op_bits_reg_vd_id : _GEN_12726; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13769 = 3'h5 == tail ? io_op_bits_reg_vd_id : _GEN_12727; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13770 = 3'h6 == tail ? io_op_bits_reg_vd_id : _GEN_12728; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13771 = 3'h7 == tail ? io_op_bits_reg_vd_id : _GEN_12729; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_13772 = io_op_bits_base_vd_valid ? _GEN_13724 : _GEN_12690; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13773 = io_op_bits_base_vd_valid ? _GEN_13725 : _GEN_12691; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13774 = io_op_bits_base_vd_valid ? _GEN_13726 : _GEN_12692; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13775 = io_op_bits_base_vd_valid ? _GEN_13727 : _GEN_12693; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13776 = io_op_bits_base_vd_valid ? _GEN_13728 : _GEN_12694; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13777 = io_op_bits_base_vd_valid ? _GEN_13729 : _GEN_12695; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13778 = io_op_bits_base_vd_valid ? _GEN_13730 : _GEN_12696; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13779 = io_op_bits_base_vd_valid ? _GEN_13731 : _GEN_12697; // @[sequencer-master.scala 362:41]
  wire  _GEN_13780 = io_op_bits_base_vd_valid ? _GEN_13732 : _GEN_12780; // @[sequencer-master.scala 362:41]
  wire  _GEN_13781 = io_op_bits_base_vd_valid ? _GEN_13733 : _GEN_12781; // @[sequencer-master.scala 362:41]
  wire  _GEN_13782 = io_op_bits_base_vd_valid ? _GEN_13734 : _GEN_12782; // @[sequencer-master.scala 362:41]
  wire  _GEN_13783 = io_op_bits_base_vd_valid ? _GEN_13735 : _GEN_12783; // @[sequencer-master.scala 362:41]
  wire  _GEN_13784 = io_op_bits_base_vd_valid ? _GEN_13736 : _GEN_12784; // @[sequencer-master.scala 362:41]
  wire  _GEN_13785 = io_op_bits_base_vd_valid ? _GEN_13737 : _GEN_12785; // @[sequencer-master.scala 362:41]
  wire  _GEN_13786 = io_op_bits_base_vd_valid ? _GEN_13738 : _GEN_12786; // @[sequencer-master.scala 362:41]
  wire  _GEN_13787 = io_op_bits_base_vd_valid ? _GEN_13739 : _GEN_12787; // @[sequencer-master.scala 362:41]
  wire  _GEN_13788 = io_op_bits_base_vd_valid ? _GEN_13740 : _GEN_12698; // @[sequencer-master.scala 362:41]
  wire  _GEN_13789 = io_op_bits_base_vd_valid ? _GEN_13741 : _GEN_12699; // @[sequencer-master.scala 362:41]
  wire  _GEN_13790 = io_op_bits_base_vd_valid ? _GEN_13742 : _GEN_12700; // @[sequencer-master.scala 362:41]
  wire  _GEN_13791 = io_op_bits_base_vd_valid ? _GEN_13743 : _GEN_12701; // @[sequencer-master.scala 362:41]
  wire  _GEN_13792 = io_op_bits_base_vd_valid ? _GEN_13744 : _GEN_12702; // @[sequencer-master.scala 362:41]
  wire  _GEN_13793 = io_op_bits_base_vd_valid ? _GEN_13745 : _GEN_12703; // @[sequencer-master.scala 362:41]
  wire  _GEN_13794 = io_op_bits_base_vd_valid ? _GEN_13746 : _GEN_12704; // @[sequencer-master.scala 362:41]
  wire  _GEN_13795 = io_op_bits_base_vd_valid ? _GEN_13747 : _GEN_12705; // @[sequencer-master.scala 362:41]
  wire  _GEN_13796 = io_op_bits_base_vd_valid ? _GEN_13748 : _GEN_12706; // @[sequencer-master.scala 362:41]
  wire  _GEN_13797 = io_op_bits_base_vd_valid ? _GEN_13749 : _GEN_12707; // @[sequencer-master.scala 362:41]
  wire  _GEN_13798 = io_op_bits_base_vd_valid ? _GEN_13750 : _GEN_12708; // @[sequencer-master.scala 362:41]
  wire  _GEN_13799 = io_op_bits_base_vd_valid ? _GEN_13751 : _GEN_12709; // @[sequencer-master.scala 362:41]
  wire  _GEN_13800 = io_op_bits_base_vd_valid ? _GEN_13752 : _GEN_12710; // @[sequencer-master.scala 362:41]
  wire  _GEN_13801 = io_op_bits_base_vd_valid ? _GEN_13753 : _GEN_12711; // @[sequencer-master.scala 362:41]
  wire  _GEN_13802 = io_op_bits_base_vd_valid ? _GEN_13754 : _GEN_12712; // @[sequencer-master.scala 362:41]
  wire  _GEN_13803 = io_op_bits_base_vd_valid ? _GEN_13755 : _GEN_12713; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13804 = io_op_bits_base_vd_valid ? _GEN_13756 : _GEN_12714; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13805 = io_op_bits_base_vd_valid ? _GEN_13757 : _GEN_12715; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13806 = io_op_bits_base_vd_valid ? _GEN_13758 : _GEN_12716; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13807 = io_op_bits_base_vd_valid ? _GEN_13759 : _GEN_12717; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13808 = io_op_bits_base_vd_valid ? _GEN_13760 : _GEN_12718; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13809 = io_op_bits_base_vd_valid ? _GEN_13761 : _GEN_12719; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13810 = io_op_bits_base_vd_valid ? _GEN_13762 : _GEN_12720; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_13811 = io_op_bits_base_vd_valid ? _GEN_13763 : _GEN_12721; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13812 = io_op_bits_base_vd_valid ? _GEN_13764 : _GEN_12722; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13813 = io_op_bits_base_vd_valid ? _GEN_13765 : _GEN_12723; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13814 = io_op_bits_base_vd_valid ? _GEN_13766 : _GEN_12724; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13815 = io_op_bits_base_vd_valid ? _GEN_13767 : _GEN_12725; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13816 = io_op_bits_base_vd_valid ? _GEN_13768 : _GEN_12726; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13817 = io_op_bits_base_vd_valid ? _GEN_13769 : _GEN_12727; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13818 = io_op_bits_base_vd_valid ? _GEN_13770 : _GEN_12728; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_13819 = io_op_bits_base_vd_valid ? _GEN_13771 : _GEN_12729; // @[sequencer-master.scala 362:41]
  wire  _GEN_13820 = _GEN_32729 | _GEN_12804; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13821 = _GEN_32730 | _GEN_12805; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13822 = _GEN_32731 | _GEN_12806; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13823 = _GEN_32732 | _GEN_12807; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13824 = _GEN_32733 | _GEN_12808; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13825 = _GEN_32734 | _GEN_12809; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13826 = _GEN_32735 | _GEN_12810; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13827 = _GEN_32736 | _GEN_12811; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13828 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13820 : _GEN_12804; // @[sequencer-master.scala 161:86]
  wire  _GEN_13829 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13821 : _GEN_12805; // @[sequencer-master.scala 161:86]
  wire  _GEN_13830 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13822 : _GEN_12806; // @[sequencer-master.scala 161:86]
  wire  _GEN_13831 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13823 : _GEN_12807; // @[sequencer-master.scala 161:86]
  wire  _GEN_13832 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13824 : _GEN_12808; // @[sequencer-master.scala 161:86]
  wire  _GEN_13833 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13825 : _GEN_12809; // @[sequencer-master.scala 161:86]
  wire  _GEN_13834 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13826 : _GEN_12810; // @[sequencer-master.scala 161:86]
  wire  _GEN_13835 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_13827 : _GEN_12811; // @[sequencer-master.scala 161:86]
  wire  _GEN_13836 = _GEN_32729 | _GEN_12828; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13837 = _GEN_32730 | _GEN_12829; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13838 = _GEN_32731 | _GEN_12830; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13839 = _GEN_32732 | _GEN_12831; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13840 = _GEN_32733 | _GEN_12832; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13841 = _GEN_32734 | _GEN_12833; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13842 = _GEN_32735 | _GEN_12834; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13843 = _GEN_32736 | _GEN_12835; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13844 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13836 : _GEN_12828; // @[sequencer-master.scala 161:86]
  wire  _GEN_13845 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13837 : _GEN_12829; // @[sequencer-master.scala 161:86]
  wire  _GEN_13846 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13838 : _GEN_12830; // @[sequencer-master.scala 161:86]
  wire  _GEN_13847 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13839 : _GEN_12831; // @[sequencer-master.scala 161:86]
  wire  _GEN_13848 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13840 : _GEN_12832; // @[sequencer-master.scala 161:86]
  wire  _GEN_13849 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13841 : _GEN_12833; // @[sequencer-master.scala 161:86]
  wire  _GEN_13850 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13842 : _GEN_12834; // @[sequencer-master.scala 161:86]
  wire  _GEN_13851 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_13843 : _GEN_12835; // @[sequencer-master.scala 161:86]
  wire  _GEN_13852 = _GEN_32729 | _GEN_12852; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13853 = _GEN_32730 | _GEN_12853; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13854 = _GEN_32731 | _GEN_12854; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13855 = _GEN_32732 | _GEN_12855; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13856 = _GEN_32733 | _GEN_12856; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13857 = _GEN_32734 | _GEN_12857; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13858 = _GEN_32735 | _GEN_12858; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13859 = _GEN_32736 | _GEN_12859; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13860 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13852 : _GEN_12852; // @[sequencer-master.scala 161:86]
  wire  _GEN_13861 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13853 : _GEN_12853; // @[sequencer-master.scala 161:86]
  wire  _GEN_13862 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13854 : _GEN_12854; // @[sequencer-master.scala 161:86]
  wire  _GEN_13863 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13855 : _GEN_12855; // @[sequencer-master.scala 161:86]
  wire  _GEN_13864 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13856 : _GEN_12856; // @[sequencer-master.scala 161:86]
  wire  _GEN_13865 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13857 : _GEN_12857; // @[sequencer-master.scala 161:86]
  wire  _GEN_13866 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13858 : _GEN_12858; // @[sequencer-master.scala 161:86]
  wire  _GEN_13867 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_13859 : _GEN_12859; // @[sequencer-master.scala 161:86]
  wire  _GEN_13868 = _GEN_32729 | _GEN_12876; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13869 = _GEN_32730 | _GEN_12877; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13870 = _GEN_32731 | _GEN_12878; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13871 = _GEN_32732 | _GEN_12879; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13872 = _GEN_32733 | _GEN_12880; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13873 = _GEN_32734 | _GEN_12881; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13874 = _GEN_32735 | _GEN_12882; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13875 = _GEN_32736 | _GEN_12883; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13876 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13868 : _GEN_12876; // @[sequencer-master.scala 161:86]
  wire  _GEN_13877 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13869 : _GEN_12877; // @[sequencer-master.scala 161:86]
  wire  _GEN_13878 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13870 : _GEN_12878; // @[sequencer-master.scala 161:86]
  wire  _GEN_13879 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13871 : _GEN_12879; // @[sequencer-master.scala 161:86]
  wire  _GEN_13880 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13872 : _GEN_12880; // @[sequencer-master.scala 161:86]
  wire  _GEN_13881 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13873 : _GEN_12881; // @[sequencer-master.scala 161:86]
  wire  _GEN_13882 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13874 : _GEN_12882; // @[sequencer-master.scala 161:86]
  wire  _GEN_13883 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_13875 : _GEN_12883; // @[sequencer-master.scala 161:86]
  wire  _GEN_13884 = _GEN_32729 | _GEN_12900; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13885 = _GEN_32730 | _GEN_12901; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13886 = _GEN_32731 | _GEN_12902; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13887 = _GEN_32732 | _GEN_12903; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13888 = _GEN_32733 | _GEN_12904; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13889 = _GEN_32734 | _GEN_12905; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13890 = _GEN_32735 | _GEN_12906; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13891 = _GEN_32736 | _GEN_12907; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13892 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13884 : _GEN_12900; // @[sequencer-master.scala 161:86]
  wire  _GEN_13893 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13885 : _GEN_12901; // @[sequencer-master.scala 161:86]
  wire  _GEN_13894 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13886 : _GEN_12902; // @[sequencer-master.scala 161:86]
  wire  _GEN_13895 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13887 : _GEN_12903; // @[sequencer-master.scala 161:86]
  wire  _GEN_13896 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13888 : _GEN_12904; // @[sequencer-master.scala 161:86]
  wire  _GEN_13897 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13889 : _GEN_12905; // @[sequencer-master.scala 161:86]
  wire  _GEN_13898 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13890 : _GEN_12906; // @[sequencer-master.scala 161:86]
  wire  _GEN_13899 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_13891 : _GEN_12907; // @[sequencer-master.scala 161:86]
  wire  _GEN_13900 = _GEN_32729 | _GEN_12924; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13901 = _GEN_32730 | _GEN_12925; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13902 = _GEN_32731 | _GEN_12926; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13903 = _GEN_32732 | _GEN_12927; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13904 = _GEN_32733 | _GEN_12928; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13905 = _GEN_32734 | _GEN_12929; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13906 = _GEN_32735 | _GEN_12930; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13907 = _GEN_32736 | _GEN_12931; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13908 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13900 : _GEN_12924; // @[sequencer-master.scala 161:86]
  wire  _GEN_13909 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13901 : _GEN_12925; // @[sequencer-master.scala 161:86]
  wire  _GEN_13910 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13902 : _GEN_12926; // @[sequencer-master.scala 161:86]
  wire  _GEN_13911 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13903 : _GEN_12927; // @[sequencer-master.scala 161:86]
  wire  _GEN_13912 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13904 : _GEN_12928; // @[sequencer-master.scala 161:86]
  wire  _GEN_13913 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13905 : _GEN_12929; // @[sequencer-master.scala 161:86]
  wire  _GEN_13914 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13906 : _GEN_12930; // @[sequencer-master.scala 161:86]
  wire  _GEN_13915 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_13907 : _GEN_12931; // @[sequencer-master.scala 161:86]
  wire  _GEN_13916 = _GEN_32729 | _GEN_12948; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13917 = _GEN_32730 | _GEN_12949; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13918 = _GEN_32731 | _GEN_12950; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13919 = _GEN_32732 | _GEN_12951; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13920 = _GEN_32733 | _GEN_12952; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13921 = _GEN_32734 | _GEN_12953; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13922 = _GEN_32735 | _GEN_12954; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13923 = _GEN_32736 | _GEN_12955; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13924 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13916 : _GEN_12948; // @[sequencer-master.scala 161:86]
  wire  _GEN_13925 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13917 : _GEN_12949; // @[sequencer-master.scala 161:86]
  wire  _GEN_13926 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13918 : _GEN_12950; // @[sequencer-master.scala 161:86]
  wire  _GEN_13927 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13919 : _GEN_12951; // @[sequencer-master.scala 161:86]
  wire  _GEN_13928 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13920 : _GEN_12952; // @[sequencer-master.scala 161:86]
  wire  _GEN_13929 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13921 : _GEN_12953; // @[sequencer-master.scala 161:86]
  wire  _GEN_13930 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13922 : _GEN_12954; // @[sequencer-master.scala 161:86]
  wire  _GEN_13931 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_13923 : _GEN_12955; // @[sequencer-master.scala 161:86]
  wire  _GEN_13932 = _GEN_32729 | _GEN_12972; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13933 = _GEN_32730 | _GEN_12973; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13934 = _GEN_32731 | _GEN_12974; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13935 = _GEN_32732 | _GEN_12975; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13936 = _GEN_32733 | _GEN_12976; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13937 = _GEN_32734 | _GEN_12977; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13938 = _GEN_32735 | _GEN_12978; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13939 = _GEN_32736 | _GEN_12979; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_13940 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13932 : _GEN_12972; // @[sequencer-master.scala 161:86]
  wire  _GEN_13941 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13933 : _GEN_12973; // @[sequencer-master.scala 161:86]
  wire  _GEN_13942 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13934 : _GEN_12974; // @[sequencer-master.scala 161:86]
  wire  _GEN_13943 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13935 : _GEN_12975; // @[sequencer-master.scala 161:86]
  wire  _GEN_13944 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13936 : _GEN_12976; // @[sequencer-master.scala 161:86]
  wire  _GEN_13945 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13937 : _GEN_12977; // @[sequencer-master.scala 161:86]
  wire  _GEN_13946 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13938 : _GEN_12978; // @[sequencer-master.scala 161:86]
  wire  _GEN_13947 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_13939 : _GEN_12979; // @[sequencer-master.scala 161:86]
  wire  _GEN_13948 = _GEN_32729 | _GEN_12812; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13949 = _GEN_32730 | _GEN_12813; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13950 = _GEN_32731 | _GEN_12814; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13951 = _GEN_32732 | _GEN_12815; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13952 = _GEN_32733 | _GEN_12816; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13953 = _GEN_32734 | _GEN_12817; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13954 = _GEN_32735 | _GEN_12818; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13955 = _GEN_32736 | _GEN_12819; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13956 = _T_1442 ? _GEN_13948 : _GEN_12812; // @[sequencer-master.scala 168:32]
  wire  _GEN_13957 = _T_1442 ? _GEN_13949 : _GEN_12813; // @[sequencer-master.scala 168:32]
  wire  _GEN_13958 = _T_1442 ? _GEN_13950 : _GEN_12814; // @[sequencer-master.scala 168:32]
  wire  _GEN_13959 = _T_1442 ? _GEN_13951 : _GEN_12815; // @[sequencer-master.scala 168:32]
  wire  _GEN_13960 = _T_1442 ? _GEN_13952 : _GEN_12816; // @[sequencer-master.scala 168:32]
  wire  _GEN_13961 = _T_1442 ? _GEN_13953 : _GEN_12817; // @[sequencer-master.scala 168:32]
  wire  _GEN_13962 = _T_1442 ? _GEN_13954 : _GEN_12818; // @[sequencer-master.scala 168:32]
  wire  _GEN_13963 = _T_1442 ? _GEN_13955 : _GEN_12819; // @[sequencer-master.scala 168:32]
  wire  _GEN_13964 = _GEN_32729 | _GEN_12836; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13965 = _GEN_32730 | _GEN_12837; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13966 = _GEN_32731 | _GEN_12838; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13967 = _GEN_32732 | _GEN_12839; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13968 = _GEN_32733 | _GEN_12840; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13969 = _GEN_32734 | _GEN_12841; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13970 = _GEN_32735 | _GEN_12842; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13971 = _GEN_32736 | _GEN_12843; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13972 = _T_1464 ? _GEN_13964 : _GEN_12836; // @[sequencer-master.scala 168:32]
  wire  _GEN_13973 = _T_1464 ? _GEN_13965 : _GEN_12837; // @[sequencer-master.scala 168:32]
  wire  _GEN_13974 = _T_1464 ? _GEN_13966 : _GEN_12838; // @[sequencer-master.scala 168:32]
  wire  _GEN_13975 = _T_1464 ? _GEN_13967 : _GEN_12839; // @[sequencer-master.scala 168:32]
  wire  _GEN_13976 = _T_1464 ? _GEN_13968 : _GEN_12840; // @[sequencer-master.scala 168:32]
  wire  _GEN_13977 = _T_1464 ? _GEN_13969 : _GEN_12841; // @[sequencer-master.scala 168:32]
  wire  _GEN_13978 = _T_1464 ? _GEN_13970 : _GEN_12842; // @[sequencer-master.scala 168:32]
  wire  _GEN_13979 = _T_1464 ? _GEN_13971 : _GEN_12843; // @[sequencer-master.scala 168:32]
  wire  _GEN_13980 = _GEN_32729 | _GEN_12860; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13981 = _GEN_32730 | _GEN_12861; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13982 = _GEN_32731 | _GEN_12862; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13983 = _GEN_32732 | _GEN_12863; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13984 = _GEN_32733 | _GEN_12864; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13985 = _GEN_32734 | _GEN_12865; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13986 = _GEN_32735 | _GEN_12866; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13987 = _GEN_32736 | _GEN_12867; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13988 = _T_1486 ? _GEN_13980 : _GEN_12860; // @[sequencer-master.scala 168:32]
  wire  _GEN_13989 = _T_1486 ? _GEN_13981 : _GEN_12861; // @[sequencer-master.scala 168:32]
  wire  _GEN_13990 = _T_1486 ? _GEN_13982 : _GEN_12862; // @[sequencer-master.scala 168:32]
  wire  _GEN_13991 = _T_1486 ? _GEN_13983 : _GEN_12863; // @[sequencer-master.scala 168:32]
  wire  _GEN_13992 = _T_1486 ? _GEN_13984 : _GEN_12864; // @[sequencer-master.scala 168:32]
  wire  _GEN_13993 = _T_1486 ? _GEN_13985 : _GEN_12865; // @[sequencer-master.scala 168:32]
  wire  _GEN_13994 = _T_1486 ? _GEN_13986 : _GEN_12866; // @[sequencer-master.scala 168:32]
  wire  _GEN_13995 = _T_1486 ? _GEN_13987 : _GEN_12867; // @[sequencer-master.scala 168:32]
  wire  _GEN_13996 = _GEN_32729 | _GEN_12884; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13997 = _GEN_32730 | _GEN_12885; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13998 = _GEN_32731 | _GEN_12886; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_13999 = _GEN_32732 | _GEN_12887; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14000 = _GEN_32733 | _GEN_12888; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14001 = _GEN_32734 | _GEN_12889; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14002 = _GEN_32735 | _GEN_12890; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14003 = _GEN_32736 | _GEN_12891; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14004 = _T_1508 ? _GEN_13996 : _GEN_12884; // @[sequencer-master.scala 168:32]
  wire  _GEN_14005 = _T_1508 ? _GEN_13997 : _GEN_12885; // @[sequencer-master.scala 168:32]
  wire  _GEN_14006 = _T_1508 ? _GEN_13998 : _GEN_12886; // @[sequencer-master.scala 168:32]
  wire  _GEN_14007 = _T_1508 ? _GEN_13999 : _GEN_12887; // @[sequencer-master.scala 168:32]
  wire  _GEN_14008 = _T_1508 ? _GEN_14000 : _GEN_12888; // @[sequencer-master.scala 168:32]
  wire  _GEN_14009 = _T_1508 ? _GEN_14001 : _GEN_12889; // @[sequencer-master.scala 168:32]
  wire  _GEN_14010 = _T_1508 ? _GEN_14002 : _GEN_12890; // @[sequencer-master.scala 168:32]
  wire  _GEN_14011 = _T_1508 ? _GEN_14003 : _GEN_12891; // @[sequencer-master.scala 168:32]
  wire  _GEN_14012 = _GEN_32729 | _GEN_12908; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14013 = _GEN_32730 | _GEN_12909; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14014 = _GEN_32731 | _GEN_12910; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14015 = _GEN_32732 | _GEN_12911; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14016 = _GEN_32733 | _GEN_12912; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14017 = _GEN_32734 | _GEN_12913; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14018 = _GEN_32735 | _GEN_12914; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14019 = _GEN_32736 | _GEN_12915; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14020 = _T_1530 ? _GEN_14012 : _GEN_12908; // @[sequencer-master.scala 168:32]
  wire  _GEN_14021 = _T_1530 ? _GEN_14013 : _GEN_12909; // @[sequencer-master.scala 168:32]
  wire  _GEN_14022 = _T_1530 ? _GEN_14014 : _GEN_12910; // @[sequencer-master.scala 168:32]
  wire  _GEN_14023 = _T_1530 ? _GEN_14015 : _GEN_12911; // @[sequencer-master.scala 168:32]
  wire  _GEN_14024 = _T_1530 ? _GEN_14016 : _GEN_12912; // @[sequencer-master.scala 168:32]
  wire  _GEN_14025 = _T_1530 ? _GEN_14017 : _GEN_12913; // @[sequencer-master.scala 168:32]
  wire  _GEN_14026 = _T_1530 ? _GEN_14018 : _GEN_12914; // @[sequencer-master.scala 168:32]
  wire  _GEN_14027 = _T_1530 ? _GEN_14019 : _GEN_12915; // @[sequencer-master.scala 168:32]
  wire  _GEN_14028 = _GEN_32729 | _GEN_12932; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14029 = _GEN_32730 | _GEN_12933; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14030 = _GEN_32731 | _GEN_12934; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14031 = _GEN_32732 | _GEN_12935; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14032 = _GEN_32733 | _GEN_12936; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14033 = _GEN_32734 | _GEN_12937; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14034 = _GEN_32735 | _GEN_12938; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14035 = _GEN_32736 | _GEN_12939; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14036 = _T_1552 ? _GEN_14028 : _GEN_12932; // @[sequencer-master.scala 168:32]
  wire  _GEN_14037 = _T_1552 ? _GEN_14029 : _GEN_12933; // @[sequencer-master.scala 168:32]
  wire  _GEN_14038 = _T_1552 ? _GEN_14030 : _GEN_12934; // @[sequencer-master.scala 168:32]
  wire  _GEN_14039 = _T_1552 ? _GEN_14031 : _GEN_12935; // @[sequencer-master.scala 168:32]
  wire  _GEN_14040 = _T_1552 ? _GEN_14032 : _GEN_12936; // @[sequencer-master.scala 168:32]
  wire  _GEN_14041 = _T_1552 ? _GEN_14033 : _GEN_12937; // @[sequencer-master.scala 168:32]
  wire  _GEN_14042 = _T_1552 ? _GEN_14034 : _GEN_12938; // @[sequencer-master.scala 168:32]
  wire  _GEN_14043 = _T_1552 ? _GEN_14035 : _GEN_12939; // @[sequencer-master.scala 168:32]
  wire  _GEN_14044 = _GEN_32729 | _GEN_12956; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14045 = _GEN_32730 | _GEN_12957; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14046 = _GEN_32731 | _GEN_12958; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14047 = _GEN_32732 | _GEN_12959; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14048 = _GEN_32733 | _GEN_12960; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14049 = _GEN_32734 | _GEN_12961; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14050 = _GEN_32735 | _GEN_12962; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14051 = _GEN_32736 | _GEN_12963; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14052 = _T_1574 ? _GEN_14044 : _GEN_12956; // @[sequencer-master.scala 168:32]
  wire  _GEN_14053 = _T_1574 ? _GEN_14045 : _GEN_12957; // @[sequencer-master.scala 168:32]
  wire  _GEN_14054 = _T_1574 ? _GEN_14046 : _GEN_12958; // @[sequencer-master.scala 168:32]
  wire  _GEN_14055 = _T_1574 ? _GEN_14047 : _GEN_12959; // @[sequencer-master.scala 168:32]
  wire  _GEN_14056 = _T_1574 ? _GEN_14048 : _GEN_12960; // @[sequencer-master.scala 168:32]
  wire  _GEN_14057 = _T_1574 ? _GEN_14049 : _GEN_12961; // @[sequencer-master.scala 168:32]
  wire  _GEN_14058 = _T_1574 ? _GEN_14050 : _GEN_12962; // @[sequencer-master.scala 168:32]
  wire  _GEN_14059 = _T_1574 ? _GEN_14051 : _GEN_12963; // @[sequencer-master.scala 168:32]
  wire  _GEN_14060 = _GEN_32729 | _GEN_12980; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14061 = _GEN_32730 | _GEN_12981; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14062 = _GEN_32731 | _GEN_12982; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14063 = _GEN_32732 | _GEN_12983; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14064 = _GEN_32733 | _GEN_12984; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14065 = _GEN_32734 | _GEN_12985; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14066 = _GEN_32735 | _GEN_12986; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14067 = _GEN_32736 | _GEN_12987; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_14068 = _T_1596 ? _GEN_14060 : _GEN_12980; // @[sequencer-master.scala 168:32]
  wire  _GEN_14069 = _T_1596 ? _GEN_14061 : _GEN_12981; // @[sequencer-master.scala 168:32]
  wire  _GEN_14070 = _T_1596 ? _GEN_14062 : _GEN_12982; // @[sequencer-master.scala 168:32]
  wire  _GEN_14071 = _T_1596 ? _GEN_14063 : _GEN_12983; // @[sequencer-master.scala 168:32]
  wire  _GEN_14072 = _T_1596 ? _GEN_14064 : _GEN_12984; // @[sequencer-master.scala 168:32]
  wire  _GEN_14073 = _T_1596 ? _GEN_14065 : _GEN_12985; // @[sequencer-master.scala 168:32]
  wire  _GEN_14074 = _T_1596 ? _GEN_14066 : _GEN_12986; // @[sequencer-master.scala 168:32]
  wire  _GEN_14075 = _T_1596 ? _GEN_14067 : _GEN_12987; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_14076 = 3'h0 == tail ? _T_1615[1:0] : _GEN_12658; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14077 = 3'h1 == tail ? _T_1615[1:0] : _GEN_12659; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14078 = 3'h2 == tail ? _T_1615[1:0] : _GEN_12660; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14079 = 3'h3 == tail ? _T_1615[1:0] : _GEN_12661; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14080 = 3'h4 == tail ? _T_1615[1:0] : _GEN_12662; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14081 = 3'h5 == tail ? _T_1615[1:0] : _GEN_12663; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14082 = 3'h6 == tail ? _T_1615[1:0] : _GEN_12664; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_14083 = 3'h7 == tail ? _T_1615[1:0] : _GEN_12665; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_14084 = 3'h0 == tail ? 4'h0 : _GEN_12666; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14085 = 3'h1 == tail ? 4'h0 : _GEN_12667; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14086 = 3'h2 == tail ? 4'h0 : _GEN_12668; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14087 = 3'h3 == tail ? 4'h0 : _GEN_12669; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14088 = 3'h4 == tail ? 4'h0 : _GEN_12670; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14089 = 3'h5 == tail ? 4'h0 : _GEN_12671; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14090 = 3'h6 == tail ? 4'h0 : _GEN_12672; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_14091 = 3'h7 == tail ? 4'h0 : _GEN_12673; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_14092 = 3'h0 == tail ? 3'h0 : _GEN_12674; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14093 = 3'h1 == tail ? 3'h0 : _GEN_12675; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14094 = 3'h2 == tail ? 3'h0 : _GEN_12676; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14095 = 3'h3 == tail ? 3'h0 : _GEN_12677; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14096 = 3'h4 == tail ? 3'h0 : _GEN_12678; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14097 = 3'h5 == tail ? 3'h0 : _GEN_12679; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14098 = 3'h6 == tail ? 3'h0 : _GEN_12680; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_14099 = 3'h7 == tail ? 3'h0 : _GEN_12681; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [3:0] _GEN_14100 = 3'h0 == tail ? _T_1792 : _GEN_14084; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14101 = 3'h1 == tail ? _T_1792 : _GEN_14085; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14102 = 3'h2 == tail ? _T_1792 : _GEN_14086; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14103 = 3'h3 == tail ? _T_1792 : _GEN_14087; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14104 = 3'h4 == tail ? _T_1792 : _GEN_14088; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14105 = 3'h5 == tail ? _T_1792 : _GEN_14089; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14106 = 3'h6 == tail ? _T_1792 : _GEN_14090; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14107 = 3'h7 == tail ? _T_1792 : _GEN_14091; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_14108 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14100 : _GEN_14084; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14109 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14101 : _GEN_14085; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14110 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14102 : _GEN_14086; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14111 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14103 : _GEN_14087; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14112 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14104 : _GEN_14088; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14113 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14105 : _GEN_14089; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14114 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14106 : _GEN_14090; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_14115 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_14107 : _GEN_14091; // @[sequencer-master.scala 235:47]
  wire [2:0] _GEN_14116 = 3'h0 == tail ? _T_1792[2:0] : _GEN_14092; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14117 = 3'h1 == tail ? _T_1792[2:0] : _GEN_14093; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14118 = 3'h2 == tail ? _T_1792[2:0] : _GEN_14094; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14119 = 3'h3 == tail ? _T_1792[2:0] : _GEN_14095; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14120 = 3'h4 == tail ? _T_1792[2:0] : _GEN_14096; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14121 = 3'h5 == tail ? _T_1792[2:0] : _GEN_14097; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14122 = 3'h6 == tail ? _T_1792[2:0] : _GEN_14098; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14123 = 3'h7 == tail ? _T_1792[2:0] : _GEN_14099; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_14124 = io_op_bits_base_vd_pred ? _GEN_14116 : _GEN_14092; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14125 = io_op_bits_base_vd_pred ? _GEN_14117 : _GEN_14093; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14126 = io_op_bits_base_vd_pred ? _GEN_14118 : _GEN_14094; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14127 = io_op_bits_base_vd_pred ? _GEN_14119 : _GEN_14095; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14128 = io_op_bits_base_vd_pred ? _GEN_14120 : _GEN_14096; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14129 = io_op_bits_base_vd_pred ? _GEN_14121 : _GEN_14097; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14130 = io_op_bits_base_vd_pred ? _GEN_14122 : _GEN_14098; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_14131 = io_op_bits_base_vd_pred ? _GEN_14123 : _GEN_14099; // @[sequencer-master.scala 236:45]
  wire  _GEN_14132 = io_op_bits_active_vfcmp ? _GEN_12732 : _GEN_12242; // @[sequencer-master.scala 646:40]
  wire  _GEN_14133 = io_op_bits_active_vfcmp ? _GEN_12733 : _GEN_12243; // @[sequencer-master.scala 646:40]
  wire  _GEN_14134 = io_op_bits_active_vfcmp ? _GEN_12734 : _GEN_12244; // @[sequencer-master.scala 646:40]
  wire  _GEN_14135 = io_op_bits_active_vfcmp ? _GEN_12735 : _GEN_12245; // @[sequencer-master.scala 646:40]
  wire  _GEN_14136 = io_op_bits_active_vfcmp ? _GEN_12736 : _GEN_12246; // @[sequencer-master.scala 646:40]
  wire  _GEN_14137 = io_op_bits_active_vfcmp ? _GEN_12737 : _GEN_12247; // @[sequencer-master.scala 646:40]
  wire  _GEN_14138 = io_op_bits_active_vfcmp ? _GEN_12738 : _GEN_12248; // @[sequencer-master.scala 646:40]
  wire  _GEN_14139 = io_op_bits_active_vfcmp ? _GEN_12739 : _GEN_12249; // @[sequencer-master.scala 646:40]
  wire  _GEN_14148 = io_op_bits_active_vfcmp ? _GEN_13068 : _GEN_12258; // @[sequencer-master.scala 646:40]
  wire  _GEN_14149 = io_op_bits_active_vfcmp ? _GEN_13069 : _GEN_12259; // @[sequencer-master.scala 646:40]
  wire  _GEN_14150 = io_op_bits_active_vfcmp ? _GEN_13070 : _GEN_12260; // @[sequencer-master.scala 646:40]
  wire  _GEN_14151 = io_op_bits_active_vfcmp ? _GEN_13071 : _GEN_12261; // @[sequencer-master.scala 646:40]
  wire  _GEN_14152 = io_op_bits_active_vfcmp ? _GEN_13072 : _GEN_12262; // @[sequencer-master.scala 646:40]
  wire  _GEN_14153 = io_op_bits_active_vfcmp ? _GEN_13073 : _GEN_12263; // @[sequencer-master.scala 646:40]
  wire  _GEN_14154 = io_op_bits_active_vfcmp ? _GEN_13074 : _GEN_12264; // @[sequencer-master.scala 646:40]
  wire  _GEN_14155 = io_op_bits_active_vfcmp ? _GEN_13075 : _GEN_12265; // @[sequencer-master.scala 646:40]
  wire  _GEN_14156 = io_op_bits_active_vfcmp ? _GEN_13300 : _GEN_12266; // @[sequencer-master.scala 646:40]
  wire  _GEN_14157 = io_op_bits_active_vfcmp ? _GEN_13301 : _GEN_12267; // @[sequencer-master.scala 646:40]
  wire  _GEN_14158 = io_op_bits_active_vfcmp ? _GEN_13302 : _GEN_12268; // @[sequencer-master.scala 646:40]
  wire  _GEN_14159 = io_op_bits_active_vfcmp ? _GEN_13303 : _GEN_12269; // @[sequencer-master.scala 646:40]
  wire  _GEN_14160 = io_op_bits_active_vfcmp ? _GEN_13304 : _GEN_12270; // @[sequencer-master.scala 646:40]
  wire  _GEN_14161 = io_op_bits_active_vfcmp ? _GEN_13305 : _GEN_12271; // @[sequencer-master.scala 646:40]
  wire  _GEN_14162 = io_op_bits_active_vfcmp ? _GEN_13306 : _GEN_12272; // @[sequencer-master.scala 646:40]
  wire  _GEN_14163 = io_op_bits_active_vfcmp ? _GEN_13307 : _GEN_12273; // @[sequencer-master.scala 646:40]
  wire  _GEN_14164 = io_op_bits_active_vfcmp ? _GEN_13548 : _GEN_12274; // @[sequencer-master.scala 646:40]
  wire  _GEN_14165 = io_op_bits_active_vfcmp ? _GEN_13549 : _GEN_12275; // @[sequencer-master.scala 646:40]
  wire  _GEN_14166 = io_op_bits_active_vfcmp ? _GEN_13550 : _GEN_12276; // @[sequencer-master.scala 646:40]
  wire  _GEN_14167 = io_op_bits_active_vfcmp ? _GEN_13551 : _GEN_12277; // @[sequencer-master.scala 646:40]
  wire  _GEN_14168 = io_op_bits_active_vfcmp ? _GEN_13552 : _GEN_12278; // @[sequencer-master.scala 646:40]
  wire  _GEN_14169 = io_op_bits_active_vfcmp ? _GEN_13553 : _GEN_12279; // @[sequencer-master.scala 646:40]
  wire  _GEN_14170 = io_op_bits_active_vfcmp ? _GEN_13554 : _GEN_12280; // @[sequencer-master.scala 646:40]
  wire  _GEN_14171 = io_op_bits_active_vfcmp ? _GEN_13555 : _GEN_12281; // @[sequencer-master.scala 646:40]
  wire  _GEN_14172 = io_op_bits_active_vfcmp ? _GEN_12772 : _GEN_12282; // @[sequencer-master.scala 646:40]
  wire  _GEN_14173 = io_op_bits_active_vfcmp ? _GEN_12773 : _GEN_12283; // @[sequencer-master.scala 646:40]
  wire  _GEN_14174 = io_op_bits_active_vfcmp ? _GEN_12774 : _GEN_12284; // @[sequencer-master.scala 646:40]
  wire  _GEN_14175 = io_op_bits_active_vfcmp ? _GEN_12775 : _GEN_12285; // @[sequencer-master.scala 646:40]
  wire  _GEN_14176 = io_op_bits_active_vfcmp ? _GEN_12776 : _GEN_12286; // @[sequencer-master.scala 646:40]
  wire  _GEN_14177 = io_op_bits_active_vfcmp ? _GEN_12777 : _GEN_12287; // @[sequencer-master.scala 646:40]
  wire  _GEN_14178 = io_op_bits_active_vfcmp ? _GEN_12778 : _GEN_12288; // @[sequencer-master.scala 646:40]
  wire  _GEN_14179 = io_op_bits_active_vfcmp ? _GEN_12779 : _GEN_12289; // @[sequencer-master.scala 646:40]
  wire  _GEN_14180 = io_op_bits_active_vfcmp ? _GEN_13780 : _GEN_12290; // @[sequencer-master.scala 646:40]
  wire  _GEN_14181 = io_op_bits_active_vfcmp ? _GEN_13781 : _GEN_12291; // @[sequencer-master.scala 646:40]
  wire  _GEN_14182 = io_op_bits_active_vfcmp ? _GEN_13782 : _GEN_12292; // @[sequencer-master.scala 646:40]
  wire  _GEN_14183 = io_op_bits_active_vfcmp ? _GEN_13783 : _GEN_12293; // @[sequencer-master.scala 646:40]
  wire  _GEN_14184 = io_op_bits_active_vfcmp ? _GEN_13784 : _GEN_12294; // @[sequencer-master.scala 646:40]
  wire  _GEN_14185 = io_op_bits_active_vfcmp ? _GEN_13785 : _GEN_12295; // @[sequencer-master.scala 646:40]
  wire  _GEN_14186 = io_op_bits_active_vfcmp ? _GEN_13786 : _GEN_12296; // @[sequencer-master.scala 646:40]
  wire  _GEN_14187 = io_op_bits_active_vfcmp ? _GEN_13787 : _GEN_12297; // @[sequencer-master.scala 646:40]
  wire  _GEN_14188 = io_op_bits_active_vfcmp ? _GEN_12788 : _GEN_12298; // @[sequencer-master.scala 646:40]
  wire  _GEN_14189 = io_op_bits_active_vfcmp ? _GEN_12789 : _GEN_12299; // @[sequencer-master.scala 646:40]
  wire  _GEN_14190 = io_op_bits_active_vfcmp ? _GEN_12790 : _GEN_12300; // @[sequencer-master.scala 646:40]
  wire  _GEN_14191 = io_op_bits_active_vfcmp ? _GEN_12791 : _GEN_12301; // @[sequencer-master.scala 646:40]
  wire  _GEN_14192 = io_op_bits_active_vfcmp ? _GEN_12792 : _GEN_12302; // @[sequencer-master.scala 646:40]
  wire  _GEN_14193 = io_op_bits_active_vfcmp ? _GEN_12793 : _GEN_12303; // @[sequencer-master.scala 646:40]
  wire  _GEN_14194 = io_op_bits_active_vfcmp ? _GEN_12794 : _GEN_12304; // @[sequencer-master.scala 646:40]
  wire  _GEN_14195 = io_op_bits_active_vfcmp ? _GEN_12795 : _GEN_12305; // @[sequencer-master.scala 646:40]
  wire  _GEN_14196 = io_op_bits_active_vfcmp ? _GEN_13604 : _GEN_12306; // @[sequencer-master.scala 646:40]
  wire  _GEN_14197 = io_op_bits_active_vfcmp ? _GEN_13605 : _GEN_12307; // @[sequencer-master.scala 646:40]
  wire  _GEN_14198 = io_op_bits_active_vfcmp ? _GEN_13606 : _GEN_12308; // @[sequencer-master.scala 646:40]
  wire  _GEN_14199 = io_op_bits_active_vfcmp ? _GEN_13607 : _GEN_12309; // @[sequencer-master.scala 646:40]
  wire  _GEN_14200 = io_op_bits_active_vfcmp ? _GEN_13608 : _GEN_12310; // @[sequencer-master.scala 646:40]
  wire  _GEN_14201 = io_op_bits_active_vfcmp ? _GEN_13609 : _GEN_12311; // @[sequencer-master.scala 646:40]
  wire  _GEN_14202 = io_op_bits_active_vfcmp ? _GEN_13610 : _GEN_12312; // @[sequencer-master.scala 646:40]
  wire  _GEN_14203 = io_op_bits_active_vfcmp ? _GEN_13611 : _GEN_12313; // @[sequencer-master.scala 646:40]
  wire  _GEN_14204 = io_op_bits_active_vfcmp ? _GEN_13828 : _GEN_12314; // @[sequencer-master.scala 646:40]
  wire  _GEN_14205 = io_op_bits_active_vfcmp ? _GEN_13829 : _GEN_12315; // @[sequencer-master.scala 646:40]
  wire  _GEN_14206 = io_op_bits_active_vfcmp ? _GEN_13830 : _GEN_12316; // @[sequencer-master.scala 646:40]
  wire  _GEN_14207 = io_op_bits_active_vfcmp ? _GEN_13831 : _GEN_12317; // @[sequencer-master.scala 646:40]
  wire  _GEN_14208 = io_op_bits_active_vfcmp ? _GEN_13832 : _GEN_12318; // @[sequencer-master.scala 646:40]
  wire  _GEN_14209 = io_op_bits_active_vfcmp ? _GEN_13833 : _GEN_12319; // @[sequencer-master.scala 646:40]
  wire  _GEN_14210 = io_op_bits_active_vfcmp ? _GEN_13834 : _GEN_12320; // @[sequencer-master.scala 646:40]
  wire  _GEN_14211 = io_op_bits_active_vfcmp ? _GEN_13835 : _GEN_12321; // @[sequencer-master.scala 646:40]
  wire  _GEN_14212 = io_op_bits_active_vfcmp ? _GEN_13956 : _GEN_12322; // @[sequencer-master.scala 646:40]
  wire  _GEN_14213 = io_op_bits_active_vfcmp ? _GEN_13957 : _GEN_12323; // @[sequencer-master.scala 646:40]
  wire  _GEN_14214 = io_op_bits_active_vfcmp ? _GEN_13958 : _GEN_12324; // @[sequencer-master.scala 646:40]
  wire  _GEN_14215 = io_op_bits_active_vfcmp ? _GEN_13959 : _GEN_12325; // @[sequencer-master.scala 646:40]
  wire  _GEN_14216 = io_op_bits_active_vfcmp ? _GEN_13960 : _GEN_12326; // @[sequencer-master.scala 646:40]
  wire  _GEN_14217 = io_op_bits_active_vfcmp ? _GEN_13961 : _GEN_12327; // @[sequencer-master.scala 646:40]
  wire  _GEN_14218 = io_op_bits_active_vfcmp ? _GEN_13962 : _GEN_12328; // @[sequencer-master.scala 646:40]
  wire  _GEN_14219 = io_op_bits_active_vfcmp ? _GEN_13963 : _GEN_12329; // @[sequencer-master.scala 646:40]
  wire  _GEN_14220 = io_op_bits_active_vfcmp ? _GEN_13620 : _GEN_12330; // @[sequencer-master.scala 646:40]
  wire  _GEN_14221 = io_op_bits_active_vfcmp ? _GEN_13621 : _GEN_12331; // @[sequencer-master.scala 646:40]
  wire  _GEN_14222 = io_op_bits_active_vfcmp ? _GEN_13622 : _GEN_12332; // @[sequencer-master.scala 646:40]
  wire  _GEN_14223 = io_op_bits_active_vfcmp ? _GEN_13623 : _GEN_12333; // @[sequencer-master.scala 646:40]
  wire  _GEN_14224 = io_op_bits_active_vfcmp ? _GEN_13624 : _GEN_12334; // @[sequencer-master.scala 646:40]
  wire  _GEN_14225 = io_op_bits_active_vfcmp ? _GEN_13625 : _GEN_12335; // @[sequencer-master.scala 646:40]
  wire  _GEN_14226 = io_op_bits_active_vfcmp ? _GEN_13626 : _GEN_12336; // @[sequencer-master.scala 646:40]
  wire  _GEN_14227 = io_op_bits_active_vfcmp ? _GEN_13627 : _GEN_12337; // @[sequencer-master.scala 646:40]
  wire  _GEN_14228 = io_op_bits_active_vfcmp ? _GEN_13844 : _GEN_12338; // @[sequencer-master.scala 646:40]
  wire  _GEN_14229 = io_op_bits_active_vfcmp ? _GEN_13845 : _GEN_12339; // @[sequencer-master.scala 646:40]
  wire  _GEN_14230 = io_op_bits_active_vfcmp ? _GEN_13846 : _GEN_12340; // @[sequencer-master.scala 646:40]
  wire  _GEN_14231 = io_op_bits_active_vfcmp ? _GEN_13847 : _GEN_12341; // @[sequencer-master.scala 646:40]
  wire  _GEN_14232 = io_op_bits_active_vfcmp ? _GEN_13848 : _GEN_12342; // @[sequencer-master.scala 646:40]
  wire  _GEN_14233 = io_op_bits_active_vfcmp ? _GEN_13849 : _GEN_12343; // @[sequencer-master.scala 646:40]
  wire  _GEN_14234 = io_op_bits_active_vfcmp ? _GEN_13850 : _GEN_12344; // @[sequencer-master.scala 646:40]
  wire  _GEN_14235 = io_op_bits_active_vfcmp ? _GEN_13851 : _GEN_12345; // @[sequencer-master.scala 646:40]
  wire  _GEN_14236 = io_op_bits_active_vfcmp ? _GEN_13972 : _GEN_12346; // @[sequencer-master.scala 646:40]
  wire  _GEN_14237 = io_op_bits_active_vfcmp ? _GEN_13973 : _GEN_12347; // @[sequencer-master.scala 646:40]
  wire  _GEN_14238 = io_op_bits_active_vfcmp ? _GEN_13974 : _GEN_12348; // @[sequencer-master.scala 646:40]
  wire  _GEN_14239 = io_op_bits_active_vfcmp ? _GEN_13975 : _GEN_12349; // @[sequencer-master.scala 646:40]
  wire  _GEN_14240 = io_op_bits_active_vfcmp ? _GEN_13976 : _GEN_12350; // @[sequencer-master.scala 646:40]
  wire  _GEN_14241 = io_op_bits_active_vfcmp ? _GEN_13977 : _GEN_12351; // @[sequencer-master.scala 646:40]
  wire  _GEN_14242 = io_op_bits_active_vfcmp ? _GEN_13978 : _GEN_12352; // @[sequencer-master.scala 646:40]
  wire  _GEN_14243 = io_op_bits_active_vfcmp ? _GEN_13979 : _GEN_12353; // @[sequencer-master.scala 646:40]
  wire  _GEN_14244 = io_op_bits_active_vfcmp ? _GEN_13636 : _GEN_12354; // @[sequencer-master.scala 646:40]
  wire  _GEN_14245 = io_op_bits_active_vfcmp ? _GEN_13637 : _GEN_12355; // @[sequencer-master.scala 646:40]
  wire  _GEN_14246 = io_op_bits_active_vfcmp ? _GEN_13638 : _GEN_12356; // @[sequencer-master.scala 646:40]
  wire  _GEN_14247 = io_op_bits_active_vfcmp ? _GEN_13639 : _GEN_12357; // @[sequencer-master.scala 646:40]
  wire  _GEN_14248 = io_op_bits_active_vfcmp ? _GEN_13640 : _GEN_12358; // @[sequencer-master.scala 646:40]
  wire  _GEN_14249 = io_op_bits_active_vfcmp ? _GEN_13641 : _GEN_12359; // @[sequencer-master.scala 646:40]
  wire  _GEN_14250 = io_op_bits_active_vfcmp ? _GEN_13642 : _GEN_12360; // @[sequencer-master.scala 646:40]
  wire  _GEN_14251 = io_op_bits_active_vfcmp ? _GEN_13643 : _GEN_12361; // @[sequencer-master.scala 646:40]
  wire  _GEN_14252 = io_op_bits_active_vfcmp ? _GEN_13860 : _GEN_12362; // @[sequencer-master.scala 646:40]
  wire  _GEN_14253 = io_op_bits_active_vfcmp ? _GEN_13861 : _GEN_12363; // @[sequencer-master.scala 646:40]
  wire  _GEN_14254 = io_op_bits_active_vfcmp ? _GEN_13862 : _GEN_12364; // @[sequencer-master.scala 646:40]
  wire  _GEN_14255 = io_op_bits_active_vfcmp ? _GEN_13863 : _GEN_12365; // @[sequencer-master.scala 646:40]
  wire  _GEN_14256 = io_op_bits_active_vfcmp ? _GEN_13864 : _GEN_12366; // @[sequencer-master.scala 646:40]
  wire  _GEN_14257 = io_op_bits_active_vfcmp ? _GEN_13865 : _GEN_12367; // @[sequencer-master.scala 646:40]
  wire  _GEN_14258 = io_op_bits_active_vfcmp ? _GEN_13866 : _GEN_12368; // @[sequencer-master.scala 646:40]
  wire  _GEN_14259 = io_op_bits_active_vfcmp ? _GEN_13867 : _GEN_12369; // @[sequencer-master.scala 646:40]
  wire  _GEN_14260 = io_op_bits_active_vfcmp ? _GEN_13988 : _GEN_12370; // @[sequencer-master.scala 646:40]
  wire  _GEN_14261 = io_op_bits_active_vfcmp ? _GEN_13989 : _GEN_12371; // @[sequencer-master.scala 646:40]
  wire  _GEN_14262 = io_op_bits_active_vfcmp ? _GEN_13990 : _GEN_12372; // @[sequencer-master.scala 646:40]
  wire  _GEN_14263 = io_op_bits_active_vfcmp ? _GEN_13991 : _GEN_12373; // @[sequencer-master.scala 646:40]
  wire  _GEN_14264 = io_op_bits_active_vfcmp ? _GEN_13992 : _GEN_12374; // @[sequencer-master.scala 646:40]
  wire  _GEN_14265 = io_op_bits_active_vfcmp ? _GEN_13993 : _GEN_12375; // @[sequencer-master.scala 646:40]
  wire  _GEN_14266 = io_op_bits_active_vfcmp ? _GEN_13994 : _GEN_12376; // @[sequencer-master.scala 646:40]
  wire  _GEN_14267 = io_op_bits_active_vfcmp ? _GEN_13995 : _GEN_12377; // @[sequencer-master.scala 646:40]
  wire  _GEN_14268 = io_op_bits_active_vfcmp ? _GEN_13652 : _GEN_12378; // @[sequencer-master.scala 646:40]
  wire  _GEN_14269 = io_op_bits_active_vfcmp ? _GEN_13653 : _GEN_12379; // @[sequencer-master.scala 646:40]
  wire  _GEN_14270 = io_op_bits_active_vfcmp ? _GEN_13654 : _GEN_12380; // @[sequencer-master.scala 646:40]
  wire  _GEN_14271 = io_op_bits_active_vfcmp ? _GEN_13655 : _GEN_12381; // @[sequencer-master.scala 646:40]
  wire  _GEN_14272 = io_op_bits_active_vfcmp ? _GEN_13656 : _GEN_12382; // @[sequencer-master.scala 646:40]
  wire  _GEN_14273 = io_op_bits_active_vfcmp ? _GEN_13657 : _GEN_12383; // @[sequencer-master.scala 646:40]
  wire  _GEN_14274 = io_op_bits_active_vfcmp ? _GEN_13658 : _GEN_12384; // @[sequencer-master.scala 646:40]
  wire  _GEN_14275 = io_op_bits_active_vfcmp ? _GEN_13659 : _GEN_12385; // @[sequencer-master.scala 646:40]
  wire  _GEN_14276 = io_op_bits_active_vfcmp ? _GEN_13876 : _GEN_12386; // @[sequencer-master.scala 646:40]
  wire  _GEN_14277 = io_op_bits_active_vfcmp ? _GEN_13877 : _GEN_12387; // @[sequencer-master.scala 646:40]
  wire  _GEN_14278 = io_op_bits_active_vfcmp ? _GEN_13878 : _GEN_12388; // @[sequencer-master.scala 646:40]
  wire  _GEN_14279 = io_op_bits_active_vfcmp ? _GEN_13879 : _GEN_12389; // @[sequencer-master.scala 646:40]
  wire  _GEN_14280 = io_op_bits_active_vfcmp ? _GEN_13880 : _GEN_12390; // @[sequencer-master.scala 646:40]
  wire  _GEN_14281 = io_op_bits_active_vfcmp ? _GEN_13881 : _GEN_12391; // @[sequencer-master.scala 646:40]
  wire  _GEN_14282 = io_op_bits_active_vfcmp ? _GEN_13882 : _GEN_12392; // @[sequencer-master.scala 646:40]
  wire  _GEN_14283 = io_op_bits_active_vfcmp ? _GEN_13883 : _GEN_12393; // @[sequencer-master.scala 646:40]
  wire  _GEN_14284 = io_op_bits_active_vfcmp ? _GEN_14004 : _GEN_12394; // @[sequencer-master.scala 646:40]
  wire  _GEN_14285 = io_op_bits_active_vfcmp ? _GEN_14005 : _GEN_12395; // @[sequencer-master.scala 646:40]
  wire  _GEN_14286 = io_op_bits_active_vfcmp ? _GEN_14006 : _GEN_12396; // @[sequencer-master.scala 646:40]
  wire  _GEN_14287 = io_op_bits_active_vfcmp ? _GEN_14007 : _GEN_12397; // @[sequencer-master.scala 646:40]
  wire  _GEN_14288 = io_op_bits_active_vfcmp ? _GEN_14008 : _GEN_12398; // @[sequencer-master.scala 646:40]
  wire  _GEN_14289 = io_op_bits_active_vfcmp ? _GEN_14009 : _GEN_12399; // @[sequencer-master.scala 646:40]
  wire  _GEN_14290 = io_op_bits_active_vfcmp ? _GEN_14010 : _GEN_12400; // @[sequencer-master.scala 646:40]
  wire  _GEN_14291 = io_op_bits_active_vfcmp ? _GEN_14011 : _GEN_12401; // @[sequencer-master.scala 646:40]
  wire  _GEN_14292 = io_op_bits_active_vfcmp ? _GEN_13668 : _GEN_12402; // @[sequencer-master.scala 646:40]
  wire  _GEN_14293 = io_op_bits_active_vfcmp ? _GEN_13669 : _GEN_12403; // @[sequencer-master.scala 646:40]
  wire  _GEN_14294 = io_op_bits_active_vfcmp ? _GEN_13670 : _GEN_12404; // @[sequencer-master.scala 646:40]
  wire  _GEN_14295 = io_op_bits_active_vfcmp ? _GEN_13671 : _GEN_12405; // @[sequencer-master.scala 646:40]
  wire  _GEN_14296 = io_op_bits_active_vfcmp ? _GEN_13672 : _GEN_12406; // @[sequencer-master.scala 646:40]
  wire  _GEN_14297 = io_op_bits_active_vfcmp ? _GEN_13673 : _GEN_12407; // @[sequencer-master.scala 646:40]
  wire  _GEN_14298 = io_op_bits_active_vfcmp ? _GEN_13674 : _GEN_12408; // @[sequencer-master.scala 646:40]
  wire  _GEN_14299 = io_op_bits_active_vfcmp ? _GEN_13675 : _GEN_12409; // @[sequencer-master.scala 646:40]
  wire  _GEN_14300 = io_op_bits_active_vfcmp ? _GEN_13892 : _GEN_12410; // @[sequencer-master.scala 646:40]
  wire  _GEN_14301 = io_op_bits_active_vfcmp ? _GEN_13893 : _GEN_12411; // @[sequencer-master.scala 646:40]
  wire  _GEN_14302 = io_op_bits_active_vfcmp ? _GEN_13894 : _GEN_12412; // @[sequencer-master.scala 646:40]
  wire  _GEN_14303 = io_op_bits_active_vfcmp ? _GEN_13895 : _GEN_12413; // @[sequencer-master.scala 646:40]
  wire  _GEN_14304 = io_op_bits_active_vfcmp ? _GEN_13896 : _GEN_12414; // @[sequencer-master.scala 646:40]
  wire  _GEN_14305 = io_op_bits_active_vfcmp ? _GEN_13897 : _GEN_12415; // @[sequencer-master.scala 646:40]
  wire  _GEN_14306 = io_op_bits_active_vfcmp ? _GEN_13898 : _GEN_12416; // @[sequencer-master.scala 646:40]
  wire  _GEN_14307 = io_op_bits_active_vfcmp ? _GEN_13899 : _GEN_12417; // @[sequencer-master.scala 646:40]
  wire  _GEN_14308 = io_op_bits_active_vfcmp ? _GEN_14020 : _GEN_12418; // @[sequencer-master.scala 646:40]
  wire  _GEN_14309 = io_op_bits_active_vfcmp ? _GEN_14021 : _GEN_12419; // @[sequencer-master.scala 646:40]
  wire  _GEN_14310 = io_op_bits_active_vfcmp ? _GEN_14022 : _GEN_12420; // @[sequencer-master.scala 646:40]
  wire  _GEN_14311 = io_op_bits_active_vfcmp ? _GEN_14023 : _GEN_12421; // @[sequencer-master.scala 646:40]
  wire  _GEN_14312 = io_op_bits_active_vfcmp ? _GEN_14024 : _GEN_12422; // @[sequencer-master.scala 646:40]
  wire  _GEN_14313 = io_op_bits_active_vfcmp ? _GEN_14025 : _GEN_12423; // @[sequencer-master.scala 646:40]
  wire  _GEN_14314 = io_op_bits_active_vfcmp ? _GEN_14026 : _GEN_12424; // @[sequencer-master.scala 646:40]
  wire  _GEN_14315 = io_op_bits_active_vfcmp ? _GEN_14027 : _GEN_12425; // @[sequencer-master.scala 646:40]
  wire  _GEN_14316 = io_op_bits_active_vfcmp ? _GEN_13684 : _GEN_12426; // @[sequencer-master.scala 646:40]
  wire  _GEN_14317 = io_op_bits_active_vfcmp ? _GEN_13685 : _GEN_12427; // @[sequencer-master.scala 646:40]
  wire  _GEN_14318 = io_op_bits_active_vfcmp ? _GEN_13686 : _GEN_12428; // @[sequencer-master.scala 646:40]
  wire  _GEN_14319 = io_op_bits_active_vfcmp ? _GEN_13687 : _GEN_12429; // @[sequencer-master.scala 646:40]
  wire  _GEN_14320 = io_op_bits_active_vfcmp ? _GEN_13688 : _GEN_12430; // @[sequencer-master.scala 646:40]
  wire  _GEN_14321 = io_op_bits_active_vfcmp ? _GEN_13689 : _GEN_12431; // @[sequencer-master.scala 646:40]
  wire  _GEN_14322 = io_op_bits_active_vfcmp ? _GEN_13690 : _GEN_12432; // @[sequencer-master.scala 646:40]
  wire  _GEN_14323 = io_op_bits_active_vfcmp ? _GEN_13691 : _GEN_12433; // @[sequencer-master.scala 646:40]
  wire  _GEN_14324 = io_op_bits_active_vfcmp ? _GEN_13908 : _GEN_12434; // @[sequencer-master.scala 646:40]
  wire  _GEN_14325 = io_op_bits_active_vfcmp ? _GEN_13909 : _GEN_12435; // @[sequencer-master.scala 646:40]
  wire  _GEN_14326 = io_op_bits_active_vfcmp ? _GEN_13910 : _GEN_12436; // @[sequencer-master.scala 646:40]
  wire  _GEN_14327 = io_op_bits_active_vfcmp ? _GEN_13911 : _GEN_12437; // @[sequencer-master.scala 646:40]
  wire  _GEN_14328 = io_op_bits_active_vfcmp ? _GEN_13912 : _GEN_12438; // @[sequencer-master.scala 646:40]
  wire  _GEN_14329 = io_op_bits_active_vfcmp ? _GEN_13913 : _GEN_12439; // @[sequencer-master.scala 646:40]
  wire  _GEN_14330 = io_op_bits_active_vfcmp ? _GEN_13914 : _GEN_12440; // @[sequencer-master.scala 646:40]
  wire  _GEN_14331 = io_op_bits_active_vfcmp ? _GEN_13915 : _GEN_12441; // @[sequencer-master.scala 646:40]
  wire  _GEN_14332 = io_op_bits_active_vfcmp ? _GEN_14036 : _GEN_12442; // @[sequencer-master.scala 646:40]
  wire  _GEN_14333 = io_op_bits_active_vfcmp ? _GEN_14037 : _GEN_12443; // @[sequencer-master.scala 646:40]
  wire  _GEN_14334 = io_op_bits_active_vfcmp ? _GEN_14038 : _GEN_12444; // @[sequencer-master.scala 646:40]
  wire  _GEN_14335 = io_op_bits_active_vfcmp ? _GEN_14039 : _GEN_12445; // @[sequencer-master.scala 646:40]
  wire  _GEN_14336 = io_op_bits_active_vfcmp ? _GEN_14040 : _GEN_12446; // @[sequencer-master.scala 646:40]
  wire  _GEN_14337 = io_op_bits_active_vfcmp ? _GEN_14041 : _GEN_12447; // @[sequencer-master.scala 646:40]
  wire  _GEN_14338 = io_op_bits_active_vfcmp ? _GEN_14042 : _GEN_12448; // @[sequencer-master.scala 646:40]
  wire  _GEN_14339 = io_op_bits_active_vfcmp ? _GEN_14043 : _GEN_12449; // @[sequencer-master.scala 646:40]
  wire  _GEN_14340 = io_op_bits_active_vfcmp ? _GEN_13700 : _GEN_12450; // @[sequencer-master.scala 646:40]
  wire  _GEN_14341 = io_op_bits_active_vfcmp ? _GEN_13701 : _GEN_12451; // @[sequencer-master.scala 646:40]
  wire  _GEN_14342 = io_op_bits_active_vfcmp ? _GEN_13702 : _GEN_12452; // @[sequencer-master.scala 646:40]
  wire  _GEN_14343 = io_op_bits_active_vfcmp ? _GEN_13703 : _GEN_12453; // @[sequencer-master.scala 646:40]
  wire  _GEN_14344 = io_op_bits_active_vfcmp ? _GEN_13704 : _GEN_12454; // @[sequencer-master.scala 646:40]
  wire  _GEN_14345 = io_op_bits_active_vfcmp ? _GEN_13705 : _GEN_12455; // @[sequencer-master.scala 646:40]
  wire  _GEN_14346 = io_op_bits_active_vfcmp ? _GEN_13706 : _GEN_12456; // @[sequencer-master.scala 646:40]
  wire  _GEN_14347 = io_op_bits_active_vfcmp ? _GEN_13707 : _GEN_12457; // @[sequencer-master.scala 646:40]
  wire  _GEN_14348 = io_op_bits_active_vfcmp ? _GEN_13924 : _GEN_12458; // @[sequencer-master.scala 646:40]
  wire  _GEN_14349 = io_op_bits_active_vfcmp ? _GEN_13925 : _GEN_12459; // @[sequencer-master.scala 646:40]
  wire  _GEN_14350 = io_op_bits_active_vfcmp ? _GEN_13926 : _GEN_12460; // @[sequencer-master.scala 646:40]
  wire  _GEN_14351 = io_op_bits_active_vfcmp ? _GEN_13927 : _GEN_12461; // @[sequencer-master.scala 646:40]
  wire  _GEN_14352 = io_op_bits_active_vfcmp ? _GEN_13928 : _GEN_12462; // @[sequencer-master.scala 646:40]
  wire  _GEN_14353 = io_op_bits_active_vfcmp ? _GEN_13929 : _GEN_12463; // @[sequencer-master.scala 646:40]
  wire  _GEN_14354 = io_op_bits_active_vfcmp ? _GEN_13930 : _GEN_12464; // @[sequencer-master.scala 646:40]
  wire  _GEN_14355 = io_op_bits_active_vfcmp ? _GEN_13931 : _GEN_12465; // @[sequencer-master.scala 646:40]
  wire  _GEN_14356 = io_op_bits_active_vfcmp ? _GEN_14052 : _GEN_12466; // @[sequencer-master.scala 646:40]
  wire  _GEN_14357 = io_op_bits_active_vfcmp ? _GEN_14053 : _GEN_12467; // @[sequencer-master.scala 646:40]
  wire  _GEN_14358 = io_op_bits_active_vfcmp ? _GEN_14054 : _GEN_12468; // @[sequencer-master.scala 646:40]
  wire  _GEN_14359 = io_op_bits_active_vfcmp ? _GEN_14055 : _GEN_12469; // @[sequencer-master.scala 646:40]
  wire  _GEN_14360 = io_op_bits_active_vfcmp ? _GEN_14056 : _GEN_12470; // @[sequencer-master.scala 646:40]
  wire  _GEN_14361 = io_op_bits_active_vfcmp ? _GEN_14057 : _GEN_12471; // @[sequencer-master.scala 646:40]
  wire  _GEN_14362 = io_op_bits_active_vfcmp ? _GEN_14058 : _GEN_12472; // @[sequencer-master.scala 646:40]
  wire  _GEN_14363 = io_op_bits_active_vfcmp ? _GEN_14059 : _GEN_12473; // @[sequencer-master.scala 646:40]
  wire  _GEN_14364 = io_op_bits_active_vfcmp ? _GEN_13716 : _GEN_12474; // @[sequencer-master.scala 646:40]
  wire  _GEN_14365 = io_op_bits_active_vfcmp ? _GEN_13717 : _GEN_12475; // @[sequencer-master.scala 646:40]
  wire  _GEN_14366 = io_op_bits_active_vfcmp ? _GEN_13718 : _GEN_12476; // @[sequencer-master.scala 646:40]
  wire  _GEN_14367 = io_op_bits_active_vfcmp ? _GEN_13719 : _GEN_12477; // @[sequencer-master.scala 646:40]
  wire  _GEN_14368 = io_op_bits_active_vfcmp ? _GEN_13720 : _GEN_12478; // @[sequencer-master.scala 646:40]
  wire  _GEN_14369 = io_op_bits_active_vfcmp ? _GEN_13721 : _GEN_12479; // @[sequencer-master.scala 646:40]
  wire  _GEN_14370 = io_op_bits_active_vfcmp ? _GEN_13722 : _GEN_12480; // @[sequencer-master.scala 646:40]
  wire  _GEN_14371 = io_op_bits_active_vfcmp ? _GEN_13723 : _GEN_12481; // @[sequencer-master.scala 646:40]
  wire  _GEN_14372 = io_op_bits_active_vfcmp ? _GEN_13940 : _GEN_12482; // @[sequencer-master.scala 646:40]
  wire  _GEN_14373 = io_op_bits_active_vfcmp ? _GEN_13941 : _GEN_12483; // @[sequencer-master.scala 646:40]
  wire  _GEN_14374 = io_op_bits_active_vfcmp ? _GEN_13942 : _GEN_12484; // @[sequencer-master.scala 646:40]
  wire  _GEN_14375 = io_op_bits_active_vfcmp ? _GEN_13943 : _GEN_12485; // @[sequencer-master.scala 646:40]
  wire  _GEN_14376 = io_op_bits_active_vfcmp ? _GEN_13944 : _GEN_12486; // @[sequencer-master.scala 646:40]
  wire  _GEN_14377 = io_op_bits_active_vfcmp ? _GEN_13945 : _GEN_12487; // @[sequencer-master.scala 646:40]
  wire  _GEN_14378 = io_op_bits_active_vfcmp ? _GEN_13946 : _GEN_12488; // @[sequencer-master.scala 646:40]
  wire  _GEN_14379 = io_op_bits_active_vfcmp ? _GEN_13947 : _GEN_12489; // @[sequencer-master.scala 646:40]
  wire  _GEN_14380 = io_op_bits_active_vfcmp ? _GEN_14068 : _GEN_12490; // @[sequencer-master.scala 646:40]
  wire  _GEN_14381 = io_op_bits_active_vfcmp ? _GEN_14069 : _GEN_12491; // @[sequencer-master.scala 646:40]
  wire  _GEN_14382 = io_op_bits_active_vfcmp ? _GEN_14070 : _GEN_12492; // @[sequencer-master.scala 646:40]
  wire  _GEN_14383 = io_op_bits_active_vfcmp ? _GEN_14071 : _GEN_12493; // @[sequencer-master.scala 646:40]
  wire  _GEN_14384 = io_op_bits_active_vfcmp ? _GEN_14072 : _GEN_12494; // @[sequencer-master.scala 646:40]
  wire  _GEN_14385 = io_op_bits_active_vfcmp ? _GEN_14073 : _GEN_12495; // @[sequencer-master.scala 646:40]
  wire  _GEN_14386 = io_op_bits_active_vfcmp ? _GEN_14074 : _GEN_12496; // @[sequencer-master.scala 646:40]
  wire  _GEN_14387 = io_op_bits_active_vfcmp ? _GEN_14075 : _GEN_12497; // @[sequencer-master.scala 646:40]
  wire  _GEN_14388 = io_op_bits_active_vfcmp ? _GEN_12988 : _GEN_12498; // @[sequencer-master.scala 646:40]
  wire  _GEN_14389 = io_op_bits_active_vfcmp ? _GEN_12989 : _GEN_12499; // @[sequencer-master.scala 646:40]
  wire  _GEN_14390 = io_op_bits_active_vfcmp ? _GEN_12990 : _GEN_12500; // @[sequencer-master.scala 646:40]
  wire  _GEN_14391 = io_op_bits_active_vfcmp ? _GEN_12991 : _GEN_12501; // @[sequencer-master.scala 646:40]
  wire  _GEN_14392 = io_op_bits_active_vfcmp ? _GEN_12992 : _GEN_12502; // @[sequencer-master.scala 646:40]
  wire  _GEN_14393 = io_op_bits_active_vfcmp ? _GEN_12993 : _GEN_12503; // @[sequencer-master.scala 646:40]
  wire  _GEN_14394 = io_op_bits_active_vfcmp ? _GEN_12994 : _GEN_12504; // @[sequencer-master.scala 646:40]
  wire  _GEN_14395 = io_op_bits_active_vfcmp ? _GEN_12995 : _GEN_12505; // @[sequencer-master.scala 646:40]
  wire  _GEN_14404 = io_op_bits_active_vfcmp ? _GEN_13004 : e_0_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14405 = io_op_bits_active_vfcmp ? _GEN_13005 : e_1_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14406 = io_op_bits_active_vfcmp ? _GEN_13006 : e_2_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14407 = io_op_bits_active_vfcmp ? _GEN_13007 : e_3_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14408 = io_op_bits_active_vfcmp ? _GEN_13008 : e_4_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14409 = io_op_bits_active_vfcmp ? _GEN_13009 : e_5_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14410 = io_op_bits_active_vfcmp ? _GEN_13010 : e_6_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire  _GEN_14411 = io_op_bits_active_vfcmp ? _GEN_13011 : e_7_active_vfcu; // @[sequencer-master.scala 646:40 sequencer-master.scala 109:14]
  wire [9:0] _GEN_14412 = io_op_bits_active_vfcmp ? _GEN_13012 : _GEN_12522; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14413 = io_op_bits_active_vfcmp ? _GEN_13013 : _GEN_12523; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14414 = io_op_bits_active_vfcmp ? _GEN_13014 : _GEN_12524; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14415 = io_op_bits_active_vfcmp ? _GEN_13015 : _GEN_12525; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14416 = io_op_bits_active_vfcmp ? _GEN_13016 : _GEN_12526; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14417 = io_op_bits_active_vfcmp ? _GEN_13017 : _GEN_12527; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14418 = io_op_bits_active_vfcmp ? _GEN_13018 : _GEN_12528; // @[sequencer-master.scala 646:40]
  wire [9:0] _GEN_14419 = io_op_bits_active_vfcmp ? _GEN_13019 : _GEN_12529; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14420 = io_op_bits_active_vfcmp ? _GEN_13060 : _GEN_12530; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14421 = io_op_bits_active_vfcmp ? _GEN_13061 : _GEN_12531; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14422 = io_op_bits_active_vfcmp ? _GEN_13062 : _GEN_12532; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14423 = io_op_bits_active_vfcmp ? _GEN_13063 : _GEN_12533; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14424 = io_op_bits_active_vfcmp ? _GEN_13064 : _GEN_12534; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14425 = io_op_bits_active_vfcmp ? _GEN_13065 : _GEN_12535; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14426 = io_op_bits_active_vfcmp ? _GEN_13066 : _GEN_12536; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14427 = io_op_bits_active_vfcmp ? _GEN_13067 : _GEN_12537; // @[sequencer-master.scala 646:40]
  wire  _GEN_14428 = io_op_bits_active_vfcmp ? _GEN_13076 : _GEN_12538; // @[sequencer-master.scala 646:40]
  wire  _GEN_14429 = io_op_bits_active_vfcmp ? _GEN_13077 : _GEN_12539; // @[sequencer-master.scala 646:40]
  wire  _GEN_14430 = io_op_bits_active_vfcmp ? _GEN_13078 : _GEN_12540; // @[sequencer-master.scala 646:40]
  wire  _GEN_14431 = io_op_bits_active_vfcmp ? _GEN_13079 : _GEN_12541; // @[sequencer-master.scala 646:40]
  wire  _GEN_14432 = io_op_bits_active_vfcmp ? _GEN_13080 : _GEN_12542; // @[sequencer-master.scala 646:40]
  wire  _GEN_14433 = io_op_bits_active_vfcmp ? _GEN_13081 : _GEN_12543; // @[sequencer-master.scala 646:40]
  wire  _GEN_14434 = io_op_bits_active_vfcmp ? _GEN_13082 : _GEN_12544; // @[sequencer-master.scala 646:40]
  wire  _GEN_14435 = io_op_bits_active_vfcmp ? _GEN_13083 : _GEN_12545; // @[sequencer-master.scala 646:40]
  wire  _GEN_14436 = io_op_bits_active_vfcmp ? _GEN_13084 : _GEN_12546; // @[sequencer-master.scala 646:40]
  wire  _GEN_14437 = io_op_bits_active_vfcmp ? _GEN_13085 : _GEN_12547; // @[sequencer-master.scala 646:40]
  wire  _GEN_14438 = io_op_bits_active_vfcmp ? _GEN_13086 : _GEN_12548; // @[sequencer-master.scala 646:40]
  wire  _GEN_14439 = io_op_bits_active_vfcmp ? _GEN_13087 : _GEN_12549; // @[sequencer-master.scala 646:40]
  wire  _GEN_14440 = io_op_bits_active_vfcmp ? _GEN_13088 : _GEN_12550; // @[sequencer-master.scala 646:40]
  wire  _GEN_14441 = io_op_bits_active_vfcmp ? _GEN_13089 : _GEN_12551; // @[sequencer-master.scala 646:40]
  wire  _GEN_14442 = io_op_bits_active_vfcmp ? _GEN_13090 : _GEN_12552; // @[sequencer-master.scala 646:40]
  wire  _GEN_14443 = io_op_bits_active_vfcmp ? _GEN_13091 : _GEN_12553; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14444 = io_op_bits_active_vfcmp ? _GEN_13092 : _GEN_12554; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14445 = io_op_bits_active_vfcmp ? _GEN_13093 : _GEN_12555; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14446 = io_op_bits_active_vfcmp ? _GEN_13094 : _GEN_12556; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14447 = io_op_bits_active_vfcmp ? _GEN_13095 : _GEN_12557; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14448 = io_op_bits_active_vfcmp ? _GEN_13096 : _GEN_12558; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14449 = io_op_bits_active_vfcmp ? _GEN_13097 : _GEN_12559; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14450 = io_op_bits_active_vfcmp ? _GEN_13098 : _GEN_12560; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14451 = io_op_bits_active_vfcmp ? _GEN_13099 : _GEN_12561; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14452 = io_op_bits_active_vfcmp ? _GEN_13292 : _GEN_12562; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14453 = io_op_bits_active_vfcmp ? _GEN_13293 : _GEN_12563; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14454 = io_op_bits_active_vfcmp ? _GEN_13294 : _GEN_12564; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14455 = io_op_bits_active_vfcmp ? _GEN_13295 : _GEN_12565; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14456 = io_op_bits_active_vfcmp ? _GEN_13296 : _GEN_12566; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14457 = io_op_bits_active_vfcmp ? _GEN_13297 : _GEN_12567; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14458 = io_op_bits_active_vfcmp ? _GEN_13298 : _GEN_12568; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14459 = io_op_bits_active_vfcmp ? _GEN_13299 : _GEN_12569; // @[sequencer-master.scala 646:40]
  wire  _GEN_14460 = io_op_bits_active_vfcmp ? _GEN_13308 : _GEN_12570; // @[sequencer-master.scala 646:40]
  wire  _GEN_14461 = io_op_bits_active_vfcmp ? _GEN_13309 : _GEN_12571; // @[sequencer-master.scala 646:40]
  wire  _GEN_14462 = io_op_bits_active_vfcmp ? _GEN_13310 : _GEN_12572; // @[sequencer-master.scala 646:40]
  wire  _GEN_14463 = io_op_bits_active_vfcmp ? _GEN_13311 : _GEN_12573; // @[sequencer-master.scala 646:40]
  wire  _GEN_14464 = io_op_bits_active_vfcmp ? _GEN_13312 : _GEN_12574; // @[sequencer-master.scala 646:40]
  wire  _GEN_14465 = io_op_bits_active_vfcmp ? _GEN_13313 : _GEN_12575; // @[sequencer-master.scala 646:40]
  wire  _GEN_14466 = io_op_bits_active_vfcmp ? _GEN_13314 : _GEN_12576; // @[sequencer-master.scala 646:40]
  wire  _GEN_14467 = io_op_bits_active_vfcmp ? _GEN_13315 : _GEN_12577; // @[sequencer-master.scala 646:40]
  wire  _GEN_14468 = io_op_bits_active_vfcmp ? _GEN_13316 : _GEN_12578; // @[sequencer-master.scala 646:40]
  wire  _GEN_14469 = io_op_bits_active_vfcmp ? _GEN_13317 : _GEN_12579; // @[sequencer-master.scala 646:40]
  wire  _GEN_14470 = io_op_bits_active_vfcmp ? _GEN_13318 : _GEN_12580; // @[sequencer-master.scala 646:40]
  wire  _GEN_14471 = io_op_bits_active_vfcmp ? _GEN_13319 : _GEN_12581; // @[sequencer-master.scala 646:40]
  wire  _GEN_14472 = io_op_bits_active_vfcmp ? _GEN_13320 : _GEN_12582; // @[sequencer-master.scala 646:40]
  wire  _GEN_14473 = io_op_bits_active_vfcmp ? _GEN_13321 : _GEN_12583; // @[sequencer-master.scala 646:40]
  wire  _GEN_14474 = io_op_bits_active_vfcmp ? _GEN_13322 : _GEN_12584; // @[sequencer-master.scala 646:40]
  wire  _GEN_14475 = io_op_bits_active_vfcmp ? _GEN_13323 : _GEN_12585; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14476 = io_op_bits_active_vfcmp ? _GEN_13324 : _GEN_12586; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14477 = io_op_bits_active_vfcmp ? _GEN_13325 : _GEN_12587; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14478 = io_op_bits_active_vfcmp ? _GEN_13326 : _GEN_12588; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14479 = io_op_bits_active_vfcmp ? _GEN_13327 : _GEN_12589; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14480 = io_op_bits_active_vfcmp ? _GEN_13328 : _GEN_12590; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14481 = io_op_bits_active_vfcmp ? _GEN_13329 : _GEN_12591; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14482 = io_op_bits_active_vfcmp ? _GEN_13330 : _GEN_12592; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14483 = io_op_bits_active_vfcmp ? _GEN_13331 : _GEN_12593; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14484 = io_op_bits_active_vfcmp ? _GEN_13332 : _GEN_12594; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14485 = io_op_bits_active_vfcmp ? _GEN_13333 : _GEN_12595; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14486 = io_op_bits_active_vfcmp ? _GEN_13334 : _GEN_12596; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14487 = io_op_bits_active_vfcmp ? _GEN_13335 : _GEN_12597; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14488 = io_op_bits_active_vfcmp ? _GEN_13336 : _GEN_12598; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14489 = io_op_bits_active_vfcmp ? _GEN_13337 : _GEN_12599; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14490 = io_op_bits_active_vfcmp ? _GEN_13338 : _GEN_12600; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14491 = io_op_bits_active_vfcmp ? _GEN_13339 : _GEN_12601; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14492 = io_op_bits_active_vfcmp ? _GEN_13340 : _GEN_12602; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14493 = io_op_bits_active_vfcmp ? _GEN_13341 : _GEN_12603; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14494 = io_op_bits_active_vfcmp ? _GEN_13342 : _GEN_12604; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14495 = io_op_bits_active_vfcmp ? _GEN_13343 : _GEN_12605; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14496 = io_op_bits_active_vfcmp ? _GEN_13344 : _GEN_12606; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14497 = io_op_bits_active_vfcmp ? _GEN_13345 : _GEN_12607; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14498 = io_op_bits_active_vfcmp ? _GEN_13346 : _GEN_12608; // @[sequencer-master.scala 646:40]
  wire [63:0] _GEN_14499 = io_op_bits_active_vfcmp ? _GEN_13347 : _GEN_12609; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14532 = io_op_bits_active_vfcmp ? _GEN_13580 : _GEN_12642; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14533 = io_op_bits_active_vfcmp ? _GEN_13581 : _GEN_12643; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14534 = io_op_bits_active_vfcmp ? _GEN_13582 : _GEN_12644; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14535 = io_op_bits_active_vfcmp ? _GEN_13583 : _GEN_12645; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14536 = io_op_bits_active_vfcmp ? _GEN_13584 : _GEN_12646; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14537 = io_op_bits_active_vfcmp ? _GEN_13585 : _GEN_12647; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14538 = io_op_bits_active_vfcmp ? _GEN_13586 : _GEN_12648; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14539 = io_op_bits_active_vfcmp ? _GEN_13587 : _GEN_12649; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14548 = io_op_bits_active_vfcmp ? _GEN_13772 : _GEN_12690; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14549 = io_op_bits_active_vfcmp ? _GEN_13773 : _GEN_12691; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14550 = io_op_bits_active_vfcmp ? _GEN_13774 : _GEN_12692; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14551 = io_op_bits_active_vfcmp ? _GEN_13775 : _GEN_12693; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14552 = io_op_bits_active_vfcmp ? _GEN_13776 : _GEN_12694; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14553 = io_op_bits_active_vfcmp ? _GEN_13777 : _GEN_12695; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14554 = io_op_bits_active_vfcmp ? _GEN_13778 : _GEN_12696; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14555 = io_op_bits_active_vfcmp ? _GEN_13779 : _GEN_12697; // @[sequencer-master.scala 646:40]
  wire  _GEN_14556 = io_op_bits_active_vfcmp ? _GEN_13788 : _GEN_12698; // @[sequencer-master.scala 646:40]
  wire  _GEN_14557 = io_op_bits_active_vfcmp ? _GEN_13789 : _GEN_12699; // @[sequencer-master.scala 646:40]
  wire  _GEN_14558 = io_op_bits_active_vfcmp ? _GEN_13790 : _GEN_12700; // @[sequencer-master.scala 646:40]
  wire  _GEN_14559 = io_op_bits_active_vfcmp ? _GEN_13791 : _GEN_12701; // @[sequencer-master.scala 646:40]
  wire  _GEN_14560 = io_op_bits_active_vfcmp ? _GEN_13792 : _GEN_12702; // @[sequencer-master.scala 646:40]
  wire  _GEN_14561 = io_op_bits_active_vfcmp ? _GEN_13793 : _GEN_12703; // @[sequencer-master.scala 646:40]
  wire  _GEN_14562 = io_op_bits_active_vfcmp ? _GEN_13794 : _GEN_12704; // @[sequencer-master.scala 646:40]
  wire  _GEN_14563 = io_op_bits_active_vfcmp ? _GEN_13795 : _GEN_12705; // @[sequencer-master.scala 646:40]
  wire  _GEN_14564 = io_op_bits_active_vfcmp ? _GEN_13796 : _GEN_12706; // @[sequencer-master.scala 646:40]
  wire  _GEN_14565 = io_op_bits_active_vfcmp ? _GEN_13797 : _GEN_12707; // @[sequencer-master.scala 646:40]
  wire  _GEN_14566 = io_op_bits_active_vfcmp ? _GEN_13798 : _GEN_12708; // @[sequencer-master.scala 646:40]
  wire  _GEN_14567 = io_op_bits_active_vfcmp ? _GEN_13799 : _GEN_12709; // @[sequencer-master.scala 646:40]
  wire  _GEN_14568 = io_op_bits_active_vfcmp ? _GEN_13800 : _GEN_12710; // @[sequencer-master.scala 646:40]
  wire  _GEN_14569 = io_op_bits_active_vfcmp ? _GEN_13801 : _GEN_12711; // @[sequencer-master.scala 646:40]
  wire  _GEN_14570 = io_op_bits_active_vfcmp ? _GEN_13802 : _GEN_12712; // @[sequencer-master.scala 646:40]
  wire  _GEN_14571 = io_op_bits_active_vfcmp ? _GEN_13803 : _GEN_12713; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14572 = io_op_bits_active_vfcmp ? _GEN_13804 : _GEN_12714; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14573 = io_op_bits_active_vfcmp ? _GEN_13805 : _GEN_12715; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14574 = io_op_bits_active_vfcmp ? _GEN_13806 : _GEN_12716; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14575 = io_op_bits_active_vfcmp ? _GEN_13807 : _GEN_12717; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14576 = io_op_bits_active_vfcmp ? _GEN_13808 : _GEN_12718; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14577 = io_op_bits_active_vfcmp ? _GEN_13809 : _GEN_12719; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14578 = io_op_bits_active_vfcmp ? _GEN_13810 : _GEN_12720; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14579 = io_op_bits_active_vfcmp ? _GEN_13811 : _GEN_12721; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14580 = io_op_bits_active_vfcmp ? _GEN_13812 : _GEN_12722; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14581 = io_op_bits_active_vfcmp ? _GEN_13813 : _GEN_12723; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14582 = io_op_bits_active_vfcmp ? _GEN_13814 : _GEN_12724; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14583 = io_op_bits_active_vfcmp ? _GEN_13815 : _GEN_12725; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14584 = io_op_bits_active_vfcmp ? _GEN_13816 : _GEN_12726; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14585 = io_op_bits_active_vfcmp ? _GEN_13817 : _GEN_12727; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14586 = io_op_bits_active_vfcmp ? _GEN_13818 : _GEN_12728; // @[sequencer-master.scala 646:40]
  wire [7:0] _GEN_14587 = io_op_bits_active_vfcmp ? _GEN_13819 : _GEN_12729; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14588 = io_op_bits_active_vfcmp ? _GEN_14076 : _GEN_12658; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14589 = io_op_bits_active_vfcmp ? _GEN_14077 : _GEN_12659; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14590 = io_op_bits_active_vfcmp ? _GEN_14078 : _GEN_12660; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14591 = io_op_bits_active_vfcmp ? _GEN_14079 : _GEN_12661; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14592 = io_op_bits_active_vfcmp ? _GEN_14080 : _GEN_12662; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14593 = io_op_bits_active_vfcmp ? _GEN_14081 : _GEN_12663; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14594 = io_op_bits_active_vfcmp ? _GEN_14082 : _GEN_12664; // @[sequencer-master.scala 646:40]
  wire [1:0] _GEN_14595 = io_op_bits_active_vfcmp ? _GEN_14083 : _GEN_12665; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14596 = io_op_bits_active_vfcmp ? _GEN_14108 : _GEN_12666; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14597 = io_op_bits_active_vfcmp ? _GEN_14109 : _GEN_12667; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14598 = io_op_bits_active_vfcmp ? _GEN_14110 : _GEN_12668; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14599 = io_op_bits_active_vfcmp ? _GEN_14111 : _GEN_12669; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14600 = io_op_bits_active_vfcmp ? _GEN_14112 : _GEN_12670; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14601 = io_op_bits_active_vfcmp ? _GEN_14113 : _GEN_12671; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14602 = io_op_bits_active_vfcmp ? _GEN_14114 : _GEN_12672; // @[sequencer-master.scala 646:40]
  wire [3:0] _GEN_14603 = io_op_bits_active_vfcmp ? _GEN_14115 : _GEN_12673; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14604 = io_op_bits_active_vfcmp ? _GEN_14124 : _GEN_12674; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14605 = io_op_bits_active_vfcmp ? _GEN_14125 : _GEN_12675; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14606 = io_op_bits_active_vfcmp ? _GEN_14126 : _GEN_12676; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14607 = io_op_bits_active_vfcmp ? _GEN_14127 : _GEN_12677; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14608 = io_op_bits_active_vfcmp ? _GEN_14128 : _GEN_12678; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14609 = io_op_bits_active_vfcmp ? _GEN_14129 : _GEN_12679; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14610 = io_op_bits_active_vfcmp ? _GEN_14130 : _GEN_12680; // @[sequencer-master.scala 646:40]
  wire [2:0] _GEN_14611 = io_op_bits_active_vfcmp ? _GEN_14131 : _GEN_12681; // @[sequencer-master.scala 646:40]
  wire  _GEN_14612 = io_op_bits_active_vfcmp | _GEN_12730; // @[sequencer-master.scala 646:40 sequencer-master.scala 265:41]
  wire [2:0] _GEN_14613 = io_op_bits_active_vfcmp ? _T_1645 : _GEN_12731; // @[sequencer-master.scala 646:40 sequencer-master.scala 265:66]
  wire  _GEN_14614 = _GEN_32729 | _GEN_14132; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14615 = _GEN_32730 | _GEN_14133; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14616 = _GEN_32731 | _GEN_14134; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14617 = _GEN_32732 | _GEN_14135; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14618 = _GEN_32733 | _GEN_14136; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14619 = _GEN_32734 | _GEN_14137; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14620 = _GEN_32735 | _GEN_14138; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14621 = _GEN_32736 | _GEN_14139; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_14630 = 3'h0 == tail ? 1'h0 : _GEN_14148; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14631 = 3'h1 == tail ? 1'h0 : _GEN_14149; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14632 = 3'h2 == tail ? 1'h0 : _GEN_14150; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14633 = 3'h3 == tail ? 1'h0 : _GEN_14151; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14634 = 3'h4 == tail ? 1'h0 : _GEN_14152; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14635 = 3'h5 == tail ? 1'h0 : _GEN_14153; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14636 = 3'h6 == tail ? 1'h0 : _GEN_14154; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14637 = 3'h7 == tail ? 1'h0 : _GEN_14155; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_14638 = 3'h0 == tail ? 1'h0 : _GEN_14156; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14639 = 3'h1 == tail ? 1'h0 : _GEN_14157; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14640 = 3'h2 == tail ? 1'h0 : _GEN_14158; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14641 = 3'h3 == tail ? 1'h0 : _GEN_14159; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14642 = 3'h4 == tail ? 1'h0 : _GEN_14160; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14643 = 3'h5 == tail ? 1'h0 : _GEN_14161; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14644 = 3'h6 == tail ? 1'h0 : _GEN_14162; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14645 = 3'h7 == tail ? 1'h0 : _GEN_14163; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_14646 = 3'h0 == tail ? 1'h0 : _GEN_14164; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14647 = 3'h1 == tail ? 1'h0 : _GEN_14165; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14648 = 3'h2 == tail ? 1'h0 : _GEN_14166; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14649 = 3'h3 == tail ? 1'h0 : _GEN_14167; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14650 = 3'h4 == tail ? 1'h0 : _GEN_14168; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14651 = 3'h5 == tail ? 1'h0 : _GEN_14169; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14652 = 3'h6 == tail ? 1'h0 : _GEN_14170; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14653 = 3'h7 == tail ? 1'h0 : _GEN_14171; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_14654 = 3'h0 == tail ? 1'h0 : _GEN_14172; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14655 = 3'h1 == tail ? 1'h0 : _GEN_14173; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14656 = 3'h2 == tail ? 1'h0 : _GEN_14174; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14657 = 3'h3 == tail ? 1'h0 : _GEN_14175; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14658 = 3'h4 == tail ? 1'h0 : _GEN_14176; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14659 = 3'h5 == tail ? 1'h0 : _GEN_14177; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14660 = 3'h6 == tail ? 1'h0 : _GEN_14178; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14661 = 3'h7 == tail ? 1'h0 : _GEN_14179; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_14662 = 3'h0 == tail ? 1'h0 : _GEN_14180; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14663 = 3'h1 == tail ? 1'h0 : _GEN_14181; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14664 = 3'h2 == tail ? 1'h0 : _GEN_14182; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14665 = 3'h3 == tail ? 1'h0 : _GEN_14183; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14666 = 3'h4 == tail ? 1'h0 : _GEN_14184; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14667 = 3'h5 == tail ? 1'h0 : _GEN_14185; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14668 = 3'h6 == tail ? 1'h0 : _GEN_14186; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14669 = 3'h7 == tail ? 1'h0 : _GEN_14187; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_14670 = _GEN_32729 | _GEN_14188; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14671 = _GEN_32730 | _GEN_14189; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14672 = _GEN_32731 | _GEN_14190; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14673 = _GEN_32732 | _GEN_14191; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14674 = _GEN_32733 | _GEN_14192; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14675 = _GEN_32734 | _GEN_14193; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14676 = _GEN_32735 | _GEN_14194; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14677 = _GEN_32736 | _GEN_14195; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_14678 = 3'h0 == tail ? 1'h0 : _GEN_14196; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14679 = 3'h1 == tail ? 1'h0 : _GEN_14197; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14680 = 3'h2 == tail ? 1'h0 : _GEN_14198; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14681 = 3'h3 == tail ? 1'h0 : _GEN_14199; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14682 = 3'h4 == tail ? 1'h0 : _GEN_14200; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14683 = 3'h5 == tail ? 1'h0 : _GEN_14201; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14684 = 3'h6 == tail ? 1'h0 : _GEN_14202; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14685 = 3'h7 == tail ? 1'h0 : _GEN_14203; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14686 = 3'h0 == tail ? 1'h0 : _GEN_14204; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14687 = 3'h1 == tail ? 1'h0 : _GEN_14205; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14688 = 3'h2 == tail ? 1'h0 : _GEN_14206; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14689 = 3'h3 == tail ? 1'h0 : _GEN_14207; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14690 = 3'h4 == tail ? 1'h0 : _GEN_14208; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14691 = 3'h5 == tail ? 1'h0 : _GEN_14209; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14692 = 3'h6 == tail ? 1'h0 : _GEN_14210; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14693 = 3'h7 == tail ? 1'h0 : _GEN_14211; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14694 = 3'h0 == tail ? 1'h0 : _GEN_14212; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14695 = 3'h1 == tail ? 1'h0 : _GEN_14213; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14696 = 3'h2 == tail ? 1'h0 : _GEN_14214; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14697 = 3'h3 == tail ? 1'h0 : _GEN_14215; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14698 = 3'h4 == tail ? 1'h0 : _GEN_14216; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14699 = 3'h5 == tail ? 1'h0 : _GEN_14217; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14700 = 3'h6 == tail ? 1'h0 : _GEN_14218; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14701 = 3'h7 == tail ? 1'h0 : _GEN_14219; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14702 = 3'h0 == tail ? 1'h0 : _GEN_14220; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14703 = 3'h1 == tail ? 1'h0 : _GEN_14221; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14704 = 3'h2 == tail ? 1'h0 : _GEN_14222; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14705 = 3'h3 == tail ? 1'h0 : _GEN_14223; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14706 = 3'h4 == tail ? 1'h0 : _GEN_14224; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14707 = 3'h5 == tail ? 1'h0 : _GEN_14225; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14708 = 3'h6 == tail ? 1'h0 : _GEN_14226; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14709 = 3'h7 == tail ? 1'h0 : _GEN_14227; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14710 = 3'h0 == tail ? 1'h0 : _GEN_14228; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14711 = 3'h1 == tail ? 1'h0 : _GEN_14229; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14712 = 3'h2 == tail ? 1'h0 : _GEN_14230; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14713 = 3'h3 == tail ? 1'h0 : _GEN_14231; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14714 = 3'h4 == tail ? 1'h0 : _GEN_14232; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14715 = 3'h5 == tail ? 1'h0 : _GEN_14233; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14716 = 3'h6 == tail ? 1'h0 : _GEN_14234; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14717 = 3'h7 == tail ? 1'h0 : _GEN_14235; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14718 = 3'h0 == tail ? 1'h0 : _GEN_14236; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14719 = 3'h1 == tail ? 1'h0 : _GEN_14237; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14720 = 3'h2 == tail ? 1'h0 : _GEN_14238; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14721 = 3'h3 == tail ? 1'h0 : _GEN_14239; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14722 = 3'h4 == tail ? 1'h0 : _GEN_14240; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14723 = 3'h5 == tail ? 1'h0 : _GEN_14241; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14724 = 3'h6 == tail ? 1'h0 : _GEN_14242; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14725 = 3'h7 == tail ? 1'h0 : _GEN_14243; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14726 = 3'h0 == tail ? 1'h0 : _GEN_14244; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14727 = 3'h1 == tail ? 1'h0 : _GEN_14245; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14728 = 3'h2 == tail ? 1'h0 : _GEN_14246; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14729 = 3'h3 == tail ? 1'h0 : _GEN_14247; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14730 = 3'h4 == tail ? 1'h0 : _GEN_14248; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14731 = 3'h5 == tail ? 1'h0 : _GEN_14249; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14732 = 3'h6 == tail ? 1'h0 : _GEN_14250; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14733 = 3'h7 == tail ? 1'h0 : _GEN_14251; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14734 = 3'h0 == tail ? 1'h0 : _GEN_14252; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14735 = 3'h1 == tail ? 1'h0 : _GEN_14253; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14736 = 3'h2 == tail ? 1'h0 : _GEN_14254; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14737 = 3'h3 == tail ? 1'h0 : _GEN_14255; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14738 = 3'h4 == tail ? 1'h0 : _GEN_14256; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14739 = 3'h5 == tail ? 1'h0 : _GEN_14257; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14740 = 3'h6 == tail ? 1'h0 : _GEN_14258; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14741 = 3'h7 == tail ? 1'h0 : _GEN_14259; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14742 = 3'h0 == tail ? 1'h0 : _GEN_14260; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14743 = 3'h1 == tail ? 1'h0 : _GEN_14261; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14744 = 3'h2 == tail ? 1'h0 : _GEN_14262; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14745 = 3'h3 == tail ? 1'h0 : _GEN_14263; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14746 = 3'h4 == tail ? 1'h0 : _GEN_14264; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14747 = 3'h5 == tail ? 1'h0 : _GEN_14265; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14748 = 3'h6 == tail ? 1'h0 : _GEN_14266; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14749 = 3'h7 == tail ? 1'h0 : _GEN_14267; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14750 = 3'h0 == tail ? 1'h0 : _GEN_14268; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14751 = 3'h1 == tail ? 1'h0 : _GEN_14269; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14752 = 3'h2 == tail ? 1'h0 : _GEN_14270; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14753 = 3'h3 == tail ? 1'h0 : _GEN_14271; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14754 = 3'h4 == tail ? 1'h0 : _GEN_14272; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14755 = 3'h5 == tail ? 1'h0 : _GEN_14273; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14756 = 3'h6 == tail ? 1'h0 : _GEN_14274; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14757 = 3'h7 == tail ? 1'h0 : _GEN_14275; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14758 = 3'h0 == tail ? 1'h0 : _GEN_14276; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14759 = 3'h1 == tail ? 1'h0 : _GEN_14277; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14760 = 3'h2 == tail ? 1'h0 : _GEN_14278; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14761 = 3'h3 == tail ? 1'h0 : _GEN_14279; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14762 = 3'h4 == tail ? 1'h0 : _GEN_14280; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14763 = 3'h5 == tail ? 1'h0 : _GEN_14281; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14764 = 3'h6 == tail ? 1'h0 : _GEN_14282; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14765 = 3'h7 == tail ? 1'h0 : _GEN_14283; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14766 = 3'h0 == tail ? 1'h0 : _GEN_14284; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14767 = 3'h1 == tail ? 1'h0 : _GEN_14285; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14768 = 3'h2 == tail ? 1'h0 : _GEN_14286; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14769 = 3'h3 == tail ? 1'h0 : _GEN_14287; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14770 = 3'h4 == tail ? 1'h0 : _GEN_14288; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14771 = 3'h5 == tail ? 1'h0 : _GEN_14289; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14772 = 3'h6 == tail ? 1'h0 : _GEN_14290; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14773 = 3'h7 == tail ? 1'h0 : _GEN_14291; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14774 = 3'h0 == tail ? 1'h0 : _GEN_14292; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14775 = 3'h1 == tail ? 1'h0 : _GEN_14293; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14776 = 3'h2 == tail ? 1'h0 : _GEN_14294; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14777 = 3'h3 == tail ? 1'h0 : _GEN_14295; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14778 = 3'h4 == tail ? 1'h0 : _GEN_14296; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14779 = 3'h5 == tail ? 1'h0 : _GEN_14297; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14780 = 3'h6 == tail ? 1'h0 : _GEN_14298; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14781 = 3'h7 == tail ? 1'h0 : _GEN_14299; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14782 = 3'h0 == tail ? 1'h0 : _GEN_14300; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14783 = 3'h1 == tail ? 1'h0 : _GEN_14301; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14784 = 3'h2 == tail ? 1'h0 : _GEN_14302; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14785 = 3'h3 == tail ? 1'h0 : _GEN_14303; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14786 = 3'h4 == tail ? 1'h0 : _GEN_14304; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14787 = 3'h5 == tail ? 1'h0 : _GEN_14305; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14788 = 3'h6 == tail ? 1'h0 : _GEN_14306; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14789 = 3'h7 == tail ? 1'h0 : _GEN_14307; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14790 = 3'h0 == tail ? 1'h0 : _GEN_14308; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14791 = 3'h1 == tail ? 1'h0 : _GEN_14309; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14792 = 3'h2 == tail ? 1'h0 : _GEN_14310; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14793 = 3'h3 == tail ? 1'h0 : _GEN_14311; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14794 = 3'h4 == tail ? 1'h0 : _GEN_14312; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14795 = 3'h5 == tail ? 1'h0 : _GEN_14313; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14796 = 3'h6 == tail ? 1'h0 : _GEN_14314; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14797 = 3'h7 == tail ? 1'h0 : _GEN_14315; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14798 = 3'h0 == tail ? 1'h0 : _GEN_14316; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14799 = 3'h1 == tail ? 1'h0 : _GEN_14317; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14800 = 3'h2 == tail ? 1'h0 : _GEN_14318; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14801 = 3'h3 == tail ? 1'h0 : _GEN_14319; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14802 = 3'h4 == tail ? 1'h0 : _GEN_14320; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14803 = 3'h5 == tail ? 1'h0 : _GEN_14321; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14804 = 3'h6 == tail ? 1'h0 : _GEN_14322; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14805 = 3'h7 == tail ? 1'h0 : _GEN_14323; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14806 = 3'h0 == tail ? 1'h0 : _GEN_14324; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14807 = 3'h1 == tail ? 1'h0 : _GEN_14325; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14808 = 3'h2 == tail ? 1'h0 : _GEN_14326; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14809 = 3'h3 == tail ? 1'h0 : _GEN_14327; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14810 = 3'h4 == tail ? 1'h0 : _GEN_14328; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14811 = 3'h5 == tail ? 1'h0 : _GEN_14329; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14812 = 3'h6 == tail ? 1'h0 : _GEN_14330; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14813 = 3'h7 == tail ? 1'h0 : _GEN_14331; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14814 = 3'h0 == tail ? 1'h0 : _GEN_14332; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14815 = 3'h1 == tail ? 1'h0 : _GEN_14333; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14816 = 3'h2 == tail ? 1'h0 : _GEN_14334; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14817 = 3'h3 == tail ? 1'h0 : _GEN_14335; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14818 = 3'h4 == tail ? 1'h0 : _GEN_14336; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14819 = 3'h5 == tail ? 1'h0 : _GEN_14337; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14820 = 3'h6 == tail ? 1'h0 : _GEN_14338; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14821 = 3'h7 == tail ? 1'h0 : _GEN_14339; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14822 = 3'h0 == tail ? 1'h0 : _GEN_14340; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14823 = 3'h1 == tail ? 1'h0 : _GEN_14341; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14824 = 3'h2 == tail ? 1'h0 : _GEN_14342; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14825 = 3'h3 == tail ? 1'h0 : _GEN_14343; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14826 = 3'h4 == tail ? 1'h0 : _GEN_14344; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14827 = 3'h5 == tail ? 1'h0 : _GEN_14345; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14828 = 3'h6 == tail ? 1'h0 : _GEN_14346; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14829 = 3'h7 == tail ? 1'h0 : _GEN_14347; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14830 = 3'h0 == tail ? 1'h0 : _GEN_14348; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14831 = 3'h1 == tail ? 1'h0 : _GEN_14349; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14832 = 3'h2 == tail ? 1'h0 : _GEN_14350; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14833 = 3'h3 == tail ? 1'h0 : _GEN_14351; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14834 = 3'h4 == tail ? 1'h0 : _GEN_14352; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14835 = 3'h5 == tail ? 1'h0 : _GEN_14353; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14836 = 3'h6 == tail ? 1'h0 : _GEN_14354; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14837 = 3'h7 == tail ? 1'h0 : _GEN_14355; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14838 = 3'h0 == tail ? 1'h0 : _GEN_14356; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14839 = 3'h1 == tail ? 1'h0 : _GEN_14357; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14840 = 3'h2 == tail ? 1'h0 : _GEN_14358; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14841 = 3'h3 == tail ? 1'h0 : _GEN_14359; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14842 = 3'h4 == tail ? 1'h0 : _GEN_14360; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14843 = 3'h5 == tail ? 1'h0 : _GEN_14361; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14844 = 3'h6 == tail ? 1'h0 : _GEN_14362; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14845 = 3'h7 == tail ? 1'h0 : _GEN_14363; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14846 = 3'h0 == tail ? 1'h0 : _GEN_14364; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14847 = 3'h1 == tail ? 1'h0 : _GEN_14365; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14848 = 3'h2 == tail ? 1'h0 : _GEN_14366; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14849 = 3'h3 == tail ? 1'h0 : _GEN_14367; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14850 = 3'h4 == tail ? 1'h0 : _GEN_14368; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14851 = 3'h5 == tail ? 1'h0 : _GEN_14369; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14852 = 3'h6 == tail ? 1'h0 : _GEN_14370; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14853 = 3'h7 == tail ? 1'h0 : _GEN_14371; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_14854 = 3'h0 == tail ? 1'h0 : _GEN_14372; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14855 = 3'h1 == tail ? 1'h0 : _GEN_14373; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14856 = 3'h2 == tail ? 1'h0 : _GEN_14374; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14857 = 3'h3 == tail ? 1'h0 : _GEN_14375; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14858 = 3'h4 == tail ? 1'h0 : _GEN_14376; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14859 = 3'h5 == tail ? 1'h0 : _GEN_14377; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14860 = 3'h6 == tail ? 1'h0 : _GEN_14378; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14861 = 3'h7 == tail ? 1'h0 : _GEN_14379; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_14862 = 3'h0 == tail ? 1'h0 : _GEN_14380; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14863 = 3'h1 == tail ? 1'h0 : _GEN_14381; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14864 = 3'h2 == tail ? 1'h0 : _GEN_14382; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14865 = 3'h3 == tail ? 1'h0 : _GEN_14383; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14866 = 3'h4 == tail ? 1'h0 : _GEN_14384; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14867 = 3'h5 == tail ? 1'h0 : _GEN_14385; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14868 = 3'h6 == tail ? 1'h0 : _GEN_14386; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14869 = 3'h7 == tail ? 1'h0 : _GEN_14387; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_14870 = 3'h0 == tail ? 1'h0 : _GEN_14388; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14871 = 3'h1 == tail ? 1'h0 : _GEN_14389; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14872 = 3'h2 == tail ? 1'h0 : _GEN_14390; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14873 = 3'h3 == tail ? 1'h0 : _GEN_14391; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14874 = 3'h4 == tail ? 1'h0 : _GEN_14392; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14875 = 3'h5 == tail ? 1'h0 : _GEN_14393; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14876 = 3'h6 == tail ? 1'h0 : _GEN_14394; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14877 = 3'h7 == tail ? 1'h0 : _GEN_14395; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_14886 = _GEN_32729 | e_0_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14887 = _GEN_32730 | e_1_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14888 = _GEN_32731 | e_2_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14889 = _GEN_32732 | e_3_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14890 = _GEN_32733 | e_4_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14891 = _GEN_32734 | e_5_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14892 = _GEN_32735 | e_6_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_14893 = _GEN_32736 | e_7_active_vfvu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_14894 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_14412; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14895 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_14413; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14896 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_14414; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14897 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_14415; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14898 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_14416; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14899 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_14417; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14900 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_14418; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_14901 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_14419; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_14902 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_14420; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14903 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_14421; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14904 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_14422; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14905 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_14423; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14906 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_14424; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14907 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_14425; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14908 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_14426; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_14909 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_14427; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14910 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_14630; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14911 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_14631; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14912 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_14632; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14913 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_14633; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14914 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_14634; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14915 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_14635; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14916 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_14636; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14917 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_14637; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14918 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_14428; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14919 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_14429; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14920 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_14430; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14921 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_14431; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14922 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_14432; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14923 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_14433; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14924 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_14434; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14925 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_14435; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14926 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_14436; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14927 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_14437; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14928 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_14438; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14929 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_14439; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14930 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_14440; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14931 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_14441; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14932 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_14442; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_14933 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_14443; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_14934 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_14444; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14935 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_14445; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14936 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_14446; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14937 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_14447; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14938 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_14448; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14939 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_14449; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14940 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_14450; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_14941 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_14451; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_14942 = io_op_bits_base_vp_valid ? _GEN_14902 : _GEN_14420; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14943 = io_op_bits_base_vp_valid ? _GEN_14903 : _GEN_14421; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14944 = io_op_bits_base_vp_valid ? _GEN_14904 : _GEN_14422; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14945 = io_op_bits_base_vp_valid ? _GEN_14905 : _GEN_14423; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14946 = io_op_bits_base_vp_valid ? _GEN_14906 : _GEN_14424; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14947 = io_op_bits_base_vp_valid ? _GEN_14907 : _GEN_14425; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14948 = io_op_bits_base_vp_valid ? _GEN_14908 : _GEN_14426; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_14949 = io_op_bits_base_vp_valid ? _GEN_14909 : _GEN_14427; // @[sequencer-master.scala 320:41]
  wire  _GEN_14950 = io_op_bits_base_vp_valid ? _GEN_14910 : _GEN_14630; // @[sequencer-master.scala 320:41]
  wire  _GEN_14951 = io_op_bits_base_vp_valid ? _GEN_14911 : _GEN_14631; // @[sequencer-master.scala 320:41]
  wire  _GEN_14952 = io_op_bits_base_vp_valid ? _GEN_14912 : _GEN_14632; // @[sequencer-master.scala 320:41]
  wire  _GEN_14953 = io_op_bits_base_vp_valid ? _GEN_14913 : _GEN_14633; // @[sequencer-master.scala 320:41]
  wire  _GEN_14954 = io_op_bits_base_vp_valid ? _GEN_14914 : _GEN_14634; // @[sequencer-master.scala 320:41]
  wire  _GEN_14955 = io_op_bits_base_vp_valid ? _GEN_14915 : _GEN_14635; // @[sequencer-master.scala 320:41]
  wire  _GEN_14956 = io_op_bits_base_vp_valid ? _GEN_14916 : _GEN_14636; // @[sequencer-master.scala 320:41]
  wire  _GEN_14957 = io_op_bits_base_vp_valid ? _GEN_14917 : _GEN_14637; // @[sequencer-master.scala 320:41]
  wire  _GEN_14958 = io_op_bits_base_vp_valid ? _GEN_14918 : _GEN_14428; // @[sequencer-master.scala 320:41]
  wire  _GEN_14959 = io_op_bits_base_vp_valid ? _GEN_14919 : _GEN_14429; // @[sequencer-master.scala 320:41]
  wire  _GEN_14960 = io_op_bits_base_vp_valid ? _GEN_14920 : _GEN_14430; // @[sequencer-master.scala 320:41]
  wire  _GEN_14961 = io_op_bits_base_vp_valid ? _GEN_14921 : _GEN_14431; // @[sequencer-master.scala 320:41]
  wire  _GEN_14962 = io_op_bits_base_vp_valid ? _GEN_14922 : _GEN_14432; // @[sequencer-master.scala 320:41]
  wire  _GEN_14963 = io_op_bits_base_vp_valid ? _GEN_14923 : _GEN_14433; // @[sequencer-master.scala 320:41]
  wire  _GEN_14964 = io_op_bits_base_vp_valid ? _GEN_14924 : _GEN_14434; // @[sequencer-master.scala 320:41]
  wire  _GEN_14965 = io_op_bits_base_vp_valid ? _GEN_14925 : _GEN_14435; // @[sequencer-master.scala 320:41]
  wire  _GEN_14966 = io_op_bits_base_vp_valid ? _GEN_14926 : _GEN_14436; // @[sequencer-master.scala 320:41]
  wire  _GEN_14967 = io_op_bits_base_vp_valid ? _GEN_14927 : _GEN_14437; // @[sequencer-master.scala 320:41]
  wire  _GEN_14968 = io_op_bits_base_vp_valid ? _GEN_14928 : _GEN_14438; // @[sequencer-master.scala 320:41]
  wire  _GEN_14969 = io_op_bits_base_vp_valid ? _GEN_14929 : _GEN_14439; // @[sequencer-master.scala 320:41]
  wire  _GEN_14970 = io_op_bits_base_vp_valid ? _GEN_14930 : _GEN_14440; // @[sequencer-master.scala 320:41]
  wire  _GEN_14971 = io_op_bits_base_vp_valid ? _GEN_14931 : _GEN_14441; // @[sequencer-master.scala 320:41]
  wire  _GEN_14972 = io_op_bits_base_vp_valid ? _GEN_14932 : _GEN_14442; // @[sequencer-master.scala 320:41]
  wire  _GEN_14973 = io_op_bits_base_vp_valid ? _GEN_14933 : _GEN_14443; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14974 = io_op_bits_base_vp_valid ? _GEN_14934 : _GEN_14444; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14975 = io_op_bits_base_vp_valid ? _GEN_14935 : _GEN_14445; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14976 = io_op_bits_base_vp_valid ? _GEN_14936 : _GEN_14446; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14977 = io_op_bits_base_vp_valid ? _GEN_14937 : _GEN_14447; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14978 = io_op_bits_base_vp_valid ? _GEN_14938 : _GEN_14448; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14979 = io_op_bits_base_vp_valid ? _GEN_14939 : _GEN_14449; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14980 = io_op_bits_base_vp_valid ? _GEN_14940 : _GEN_14450; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_14981 = io_op_bits_base_vp_valid ? _GEN_14941 : _GEN_14451; // @[sequencer-master.scala 320:41]
  wire  _GEN_14982 = _GEN_32729 | _GEN_14678; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14983 = _GEN_32730 | _GEN_14679; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14984 = _GEN_32731 | _GEN_14680; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14985 = _GEN_32732 | _GEN_14681; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14986 = _GEN_32733 | _GEN_14682; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14987 = _GEN_32734 | _GEN_14683; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14988 = _GEN_32735 | _GEN_14684; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14989 = _GEN_32736 | _GEN_14685; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14990 = _T_26 ? _GEN_14982 : _GEN_14678; // @[sequencer-master.scala 154:24]
  wire  _GEN_14991 = _T_26 ? _GEN_14983 : _GEN_14679; // @[sequencer-master.scala 154:24]
  wire  _GEN_14992 = _T_26 ? _GEN_14984 : _GEN_14680; // @[sequencer-master.scala 154:24]
  wire  _GEN_14993 = _T_26 ? _GEN_14985 : _GEN_14681; // @[sequencer-master.scala 154:24]
  wire  _GEN_14994 = _T_26 ? _GEN_14986 : _GEN_14682; // @[sequencer-master.scala 154:24]
  wire  _GEN_14995 = _T_26 ? _GEN_14987 : _GEN_14683; // @[sequencer-master.scala 154:24]
  wire  _GEN_14996 = _T_26 ? _GEN_14988 : _GEN_14684; // @[sequencer-master.scala 154:24]
  wire  _GEN_14997 = _T_26 ? _GEN_14989 : _GEN_14685; // @[sequencer-master.scala 154:24]
  wire  _GEN_14998 = _GEN_32729 | _GEN_14702; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_14999 = _GEN_32730 | _GEN_14703; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15000 = _GEN_32731 | _GEN_14704; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15001 = _GEN_32732 | _GEN_14705; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15002 = _GEN_32733 | _GEN_14706; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15003 = _GEN_32734 | _GEN_14707; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15004 = _GEN_32735 | _GEN_14708; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15005 = _GEN_32736 | _GEN_14709; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15006 = _T_48 ? _GEN_14998 : _GEN_14702; // @[sequencer-master.scala 154:24]
  wire  _GEN_15007 = _T_48 ? _GEN_14999 : _GEN_14703; // @[sequencer-master.scala 154:24]
  wire  _GEN_15008 = _T_48 ? _GEN_15000 : _GEN_14704; // @[sequencer-master.scala 154:24]
  wire  _GEN_15009 = _T_48 ? _GEN_15001 : _GEN_14705; // @[sequencer-master.scala 154:24]
  wire  _GEN_15010 = _T_48 ? _GEN_15002 : _GEN_14706; // @[sequencer-master.scala 154:24]
  wire  _GEN_15011 = _T_48 ? _GEN_15003 : _GEN_14707; // @[sequencer-master.scala 154:24]
  wire  _GEN_15012 = _T_48 ? _GEN_15004 : _GEN_14708; // @[sequencer-master.scala 154:24]
  wire  _GEN_15013 = _T_48 ? _GEN_15005 : _GEN_14709; // @[sequencer-master.scala 154:24]
  wire  _GEN_15014 = _GEN_32729 | _GEN_14726; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15015 = _GEN_32730 | _GEN_14727; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15016 = _GEN_32731 | _GEN_14728; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15017 = _GEN_32732 | _GEN_14729; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15018 = _GEN_32733 | _GEN_14730; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15019 = _GEN_32734 | _GEN_14731; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15020 = _GEN_32735 | _GEN_14732; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15021 = _GEN_32736 | _GEN_14733; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15022 = _T_70 ? _GEN_15014 : _GEN_14726; // @[sequencer-master.scala 154:24]
  wire  _GEN_15023 = _T_70 ? _GEN_15015 : _GEN_14727; // @[sequencer-master.scala 154:24]
  wire  _GEN_15024 = _T_70 ? _GEN_15016 : _GEN_14728; // @[sequencer-master.scala 154:24]
  wire  _GEN_15025 = _T_70 ? _GEN_15017 : _GEN_14729; // @[sequencer-master.scala 154:24]
  wire  _GEN_15026 = _T_70 ? _GEN_15018 : _GEN_14730; // @[sequencer-master.scala 154:24]
  wire  _GEN_15027 = _T_70 ? _GEN_15019 : _GEN_14731; // @[sequencer-master.scala 154:24]
  wire  _GEN_15028 = _T_70 ? _GEN_15020 : _GEN_14732; // @[sequencer-master.scala 154:24]
  wire  _GEN_15029 = _T_70 ? _GEN_15021 : _GEN_14733; // @[sequencer-master.scala 154:24]
  wire  _GEN_15030 = _GEN_32729 | _GEN_14750; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15031 = _GEN_32730 | _GEN_14751; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15032 = _GEN_32731 | _GEN_14752; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15033 = _GEN_32732 | _GEN_14753; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15034 = _GEN_32733 | _GEN_14754; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15035 = _GEN_32734 | _GEN_14755; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15036 = _GEN_32735 | _GEN_14756; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15037 = _GEN_32736 | _GEN_14757; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15038 = _T_92 ? _GEN_15030 : _GEN_14750; // @[sequencer-master.scala 154:24]
  wire  _GEN_15039 = _T_92 ? _GEN_15031 : _GEN_14751; // @[sequencer-master.scala 154:24]
  wire  _GEN_15040 = _T_92 ? _GEN_15032 : _GEN_14752; // @[sequencer-master.scala 154:24]
  wire  _GEN_15041 = _T_92 ? _GEN_15033 : _GEN_14753; // @[sequencer-master.scala 154:24]
  wire  _GEN_15042 = _T_92 ? _GEN_15034 : _GEN_14754; // @[sequencer-master.scala 154:24]
  wire  _GEN_15043 = _T_92 ? _GEN_15035 : _GEN_14755; // @[sequencer-master.scala 154:24]
  wire  _GEN_15044 = _T_92 ? _GEN_15036 : _GEN_14756; // @[sequencer-master.scala 154:24]
  wire  _GEN_15045 = _T_92 ? _GEN_15037 : _GEN_14757; // @[sequencer-master.scala 154:24]
  wire  _GEN_15046 = _GEN_32729 | _GEN_14774; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15047 = _GEN_32730 | _GEN_14775; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15048 = _GEN_32731 | _GEN_14776; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15049 = _GEN_32732 | _GEN_14777; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15050 = _GEN_32733 | _GEN_14778; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15051 = _GEN_32734 | _GEN_14779; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15052 = _GEN_32735 | _GEN_14780; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15053 = _GEN_32736 | _GEN_14781; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15054 = _T_114 ? _GEN_15046 : _GEN_14774; // @[sequencer-master.scala 154:24]
  wire  _GEN_15055 = _T_114 ? _GEN_15047 : _GEN_14775; // @[sequencer-master.scala 154:24]
  wire  _GEN_15056 = _T_114 ? _GEN_15048 : _GEN_14776; // @[sequencer-master.scala 154:24]
  wire  _GEN_15057 = _T_114 ? _GEN_15049 : _GEN_14777; // @[sequencer-master.scala 154:24]
  wire  _GEN_15058 = _T_114 ? _GEN_15050 : _GEN_14778; // @[sequencer-master.scala 154:24]
  wire  _GEN_15059 = _T_114 ? _GEN_15051 : _GEN_14779; // @[sequencer-master.scala 154:24]
  wire  _GEN_15060 = _T_114 ? _GEN_15052 : _GEN_14780; // @[sequencer-master.scala 154:24]
  wire  _GEN_15061 = _T_114 ? _GEN_15053 : _GEN_14781; // @[sequencer-master.scala 154:24]
  wire  _GEN_15062 = _GEN_32729 | _GEN_14798; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15063 = _GEN_32730 | _GEN_14799; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15064 = _GEN_32731 | _GEN_14800; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15065 = _GEN_32732 | _GEN_14801; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15066 = _GEN_32733 | _GEN_14802; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15067 = _GEN_32734 | _GEN_14803; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15068 = _GEN_32735 | _GEN_14804; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15069 = _GEN_32736 | _GEN_14805; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15070 = _T_136 ? _GEN_15062 : _GEN_14798; // @[sequencer-master.scala 154:24]
  wire  _GEN_15071 = _T_136 ? _GEN_15063 : _GEN_14799; // @[sequencer-master.scala 154:24]
  wire  _GEN_15072 = _T_136 ? _GEN_15064 : _GEN_14800; // @[sequencer-master.scala 154:24]
  wire  _GEN_15073 = _T_136 ? _GEN_15065 : _GEN_14801; // @[sequencer-master.scala 154:24]
  wire  _GEN_15074 = _T_136 ? _GEN_15066 : _GEN_14802; // @[sequencer-master.scala 154:24]
  wire  _GEN_15075 = _T_136 ? _GEN_15067 : _GEN_14803; // @[sequencer-master.scala 154:24]
  wire  _GEN_15076 = _T_136 ? _GEN_15068 : _GEN_14804; // @[sequencer-master.scala 154:24]
  wire  _GEN_15077 = _T_136 ? _GEN_15069 : _GEN_14805; // @[sequencer-master.scala 154:24]
  wire  _GEN_15078 = _GEN_32729 | _GEN_14822; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15079 = _GEN_32730 | _GEN_14823; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15080 = _GEN_32731 | _GEN_14824; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15081 = _GEN_32732 | _GEN_14825; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15082 = _GEN_32733 | _GEN_14826; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15083 = _GEN_32734 | _GEN_14827; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15084 = _GEN_32735 | _GEN_14828; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15085 = _GEN_32736 | _GEN_14829; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15086 = _T_158 ? _GEN_15078 : _GEN_14822; // @[sequencer-master.scala 154:24]
  wire  _GEN_15087 = _T_158 ? _GEN_15079 : _GEN_14823; // @[sequencer-master.scala 154:24]
  wire  _GEN_15088 = _T_158 ? _GEN_15080 : _GEN_14824; // @[sequencer-master.scala 154:24]
  wire  _GEN_15089 = _T_158 ? _GEN_15081 : _GEN_14825; // @[sequencer-master.scala 154:24]
  wire  _GEN_15090 = _T_158 ? _GEN_15082 : _GEN_14826; // @[sequencer-master.scala 154:24]
  wire  _GEN_15091 = _T_158 ? _GEN_15083 : _GEN_14827; // @[sequencer-master.scala 154:24]
  wire  _GEN_15092 = _T_158 ? _GEN_15084 : _GEN_14828; // @[sequencer-master.scala 154:24]
  wire  _GEN_15093 = _T_158 ? _GEN_15085 : _GEN_14829; // @[sequencer-master.scala 154:24]
  wire  _GEN_15094 = _GEN_32729 | _GEN_14846; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15095 = _GEN_32730 | _GEN_14847; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15096 = _GEN_32731 | _GEN_14848; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15097 = _GEN_32732 | _GEN_14849; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15098 = _GEN_32733 | _GEN_14850; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15099 = _GEN_32734 | _GEN_14851; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15100 = _GEN_32735 | _GEN_14852; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15101 = _GEN_32736 | _GEN_14853; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15102 = _T_180 ? _GEN_15094 : _GEN_14846; // @[sequencer-master.scala 154:24]
  wire  _GEN_15103 = _T_180 ? _GEN_15095 : _GEN_14847; // @[sequencer-master.scala 154:24]
  wire  _GEN_15104 = _T_180 ? _GEN_15096 : _GEN_14848; // @[sequencer-master.scala 154:24]
  wire  _GEN_15105 = _T_180 ? _GEN_15097 : _GEN_14849; // @[sequencer-master.scala 154:24]
  wire  _GEN_15106 = _T_180 ? _GEN_15098 : _GEN_14850; // @[sequencer-master.scala 154:24]
  wire  _GEN_15107 = _T_180 ? _GEN_15099 : _GEN_14851; // @[sequencer-master.scala 154:24]
  wire  _GEN_15108 = _T_180 ? _GEN_15100 : _GEN_14852; // @[sequencer-master.scala 154:24]
  wire  _GEN_15109 = _T_180 ? _GEN_15101 : _GEN_14853; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_15110 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_14452; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15111 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_14453; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15112 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_14454; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15113 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_14455; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15114 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_14456; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15115 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_14457; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15116 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_14458; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15117 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_14459; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15118 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_14638; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15119 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_14639; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15120 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_14640; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15121 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_14641; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15122 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_14642; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15123 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_14643; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15124 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_14644; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15125 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_14645; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15126 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_14460; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15127 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_14461; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15128 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_14462; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15129 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_14463; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15130 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_14464; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15131 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_14465; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15132 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_14466; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15133 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_14467; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15134 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_14468; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15135 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_14469; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15136 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_14470; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15137 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_14471; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15138 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_14472; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15139 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_14473; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15140 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_14474; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_15141 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_14475; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15142 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_14476; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15143 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_14477; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15144 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_14478; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15145 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_14479; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15146 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_14480; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15147 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_14481; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15148 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_14482; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_15149 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_14483; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_15150 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_14484; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15151 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_14485; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15152 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_14486; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15153 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_14487; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15154 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_14488; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15155 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_14489; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15156 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_14490; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_15157 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_14491; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_15158 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_14492; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15159 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_14493; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15160 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_14494; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15161 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_14495; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15162 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_14496; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15163 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_14497; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15164 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_14498; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15165 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_14499; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_15166 = _T_189 ? _GEN_15158 : _GEN_14492; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15167 = _T_189 ? _GEN_15159 : _GEN_14493; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15168 = _T_189 ? _GEN_15160 : _GEN_14494; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15169 = _T_189 ? _GEN_15161 : _GEN_14495; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15170 = _T_189 ? _GEN_15162 : _GEN_14496; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15171 = _T_189 ? _GEN_15163 : _GEN_14497; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15172 = _T_189 ? _GEN_15164 : _GEN_14498; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_15173 = _T_189 ? _GEN_15165 : _GEN_14499; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_15174 = io_op_bits_base_vs1_valid ? _GEN_15110 : _GEN_14452; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15175 = io_op_bits_base_vs1_valid ? _GEN_15111 : _GEN_14453; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15176 = io_op_bits_base_vs1_valid ? _GEN_15112 : _GEN_14454; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15177 = io_op_bits_base_vs1_valid ? _GEN_15113 : _GEN_14455; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15178 = io_op_bits_base_vs1_valid ? _GEN_15114 : _GEN_14456; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15179 = io_op_bits_base_vs1_valid ? _GEN_15115 : _GEN_14457; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15180 = io_op_bits_base_vs1_valid ? _GEN_15116 : _GEN_14458; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15181 = io_op_bits_base_vs1_valid ? _GEN_15117 : _GEN_14459; // @[sequencer-master.scala 328:47]
  wire  _GEN_15182 = io_op_bits_base_vs1_valid ? _GEN_15118 : _GEN_14638; // @[sequencer-master.scala 328:47]
  wire  _GEN_15183 = io_op_bits_base_vs1_valid ? _GEN_15119 : _GEN_14639; // @[sequencer-master.scala 328:47]
  wire  _GEN_15184 = io_op_bits_base_vs1_valid ? _GEN_15120 : _GEN_14640; // @[sequencer-master.scala 328:47]
  wire  _GEN_15185 = io_op_bits_base_vs1_valid ? _GEN_15121 : _GEN_14641; // @[sequencer-master.scala 328:47]
  wire  _GEN_15186 = io_op_bits_base_vs1_valid ? _GEN_15122 : _GEN_14642; // @[sequencer-master.scala 328:47]
  wire  _GEN_15187 = io_op_bits_base_vs1_valid ? _GEN_15123 : _GEN_14643; // @[sequencer-master.scala 328:47]
  wire  _GEN_15188 = io_op_bits_base_vs1_valid ? _GEN_15124 : _GEN_14644; // @[sequencer-master.scala 328:47]
  wire  _GEN_15189 = io_op_bits_base_vs1_valid ? _GEN_15125 : _GEN_14645; // @[sequencer-master.scala 328:47]
  wire  _GEN_15190 = io_op_bits_base_vs1_valid ? _GEN_15126 : _GEN_14460; // @[sequencer-master.scala 328:47]
  wire  _GEN_15191 = io_op_bits_base_vs1_valid ? _GEN_15127 : _GEN_14461; // @[sequencer-master.scala 328:47]
  wire  _GEN_15192 = io_op_bits_base_vs1_valid ? _GEN_15128 : _GEN_14462; // @[sequencer-master.scala 328:47]
  wire  _GEN_15193 = io_op_bits_base_vs1_valid ? _GEN_15129 : _GEN_14463; // @[sequencer-master.scala 328:47]
  wire  _GEN_15194 = io_op_bits_base_vs1_valid ? _GEN_15130 : _GEN_14464; // @[sequencer-master.scala 328:47]
  wire  _GEN_15195 = io_op_bits_base_vs1_valid ? _GEN_15131 : _GEN_14465; // @[sequencer-master.scala 328:47]
  wire  _GEN_15196 = io_op_bits_base_vs1_valid ? _GEN_15132 : _GEN_14466; // @[sequencer-master.scala 328:47]
  wire  _GEN_15197 = io_op_bits_base_vs1_valid ? _GEN_15133 : _GEN_14467; // @[sequencer-master.scala 328:47]
  wire  _GEN_15198 = io_op_bits_base_vs1_valid ? _GEN_15134 : _GEN_14468; // @[sequencer-master.scala 328:47]
  wire  _GEN_15199 = io_op_bits_base_vs1_valid ? _GEN_15135 : _GEN_14469; // @[sequencer-master.scala 328:47]
  wire  _GEN_15200 = io_op_bits_base_vs1_valid ? _GEN_15136 : _GEN_14470; // @[sequencer-master.scala 328:47]
  wire  _GEN_15201 = io_op_bits_base_vs1_valid ? _GEN_15137 : _GEN_14471; // @[sequencer-master.scala 328:47]
  wire  _GEN_15202 = io_op_bits_base_vs1_valid ? _GEN_15138 : _GEN_14472; // @[sequencer-master.scala 328:47]
  wire  _GEN_15203 = io_op_bits_base_vs1_valid ? _GEN_15139 : _GEN_14473; // @[sequencer-master.scala 328:47]
  wire  _GEN_15204 = io_op_bits_base_vs1_valid ? _GEN_15140 : _GEN_14474; // @[sequencer-master.scala 328:47]
  wire  _GEN_15205 = io_op_bits_base_vs1_valid ? _GEN_15141 : _GEN_14475; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15206 = io_op_bits_base_vs1_valid ? _GEN_15142 : _GEN_14476; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15207 = io_op_bits_base_vs1_valid ? _GEN_15143 : _GEN_14477; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15208 = io_op_bits_base_vs1_valid ? _GEN_15144 : _GEN_14478; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15209 = io_op_bits_base_vs1_valid ? _GEN_15145 : _GEN_14479; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15210 = io_op_bits_base_vs1_valid ? _GEN_15146 : _GEN_14480; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15211 = io_op_bits_base_vs1_valid ? _GEN_15147 : _GEN_14481; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15212 = io_op_bits_base_vs1_valid ? _GEN_15148 : _GEN_14482; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_15213 = io_op_bits_base_vs1_valid ? _GEN_15149 : _GEN_14483; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15214 = io_op_bits_base_vs1_valid ? _GEN_15150 : _GEN_14484; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15215 = io_op_bits_base_vs1_valid ? _GEN_15151 : _GEN_14485; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15216 = io_op_bits_base_vs1_valid ? _GEN_15152 : _GEN_14486; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15217 = io_op_bits_base_vs1_valid ? _GEN_15153 : _GEN_14487; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15218 = io_op_bits_base_vs1_valid ? _GEN_15154 : _GEN_14488; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15219 = io_op_bits_base_vs1_valid ? _GEN_15155 : _GEN_14489; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15220 = io_op_bits_base_vs1_valid ? _GEN_15156 : _GEN_14490; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_15221 = io_op_bits_base_vs1_valid ? _GEN_15157 : _GEN_14491; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15222 = io_op_bits_base_vs1_valid ? _GEN_15166 : _GEN_14492; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15223 = io_op_bits_base_vs1_valid ? _GEN_15167 : _GEN_14493; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15224 = io_op_bits_base_vs1_valid ? _GEN_15168 : _GEN_14494; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15225 = io_op_bits_base_vs1_valid ? _GEN_15169 : _GEN_14495; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15226 = io_op_bits_base_vs1_valid ? _GEN_15170 : _GEN_14496; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15227 = io_op_bits_base_vs1_valid ? _GEN_15171 : _GEN_14497; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15228 = io_op_bits_base_vs1_valid ? _GEN_15172 : _GEN_14498; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_15229 = io_op_bits_base_vs1_valid ? _GEN_15173 : _GEN_14499; // @[sequencer-master.scala 328:47]
  wire  _GEN_15230 = _GEN_32729 | _GEN_14990; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15231 = _GEN_32730 | _GEN_14991; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15232 = _GEN_32731 | _GEN_14992; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15233 = _GEN_32732 | _GEN_14993; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15234 = _GEN_32733 | _GEN_14994; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15235 = _GEN_32734 | _GEN_14995; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15236 = _GEN_32735 | _GEN_14996; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15237 = _GEN_32736 | _GEN_14997; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15238 = _T_203 ? _GEN_15230 : _GEN_14990; // @[sequencer-master.scala 154:24]
  wire  _GEN_15239 = _T_203 ? _GEN_15231 : _GEN_14991; // @[sequencer-master.scala 154:24]
  wire  _GEN_15240 = _T_203 ? _GEN_15232 : _GEN_14992; // @[sequencer-master.scala 154:24]
  wire  _GEN_15241 = _T_203 ? _GEN_15233 : _GEN_14993; // @[sequencer-master.scala 154:24]
  wire  _GEN_15242 = _T_203 ? _GEN_15234 : _GEN_14994; // @[sequencer-master.scala 154:24]
  wire  _GEN_15243 = _T_203 ? _GEN_15235 : _GEN_14995; // @[sequencer-master.scala 154:24]
  wire  _GEN_15244 = _T_203 ? _GEN_15236 : _GEN_14996; // @[sequencer-master.scala 154:24]
  wire  _GEN_15245 = _T_203 ? _GEN_15237 : _GEN_14997; // @[sequencer-master.scala 154:24]
  wire  _GEN_15246 = _GEN_32729 | _GEN_15006; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15247 = _GEN_32730 | _GEN_15007; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15248 = _GEN_32731 | _GEN_15008; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15249 = _GEN_32732 | _GEN_15009; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15250 = _GEN_32733 | _GEN_15010; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15251 = _GEN_32734 | _GEN_15011; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15252 = _GEN_32735 | _GEN_15012; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15253 = _GEN_32736 | _GEN_15013; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15254 = _T_225 ? _GEN_15246 : _GEN_15006; // @[sequencer-master.scala 154:24]
  wire  _GEN_15255 = _T_225 ? _GEN_15247 : _GEN_15007; // @[sequencer-master.scala 154:24]
  wire  _GEN_15256 = _T_225 ? _GEN_15248 : _GEN_15008; // @[sequencer-master.scala 154:24]
  wire  _GEN_15257 = _T_225 ? _GEN_15249 : _GEN_15009; // @[sequencer-master.scala 154:24]
  wire  _GEN_15258 = _T_225 ? _GEN_15250 : _GEN_15010; // @[sequencer-master.scala 154:24]
  wire  _GEN_15259 = _T_225 ? _GEN_15251 : _GEN_15011; // @[sequencer-master.scala 154:24]
  wire  _GEN_15260 = _T_225 ? _GEN_15252 : _GEN_15012; // @[sequencer-master.scala 154:24]
  wire  _GEN_15261 = _T_225 ? _GEN_15253 : _GEN_15013; // @[sequencer-master.scala 154:24]
  wire  _GEN_15262 = _GEN_32729 | _GEN_15022; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15263 = _GEN_32730 | _GEN_15023; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15264 = _GEN_32731 | _GEN_15024; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15265 = _GEN_32732 | _GEN_15025; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15266 = _GEN_32733 | _GEN_15026; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15267 = _GEN_32734 | _GEN_15027; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15268 = _GEN_32735 | _GEN_15028; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15269 = _GEN_32736 | _GEN_15029; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15270 = _T_247 ? _GEN_15262 : _GEN_15022; // @[sequencer-master.scala 154:24]
  wire  _GEN_15271 = _T_247 ? _GEN_15263 : _GEN_15023; // @[sequencer-master.scala 154:24]
  wire  _GEN_15272 = _T_247 ? _GEN_15264 : _GEN_15024; // @[sequencer-master.scala 154:24]
  wire  _GEN_15273 = _T_247 ? _GEN_15265 : _GEN_15025; // @[sequencer-master.scala 154:24]
  wire  _GEN_15274 = _T_247 ? _GEN_15266 : _GEN_15026; // @[sequencer-master.scala 154:24]
  wire  _GEN_15275 = _T_247 ? _GEN_15267 : _GEN_15027; // @[sequencer-master.scala 154:24]
  wire  _GEN_15276 = _T_247 ? _GEN_15268 : _GEN_15028; // @[sequencer-master.scala 154:24]
  wire  _GEN_15277 = _T_247 ? _GEN_15269 : _GEN_15029; // @[sequencer-master.scala 154:24]
  wire  _GEN_15278 = _GEN_32729 | _GEN_15038; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15279 = _GEN_32730 | _GEN_15039; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15280 = _GEN_32731 | _GEN_15040; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15281 = _GEN_32732 | _GEN_15041; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15282 = _GEN_32733 | _GEN_15042; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15283 = _GEN_32734 | _GEN_15043; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15284 = _GEN_32735 | _GEN_15044; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15285 = _GEN_32736 | _GEN_15045; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15286 = _T_269 ? _GEN_15278 : _GEN_15038; // @[sequencer-master.scala 154:24]
  wire  _GEN_15287 = _T_269 ? _GEN_15279 : _GEN_15039; // @[sequencer-master.scala 154:24]
  wire  _GEN_15288 = _T_269 ? _GEN_15280 : _GEN_15040; // @[sequencer-master.scala 154:24]
  wire  _GEN_15289 = _T_269 ? _GEN_15281 : _GEN_15041; // @[sequencer-master.scala 154:24]
  wire  _GEN_15290 = _T_269 ? _GEN_15282 : _GEN_15042; // @[sequencer-master.scala 154:24]
  wire  _GEN_15291 = _T_269 ? _GEN_15283 : _GEN_15043; // @[sequencer-master.scala 154:24]
  wire  _GEN_15292 = _T_269 ? _GEN_15284 : _GEN_15044; // @[sequencer-master.scala 154:24]
  wire  _GEN_15293 = _T_269 ? _GEN_15285 : _GEN_15045; // @[sequencer-master.scala 154:24]
  wire  _GEN_15294 = _GEN_32729 | _GEN_15054; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15295 = _GEN_32730 | _GEN_15055; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15296 = _GEN_32731 | _GEN_15056; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15297 = _GEN_32732 | _GEN_15057; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15298 = _GEN_32733 | _GEN_15058; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15299 = _GEN_32734 | _GEN_15059; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15300 = _GEN_32735 | _GEN_15060; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15301 = _GEN_32736 | _GEN_15061; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15302 = _T_291 ? _GEN_15294 : _GEN_15054; // @[sequencer-master.scala 154:24]
  wire  _GEN_15303 = _T_291 ? _GEN_15295 : _GEN_15055; // @[sequencer-master.scala 154:24]
  wire  _GEN_15304 = _T_291 ? _GEN_15296 : _GEN_15056; // @[sequencer-master.scala 154:24]
  wire  _GEN_15305 = _T_291 ? _GEN_15297 : _GEN_15057; // @[sequencer-master.scala 154:24]
  wire  _GEN_15306 = _T_291 ? _GEN_15298 : _GEN_15058; // @[sequencer-master.scala 154:24]
  wire  _GEN_15307 = _T_291 ? _GEN_15299 : _GEN_15059; // @[sequencer-master.scala 154:24]
  wire  _GEN_15308 = _T_291 ? _GEN_15300 : _GEN_15060; // @[sequencer-master.scala 154:24]
  wire  _GEN_15309 = _T_291 ? _GEN_15301 : _GEN_15061; // @[sequencer-master.scala 154:24]
  wire  _GEN_15310 = _GEN_32729 | _GEN_15070; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15311 = _GEN_32730 | _GEN_15071; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15312 = _GEN_32731 | _GEN_15072; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15313 = _GEN_32732 | _GEN_15073; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15314 = _GEN_32733 | _GEN_15074; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15315 = _GEN_32734 | _GEN_15075; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15316 = _GEN_32735 | _GEN_15076; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15317 = _GEN_32736 | _GEN_15077; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15318 = _T_313 ? _GEN_15310 : _GEN_15070; // @[sequencer-master.scala 154:24]
  wire  _GEN_15319 = _T_313 ? _GEN_15311 : _GEN_15071; // @[sequencer-master.scala 154:24]
  wire  _GEN_15320 = _T_313 ? _GEN_15312 : _GEN_15072; // @[sequencer-master.scala 154:24]
  wire  _GEN_15321 = _T_313 ? _GEN_15313 : _GEN_15073; // @[sequencer-master.scala 154:24]
  wire  _GEN_15322 = _T_313 ? _GEN_15314 : _GEN_15074; // @[sequencer-master.scala 154:24]
  wire  _GEN_15323 = _T_313 ? _GEN_15315 : _GEN_15075; // @[sequencer-master.scala 154:24]
  wire  _GEN_15324 = _T_313 ? _GEN_15316 : _GEN_15076; // @[sequencer-master.scala 154:24]
  wire  _GEN_15325 = _T_313 ? _GEN_15317 : _GEN_15077; // @[sequencer-master.scala 154:24]
  wire  _GEN_15326 = _GEN_32729 | _GEN_15086; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15327 = _GEN_32730 | _GEN_15087; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15328 = _GEN_32731 | _GEN_15088; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15329 = _GEN_32732 | _GEN_15089; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15330 = _GEN_32733 | _GEN_15090; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15331 = _GEN_32734 | _GEN_15091; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15332 = _GEN_32735 | _GEN_15092; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15333 = _GEN_32736 | _GEN_15093; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15334 = _T_335 ? _GEN_15326 : _GEN_15086; // @[sequencer-master.scala 154:24]
  wire  _GEN_15335 = _T_335 ? _GEN_15327 : _GEN_15087; // @[sequencer-master.scala 154:24]
  wire  _GEN_15336 = _T_335 ? _GEN_15328 : _GEN_15088; // @[sequencer-master.scala 154:24]
  wire  _GEN_15337 = _T_335 ? _GEN_15329 : _GEN_15089; // @[sequencer-master.scala 154:24]
  wire  _GEN_15338 = _T_335 ? _GEN_15330 : _GEN_15090; // @[sequencer-master.scala 154:24]
  wire  _GEN_15339 = _T_335 ? _GEN_15331 : _GEN_15091; // @[sequencer-master.scala 154:24]
  wire  _GEN_15340 = _T_335 ? _GEN_15332 : _GEN_15092; // @[sequencer-master.scala 154:24]
  wire  _GEN_15341 = _T_335 ? _GEN_15333 : _GEN_15093; // @[sequencer-master.scala 154:24]
  wire  _GEN_15342 = _GEN_32729 | _GEN_15102; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15343 = _GEN_32730 | _GEN_15103; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15344 = _GEN_32731 | _GEN_15104; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15345 = _GEN_32732 | _GEN_15105; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15346 = _GEN_32733 | _GEN_15106; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15347 = _GEN_32734 | _GEN_15107; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15348 = _GEN_32735 | _GEN_15108; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15349 = _GEN_32736 | _GEN_15109; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_15350 = _T_357 ? _GEN_15342 : _GEN_15102; // @[sequencer-master.scala 154:24]
  wire  _GEN_15351 = _T_357 ? _GEN_15343 : _GEN_15103; // @[sequencer-master.scala 154:24]
  wire  _GEN_15352 = _T_357 ? _GEN_15344 : _GEN_15104; // @[sequencer-master.scala 154:24]
  wire  _GEN_15353 = _T_357 ? _GEN_15345 : _GEN_15105; // @[sequencer-master.scala 154:24]
  wire  _GEN_15354 = _T_357 ? _GEN_15346 : _GEN_15106; // @[sequencer-master.scala 154:24]
  wire  _GEN_15355 = _T_357 ? _GEN_15347 : _GEN_15107; // @[sequencer-master.scala 154:24]
  wire  _GEN_15356 = _T_357 ? _GEN_15348 : _GEN_15108; // @[sequencer-master.scala 154:24]
  wire  _GEN_15357 = _T_357 ? _GEN_15349 : _GEN_15109; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_15358 = 3'h0 == tail ? io_op_bits_base_vd_id : _GEN_14548; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15359 = 3'h1 == tail ? io_op_bits_base_vd_id : _GEN_14549; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15360 = 3'h2 == tail ? io_op_bits_base_vd_id : _GEN_14550; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15361 = 3'h3 == tail ? io_op_bits_base_vd_id : _GEN_14551; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15362 = 3'h4 == tail ? io_op_bits_base_vd_id : _GEN_14552; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15363 = 3'h5 == tail ? io_op_bits_base_vd_id : _GEN_14553; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15364 = 3'h6 == tail ? io_op_bits_base_vd_id : _GEN_14554; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15365 = 3'h7 == tail ? io_op_bits_base_vd_id : _GEN_14555; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15366 = 3'h0 == tail ? io_op_bits_base_vd_valid : _GEN_14662; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15367 = 3'h1 == tail ? io_op_bits_base_vd_valid : _GEN_14663; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15368 = 3'h2 == tail ? io_op_bits_base_vd_valid : _GEN_14664; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15369 = 3'h3 == tail ? io_op_bits_base_vd_valid : _GEN_14665; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15370 = 3'h4 == tail ? io_op_bits_base_vd_valid : _GEN_14666; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15371 = 3'h5 == tail ? io_op_bits_base_vd_valid : _GEN_14667; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15372 = 3'h6 == tail ? io_op_bits_base_vd_valid : _GEN_14668; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15373 = 3'h7 == tail ? io_op_bits_base_vd_valid : _GEN_14669; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15374 = 3'h0 == tail ? io_op_bits_base_vd_scalar : _GEN_14556; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15375 = 3'h1 == tail ? io_op_bits_base_vd_scalar : _GEN_14557; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15376 = 3'h2 == tail ? io_op_bits_base_vd_scalar : _GEN_14558; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15377 = 3'h3 == tail ? io_op_bits_base_vd_scalar : _GEN_14559; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15378 = 3'h4 == tail ? io_op_bits_base_vd_scalar : _GEN_14560; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15379 = 3'h5 == tail ? io_op_bits_base_vd_scalar : _GEN_14561; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15380 = 3'h6 == tail ? io_op_bits_base_vd_scalar : _GEN_14562; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15381 = 3'h7 == tail ? io_op_bits_base_vd_scalar : _GEN_14563; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15382 = 3'h0 == tail ? io_op_bits_base_vd_pred : _GEN_14564; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15383 = 3'h1 == tail ? io_op_bits_base_vd_pred : _GEN_14565; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15384 = 3'h2 == tail ? io_op_bits_base_vd_pred : _GEN_14566; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15385 = 3'h3 == tail ? io_op_bits_base_vd_pred : _GEN_14567; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15386 = 3'h4 == tail ? io_op_bits_base_vd_pred : _GEN_14568; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15387 = 3'h5 == tail ? io_op_bits_base_vd_pred : _GEN_14569; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15388 = 3'h6 == tail ? io_op_bits_base_vd_pred : _GEN_14570; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_15389 = 3'h7 == tail ? io_op_bits_base_vd_pred : _GEN_14571; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15390 = 3'h0 == tail ? io_op_bits_base_vd_prec : _GEN_14572; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15391 = 3'h1 == tail ? io_op_bits_base_vd_prec : _GEN_14573; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15392 = 3'h2 == tail ? io_op_bits_base_vd_prec : _GEN_14574; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15393 = 3'h3 == tail ? io_op_bits_base_vd_prec : _GEN_14575; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15394 = 3'h4 == tail ? io_op_bits_base_vd_prec : _GEN_14576; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15395 = 3'h5 == tail ? io_op_bits_base_vd_prec : _GEN_14577; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15396 = 3'h6 == tail ? io_op_bits_base_vd_prec : _GEN_14578; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_15397 = 3'h7 == tail ? io_op_bits_base_vd_prec : _GEN_14579; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_15398 = 3'h0 == tail ? io_op_bits_reg_vd_id : _GEN_14580; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15399 = 3'h1 == tail ? io_op_bits_reg_vd_id : _GEN_14581; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15400 = 3'h2 == tail ? io_op_bits_reg_vd_id : _GEN_14582; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15401 = 3'h3 == tail ? io_op_bits_reg_vd_id : _GEN_14583; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15402 = 3'h4 == tail ? io_op_bits_reg_vd_id : _GEN_14584; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15403 = 3'h5 == tail ? io_op_bits_reg_vd_id : _GEN_14585; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15404 = 3'h6 == tail ? io_op_bits_reg_vd_id : _GEN_14586; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15405 = 3'h7 == tail ? io_op_bits_reg_vd_id : _GEN_14587; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_15406 = io_op_bits_base_vd_valid ? _GEN_15358 : _GEN_14548; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15407 = io_op_bits_base_vd_valid ? _GEN_15359 : _GEN_14549; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15408 = io_op_bits_base_vd_valid ? _GEN_15360 : _GEN_14550; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15409 = io_op_bits_base_vd_valid ? _GEN_15361 : _GEN_14551; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15410 = io_op_bits_base_vd_valid ? _GEN_15362 : _GEN_14552; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15411 = io_op_bits_base_vd_valid ? _GEN_15363 : _GEN_14553; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15412 = io_op_bits_base_vd_valid ? _GEN_15364 : _GEN_14554; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15413 = io_op_bits_base_vd_valid ? _GEN_15365 : _GEN_14555; // @[sequencer-master.scala 362:41]
  wire  _GEN_15414 = io_op_bits_base_vd_valid ? _GEN_15366 : _GEN_14662; // @[sequencer-master.scala 362:41]
  wire  _GEN_15415 = io_op_bits_base_vd_valid ? _GEN_15367 : _GEN_14663; // @[sequencer-master.scala 362:41]
  wire  _GEN_15416 = io_op_bits_base_vd_valid ? _GEN_15368 : _GEN_14664; // @[sequencer-master.scala 362:41]
  wire  _GEN_15417 = io_op_bits_base_vd_valid ? _GEN_15369 : _GEN_14665; // @[sequencer-master.scala 362:41]
  wire  _GEN_15418 = io_op_bits_base_vd_valid ? _GEN_15370 : _GEN_14666; // @[sequencer-master.scala 362:41]
  wire  _GEN_15419 = io_op_bits_base_vd_valid ? _GEN_15371 : _GEN_14667; // @[sequencer-master.scala 362:41]
  wire  _GEN_15420 = io_op_bits_base_vd_valid ? _GEN_15372 : _GEN_14668; // @[sequencer-master.scala 362:41]
  wire  _GEN_15421 = io_op_bits_base_vd_valid ? _GEN_15373 : _GEN_14669; // @[sequencer-master.scala 362:41]
  wire  _GEN_15422 = io_op_bits_base_vd_valid ? _GEN_15374 : _GEN_14556; // @[sequencer-master.scala 362:41]
  wire  _GEN_15423 = io_op_bits_base_vd_valid ? _GEN_15375 : _GEN_14557; // @[sequencer-master.scala 362:41]
  wire  _GEN_15424 = io_op_bits_base_vd_valid ? _GEN_15376 : _GEN_14558; // @[sequencer-master.scala 362:41]
  wire  _GEN_15425 = io_op_bits_base_vd_valid ? _GEN_15377 : _GEN_14559; // @[sequencer-master.scala 362:41]
  wire  _GEN_15426 = io_op_bits_base_vd_valid ? _GEN_15378 : _GEN_14560; // @[sequencer-master.scala 362:41]
  wire  _GEN_15427 = io_op_bits_base_vd_valid ? _GEN_15379 : _GEN_14561; // @[sequencer-master.scala 362:41]
  wire  _GEN_15428 = io_op_bits_base_vd_valid ? _GEN_15380 : _GEN_14562; // @[sequencer-master.scala 362:41]
  wire  _GEN_15429 = io_op_bits_base_vd_valid ? _GEN_15381 : _GEN_14563; // @[sequencer-master.scala 362:41]
  wire  _GEN_15430 = io_op_bits_base_vd_valid ? _GEN_15382 : _GEN_14564; // @[sequencer-master.scala 362:41]
  wire  _GEN_15431 = io_op_bits_base_vd_valid ? _GEN_15383 : _GEN_14565; // @[sequencer-master.scala 362:41]
  wire  _GEN_15432 = io_op_bits_base_vd_valid ? _GEN_15384 : _GEN_14566; // @[sequencer-master.scala 362:41]
  wire  _GEN_15433 = io_op_bits_base_vd_valid ? _GEN_15385 : _GEN_14567; // @[sequencer-master.scala 362:41]
  wire  _GEN_15434 = io_op_bits_base_vd_valid ? _GEN_15386 : _GEN_14568; // @[sequencer-master.scala 362:41]
  wire  _GEN_15435 = io_op_bits_base_vd_valid ? _GEN_15387 : _GEN_14569; // @[sequencer-master.scala 362:41]
  wire  _GEN_15436 = io_op_bits_base_vd_valid ? _GEN_15388 : _GEN_14570; // @[sequencer-master.scala 362:41]
  wire  _GEN_15437 = io_op_bits_base_vd_valid ? _GEN_15389 : _GEN_14571; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15438 = io_op_bits_base_vd_valid ? _GEN_15390 : _GEN_14572; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15439 = io_op_bits_base_vd_valid ? _GEN_15391 : _GEN_14573; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15440 = io_op_bits_base_vd_valid ? _GEN_15392 : _GEN_14574; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15441 = io_op_bits_base_vd_valid ? _GEN_15393 : _GEN_14575; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15442 = io_op_bits_base_vd_valid ? _GEN_15394 : _GEN_14576; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15443 = io_op_bits_base_vd_valid ? _GEN_15395 : _GEN_14577; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15444 = io_op_bits_base_vd_valid ? _GEN_15396 : _GEN_14578; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_15445 = io_op_bits_base_vd_valid ? _GEN_15397 : _GEN_14579; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15446 = io_op_bits_base_vd_valid ? _GEN_15398 : _GEN_14580; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15447 = io_op_bits_base_vd_valid ? _GEN_15399 : _GEN_14581; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15448 = io_op_bits_base_vd_valid ? _GEN_15400 : _GEN_14582; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15449 = io_op_bits_base_vd_valid ? _GEN_15401 : _GEN_14583; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15450 = io_op_bits_base_vd_valid ? _GEN_15402 : _GEN_14584; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15451 = io_op_bits_base_vd_valid ? _GEN_15403 : _GEN_14585; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15452 = io_op_bits_base_vd_valid ? _GEN_15404 : _GEN_14586; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_15453 = io_op_bits_base_vd_valid ? _GEN_15405 : _GEN_14587; // @[sequencer-master.scala 362:41]
  wire  _GEN_15454 = _GEN_32729 | _GEN_14686; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15455 = _GEN_32730 | _GEN_14687; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15456 = _GEN_32731 | _GEN_14688; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15457 = _GEN_32732 | _GEN_14689; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15458 = _GEN_32733 | _GEN_14690; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15459 = _GEN_32734 | _GEN_14691; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15460 = _GEN_32735 | _GEN_14692; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15461 = _GEN_32736 | _GEN_14693; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15462 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15454 : _GEN_14686; // @[sequencer-master.scala 161:86]
  wire  _GEN_15463 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15455 : _GEN_14687; // @[sequencer-master.scala 161:86]
  wire  _GEN_15464 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15456 : _GEN_14688; // @[sequencer-master.scala 161:86]
  wire  _GEN_15465 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15457 : _GEN_14689; // @[sequencer-master.scala 161:86]
  wire  _GEN_15466 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15458 : _GEN_14690; // @[sequencer-master.scala 161:86]
  wire  _GEN_15467 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15459 : _GEN_14691; // @[sequencer-master.scala 161:86]
  wire  _GEN_15468 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15460 : _GEN_14692; // @[sequencer-master.scala 161:86]
  wire  _GEN_15469 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_15461 : _GEN_14693; // @[sequencer-master.scala 161:86]
  wire  _GEN_15470 = _GEN_32729 | _GEN_14710; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15471 = _GEN_32730 | _GEN_14711; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15472 = _GEN_32731 | _GEN_14712; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15473 = _GEN_32732 | _GEN_14713; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15474 = _GEN_32733 | _GEN_14714; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15475 = _GEN_32734 | _GEN_14715; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15476 = _GEN_32735 | _GEN_14716; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15477 = _GEN_32736 | _GEN_14717; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15478 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15470 : _GEN_14710; // @[sequencer-master.scala 161:86]
  wire  _GEN_15479 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15471 : _GEN_14711; // @[sequencer-master.scala 161:86]
  wire  _GEN_15480 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15472 : _GEN_14712; // @[sequencer-master.scala 161:86]
  wire  _GEN_15481 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15473 : _GEN_14713; // @[sequencer-master.scala 161:86]
  wire  _GEN_15482 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15474 : _GEN_14714; // @[sequencer-master.scala 161:86]
  wire  _GEN_15483 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15475 : _GEN_14715; // @[sequencer-master.scala 161:86]
  wire  _GEN_15484 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15476 : _GEN_14716; // @[sequencer-master.scala 161:86]
  wire  _GEN_15485 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_15477 : _GEN_14717; // @[sequencer-master.scala 161:86]
  wire  _GEN_15486 = _GEN_32729 | _GEN_14734; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15487 = _GEN_32730 | _GEN_14735; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15488 = _GEN_32731 | _GEN_14736; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15489 = _GEN_32732 | _GEN_14737; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15490 = _GEN_32733 | _GEN_14738; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15491 = _GEN_32734 | _GEN_14739; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15492 = _GEN_32735 | _GEN_14740; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15493 = _GEN_32736 | _GEN_14741; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15494 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15486 : _GEN_14734; // @[sequencer-master.scala 161:86]
  wire  _GEN_15495 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15487 : _GEN_14735; // @[sequencer-master.scala 161:86]
  wire  _GEN_15496 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15488 : _GEN_14736; // @[sequencer-master.scala 161:86]
  wire  _GEN_15497 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15489 : _GEN_14737; // @[sequencer-master.scala 161:86]
  wire  _GEN_15498 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15490 : _GEN_14738; // @[sequencer-master.scala 161:86]
  wire  _GEN_15499 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15491 : _GEN_14739; // @[sequencer-master.scala 161:86]
  wire  _GEN_15500 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15492 : _GEN_14740; // @[sequencer-master.scala 161:86]
  wire  _GEN_15501 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_15493 : _GEN_14741; // @[sequencer-master.scala 161:86]
  wire  _GEN_15502 = _GEN_32729 | _GEN_14758; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15503 = _GEN_32730 | _GEN_14759; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15504 = _GEN_32731 | _GEN_14760; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15505 = _GEN_32732 | _GEN_14761; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15506 = _GEN_32733 | _GEN_14762; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15507 = _GEN_32734 | _GEN_14763; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15508 = _GEN_32735 | _GEN_14764; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15509 = _GEN_32736 | _GEN_14765; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15510 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15502 : _GEN_14758; // @[sequencer-master.scala 161:86]
  wire  _GEN_15511 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15503 : _GEN_14759; // @[sequencer-master.scala 161:86]
  wire  _GEN_15512 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15504 : _GEN_14760; // @[sequencer-master.scala 161:86]
  wire  _GEN_15513 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15505 : _GEN_14761; // @[sequencer-master.scala 161:86]
  wire  _GEN_15514 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15506 : _GEN_14762; // @[sequencer-master.scala 161:86]
  wire  _GEN_15515 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15507 : _GEN_14763; // @[sequencer-master.scala 161:86]
  wire  _GEN_15516 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15508 : _GEN_14764; // @[sequencer-master.scala 161:86]
  wire  _GEN_15517 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_15509 : _GEN_14765; // @[sequencer-master.scala 161:86]
  wire  _GEN_15518 = _GEN_32729 | _GEN_14782; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15519 = _GEN_32730 | _GEN_14783; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15520 = _GEN_32731 | _GEN_14784; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15521 = _GEN_32732 | _GEN_14785; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15522 = _GEN_32733 | _GEN_14786; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15523 = _GEN_32734 | _GEN_14787; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15524 = _GEN_32735 | _GEN_14788; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15525 = _GEN_32736 | _GEN_14789; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15526 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15518 : _GEN_14782; // @[sequencer-master.scala 161:86]
  wire  _GEN_15527 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15519 : _GEN_14783; // @[sequencer-master.scala 161:86]
  wire  _GEN_15528 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15520 : _GEN_14784; // @[sequencer-master.scala 161:86]
  wire  _GEN_15529 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15521 : _GEN_14785; // @[sequencer-master.scala 161:86]
  wire  _GEN_15530 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15522 : _GEN_14786; // @[sequencer-master.scala 161:86]
  wire  _GEN_15531 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15523 : _GEN_14787; // @[sequencer-master.scala 161:86]
  wire  _GEN_15532 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15524 : _GEN_14788; // @[sequencer-master.scala 161:86]
  wire  _GEN_15533 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_15525 : _GEN_14789; // @[sequencer-master.scala 161:86]
  wire  _GEN_15534 = _GEN_32729 | _GEN_14806; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15535 = _GEN_32730 | _GEN_14807; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15536 = _GEN_32731 | _GEN_14808; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15537 = _GEN_32732 | _GEN_14809; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15538 = _GEN_32733 | _GEN_14810; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15539 = _GEN_32734 | _GEN_14811; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15540 = _GEN_32735 | _GEN_14812; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15541 = _GEN_32736 | _GEN_14813; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15542 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15534 : _GEN_14806; // @[sequencer-master.scala 161:86]
  wire  _GEN_15543 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15535 : _GEN_14807; // @[sequencer-master.scala 161:86]
  wire  _GEN_15544 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15536 : _GEN_14808; // @[sequencer-master.scala 161:86]
  wire  _GEN_15545 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15537 : _GEN_14809; // @[sequencer-master.scala 161:86]
  wire  _GEN_15546 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15538 : _GEN_14810; // @[sequencer-master.scala 161:86]
  wire  _GEN_15547 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15539 : _GEN_14811; // @[sequencer-master.scala 161:86]
  wire  _GEN_15548 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15540 : _GEN_14812; // @[sequencer-master.scala 161:86]
  wire  _GEN_15549 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_15541 : _GEN_14813; // @[sequencer-master.scala 161:86]
  wire  _GEN_15550 = _GEN_32729 | _GEN_14830; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15551 = _GEN_32730 | _GEN_14831; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15552 = _GEN_32731 | _GEN_14832; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15553 = _GEN_32732 | _GEN_14833; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15554 = _GEN_32733 | _GEN_14834; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15555 = _GEN_32734 | _GEN_14835; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15556 = _GEN_32735 | _GEN_14836; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15557 = _GEN_32736 | _GEN_14837; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15558 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15550 : _GEN_14830; // @[sequencer-master.scala 161:86]
  wire  _GEN_15559 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15551 : _GEN_14831; // @[sequencer-master.scala 161:86]
  wire  _GEN_15560 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15552 : _GEN_14832; // @[sequencer-master.scala 161:86]
  wire  _GEN_15561 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15553 : _GEN_14833; // @[sequencer-master.scala 161:86]
  wire  _GEN_15562 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15554 : _GEN_14834; // @[sequencer-master.scala 161:86]
  wire  _GEN_15563 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15555 : _GEN_14835; // @[sequencer-master.scala 161:86]
  wire  _GEN_15564 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15556 : _GEN_14836; // @[sequencer-master.scala 161:86]
  wire  _GEN_15565 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_15557 : _GEN_14837; // @[sequencer-master.scala 161:86]
  wire  _GEN_15566 = _GEN_32729 | _GEN_14854; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15567 = _GEN_32730 | _GEN_14855; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15568 = _GEN_32731 | _GEN_14856; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15569 = _GEN_32732 | _GEN_14857; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15570 = _GEN_32733 | _GEN_14858; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15571 = _GEN_32734 | _GEN_14859; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15572 = _GEN_32735 | _GEN_14860; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15573 = _GEN_32736 | _GEN_14861; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_15574 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15566 : _GEN_14854; // @[sequencer-master.scala 161:86]
  wire  _GEN_15575 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15567 : _GEN_14855; // @[sequencer-master.scala 161:86]
  wire  _GEN_15576 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15568 : _GEN_14856; // @[sequencer-master.scala 161:86]
  wire  _GEN_15577 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15569 : _GEN_14857; // @[sequencer-master.scala 161:86]
  wire  _GEN_15578 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15570 : _GEN_14858; // @[sequencer-master.scala 161:86]
  wire  _GEN_15579 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15571 : _GEN_14859; // @[sequencer-master.scala 161:86]
  wire  _GEN_15580 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15572 : _GEN_14860; // @[sequencer-master.scala 161:86]
  wire  _GEN_15581 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_15573 : _GEN_14861; // @[sequencer-master.scala 161:86]
  wire  _GEN_15582 = _GEN_32729 | _GEN_14694; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15583 = _GEN_32730 | _GEN_14695; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15584 = _GEN_32731 | _GEN_14696; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15585 = _GEN_32732 | _GEN_14697; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15586 = _GEN_32733 | _GEN_14698; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15587 = _GEN_32734 | _GEN_14699; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15588 = _GEN_32735 | _GEN_14700; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15589 = _GEN_32736 | _GEN_14701; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15590 = _T_1442 ? _GEN_15582 : _GEN_14694; // @[sequencer-master.scala 168:32]
  wire  _GEN_15591 = _T_1442 ? _GEN_15583 : _GEN_14695; // @[sequencer-master.scala 168:32]
  wire  _GEN_15592 = _T_1442 ? _GEN_15584 : _GEN_14696; // @[sequencer-master.scala 168:32]
  wire  _GEN_15593 = _T_1442 ? _GEN_15585 : _GEN_14697; // @[sequencer-master.scala 168:32]
  wire  _GEN_15594 = _T_1442 ? _GEN_15586 : _GEN_14698; // @[sequencer-master.scala 168:32]
  wire  _GEN_15595 = _T_1442 ? _GEN_15587 : _GEN_14699; // @[sequencer-master.scala 168:32]
  wire  _GEN_15596 = _T_1442 ? _GEN_15588 : _GEN_14700; // @[sequencer-master.scala 168:32]
  wire  _GEN_15597 = _T_1442 ? _GEN_15589 : _GEN_14701; // @[sequencer-master.scala 168:32]
  wire  _GEN_15598 = _GEN_32729 | _GEN_14718; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15599 = _GEN_32730 | _GEN_14719; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15600 = _GEN_32731 | _GEN_14720; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15601 = _GEN_32732 | _GEN_14721; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15602 = _GEN_32733 | _GEN_14722; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15603 = _GEN_32734 | _GEN_14723; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15604 = _GEN_32735 | _GEN_14724; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15605 = _GEN_32736 | _GEN_14725; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15606 = _T_1464 ? _GEN_15598 : _GEN_14718; // @[sequencer-master.scala 168:32]
  wire  _GEN_15607 = _T_1464 ? _GEN_15599 : _GEN_14719; // @[sequencer-master.scala 168:32]
  wire  _GEN_15608 = _T_1464 ? _GEN_15600 : _GEN_14720; // @[sequencer-master.scala 168:32]
  wire  _GEN_15609 = _T_1464 ? _GEN_15601 : _GEN_14721; // @[sequencer-master.scala 168:32]
  wire  _GEN_15610 = _T_1464 ? _GEN_15602 : _GEN_14722; // @[sequencer-master.scala 168:32]
  wire  _GEN_15611 = _T_1464 ? _GEN_15603 : _GEN_14723; // @[sequencer-master.scala 168:32]
  wire  _GEN_15612 = _T_1464 ? _GEN_15604 : _GEN_14724; // @[sequencer-master.scala 168:32]
  wire  _GEN_15613 = _T_1464 ? _GEN_15605 : _GEN_14725; // @[sequencer-master.scala 168:32]
  wire  _GEN_15614 = _GEN_32729 | _GEN_14742; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15615 = _GEN_32730 | _GEN_14743; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15616 = _GEN_32731 | _GEN_14744; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15617 = _GEN_32732 | _GEN_14745; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15618 = _GEN_32733 | _GEN_14746; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15619 = _GEN_32734 | _GEN_14747; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15620 = _GEN_32735 | _GEN_14748; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15621 = _GEN_32736 | _GEN_14749; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15622 = _T_1486 ? _GEN_15614 : _GEN_14742; // @[sequencer-master.scala 168:32]
  wire  _GEN_15623 = _T_1486 ? _GEN_15615 : _GEN_14743; // @[sequencer-master.scala 168:32]
  wire  _GEN_15624 = _T_1486 ? _GEN_15616 : _GEN_14744; // @[sequencer-master.scala 168:32]
  wire  _GEN_15625 = _T_1486 ? _GEN_15617 : _GEN_14745; // @[sequencer-master.scala 168:32]
  wire  _GEN_15626 = _T_1486 ? _GEN_15618 : _GEN_14746; // @[sequencer-master.scala 168:32]
  wire  _GEN_15627 = _T_1486 ? _GEN_15619 : _GEN_14747; // @[sequencer-master.scala 168:32]
  wire  _GEN_15628 = _T_1486 ? _GEN_15620 : _GEN_14748; // @[sequencer-master.scala 168:32]
  wire  _GEN_15629 = _T_1486 ? _GEN_15621 : _GEN_14749; // @[sequencer-master.scala 168:32]
  wire  _GEN_15630 = _GEN_32729 | _GEN_14766; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15631 = _GEN_32730 | _GEN_14767; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15632 = _GEN_32731 | _GEN_14768; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15633 = _GEN_32732 | _GEN_14769; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15634 = _GEN_32733 | _GEN_14770; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15635 = _GEN_32734 | _GEN_14771; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15636 = _GEN_32735 | _GEN_14772; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15637 = _GEN_32736 | _GEN_14773; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15638 = _T_1508 ? _GEN_15630 : _GEN_14766; // @[sequencer-master.scala 168:32]
  wire  _GEN_15639 = _T_1508 ? _GEN_15631 : _GEN_14767; // @[sequencer-master.scala 168:32]
  wire  _GEN_15640 = _T_1508 ? _GEN_15632 : _GEN_14768; // @[sequencer-master.scala 168:32]
  wire  _GEN_15641 = _T_1508 ? _GEN_15633 : _GEN_14769; // @[sequencer-master.scala 168:32]
  wire  _GEN_15642 = _T_1508 ? _GEN_15634 : _GEN_14770; // @[sequencer-master.scala 168:32]
  wire  _GEN_15643 = _T_1508 ? _GEN_15635 : _GEN_14771; // @[sequencer-master.scala 168:32]
  wire  _GEN_15644 = _T_1508 ? _GEN_15636 : _GEN_14772; // @[sequencer-master.scala 168:32]
  wire  _GEN_15645 = _T_1508 ? _GEN_15637 : _GEN_14773; // @[sequencer-master.scala 168:32]
  wire  _GEN_15646 = _GEN_32729 | _GEN_14790; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15647 = _GEN_32730 | _GEN_14791; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15648 = _GEN_32731 | _GEN_14792; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15649 = _GEN_32732 | _GEN_14793; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15650 = _GEN_32733 | _GEN_14794; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15651 = _GEN_32734 | _GEN_14795; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15652 = _GEN_32735 | _GEN_14796; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15653 = _GEN_32736 | _GEN_14797; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15654 = _T_1530 ? _GEN_15646 : _GEN_14790; // @[sequencer-master.scala 168:32]
  wire  _GEN_15655 = _T_1530 ? _GEN_15647 : _GEN_14791; // @[sequencer-master.scala 168:32]
  wire  _GEN_15656 = _T_1530 ? _GEN_15648 : _GEN_14792; // @[sequencer-master.scala 168:32]
  wire  _GEN_15657 = _T_1530 ? _GEN_15649 : _GEN_14793; // @[sequencer-master.scala 168:32]
  wire  _GEN_15658 = _T_1530 ? _GEN_15650 : _GEN_14794; // @[sequencer-master.scala 168:32]
  wire  _GEN_15659 = _T_1530 ? _GEN_15651 : _GEN_14795; // @[sequencer-master.scala 168:32]
  wire  _GEN_15660 = _T_1530 ? _GEN_15652 : _GEN_14796; // @[sequencer-master.scala 168:32]
  wire  _GEN_15661 = _T_1530 ? _GEN_15653 : _GEN_14797; // @[sequencer-master.scala 168:32]
  wire  _GEN_15662 = _GEN_32729 | _GEN_14814; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15663 = _GEN_32730 | _GEN_14815; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15664 = _GEN_32731 | _GEN_14816; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15665 = _GEN_32732 | _GEN_14817; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15666 = _GEN_32733 | _GEN_14818; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15667 = _GEN_32734 | _GEN_14819; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15668 = _GEN_32735 | _GEN_14820; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15669 = _GEN_32736 | _GEN_14821; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15670 = _T_1552 ? _GEN_15662 : _GEN_14814; // @[sequencer-master.scala 168:32]
  wire  _GEN_15671 = _T_1552 ? _GEN_15663 : _GEN_14815; // @[sequencer-master.scala 168:32]
  wire  _GEN_15672 = _T_1552 ? _GEN_15664 : _GEN_14816; // @[sequencer-master.scala 168:32]
  wire  _GEN_15673 = _T_1552 ? _GEN_15665 : _GEN_14817; // @[sequencer-master.scala 168:32]
  wire  _GEN_15674 = _T_1552 ? _GEN_15666 : _GEN_14818; // @[sequencer-master.scala 168:32]
  wire  _GEN_15675 = _T_1552 ? _GEN_15667 : _GEN_14819; // @[sequencer-master.scala 168:32]
  wire  _GEN_15676 = _T_1552 ? _GEN_15668 : _GEN_14820; // @[sequencer-master.scala 168:32]
  wire  _GEN_15677 = _T_1552 ? _GEN_15669 : _GEN_14821; // @[sequencer-master.scala 168:32]
  wire  _GEN_15678 = _GEN_32729 | _GEN_14838; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15679 = _GEN_32730 | _GEN_14839; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15680 = _GEN_32731 | _GEN_14840; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15681 = _GEN_32732 | _GEN_14841; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15682 = _GEN_32733 | _GEN_14842; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15683 = _GEN_32734 | _GEN_14843; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15684 = _GEN_32735 | _GEN_14844; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15685 = _GEN_32736 | _GEN_14845; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15686 = _T_1574 ? _GEN_15678 : _GEN_14838; // @[sequencer-master.scala 168:32]
  wire  _GEN_15687 = _T_1574 ? _GEN_15679 : _GEN_14839; // @[sequencer-master.scala 168:32]
  wire  _GEN_15688 = _T_1574 ? _GEN_15680 : _GEN_14840; // @[sequencer-master.scala 168:32]
  wire  _GEN_15689 = _T_1574 ? _GEN_15681 : _GEN_14841; // @[sequencer-master.scala 168:32]
  wire  _GEN_15690 = _T_1574 ? _GEN_15682 : _GEN_14842; // @[sequencer-master.scala 168:32]
  wire  _GEN_15691 = _T_1574 ? _GEN_15683 : _GEN_14843; // @[sequencer-master.scala 168:32]
  wire  _GEN_15692 = _T_1574 ? _GEN_15684 : _GEN_14844; // @[sequencer-master.scala 168:32]
  wire  _GEN_15693 = _T_1574 ? _GEN_15685 : _GEN_14845; // @[sequencer-master.scala 168:32]
  wire  _GEN_15694 = _GEN_32729 | _GEN_14862; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15695 = _GEN_32730 | _GEN_14863; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15696 = _GEN_32731 | _GEN_14864; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15697 = _GEN_32732 | _GEN_14865; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15698 = _GEN_32733 | _GEN_14866; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15699 = _GEN_32734 | _GEN_14867; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15700 = _GEN_32735 | _GEN_14868; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15701 = _GEN_32736 | _GEN_14869; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_15702 = _T_1596 ? _GEN_15694 : _GEN_14862; // @[sequencer-master.scala 168:32]
  wire  _GEN_15703 = _T_1596 ? _GEN_15695 : _GEN_14863; // @[sequencer-master.scala 168:32]
  wire  _GEN_15704 = _T_1596 ? _GEN_15696 : _GEN_14864; // @[sequencer-master.scala 168:32]
  wire  _GEN_15705 = _T_1596 ? _GEN_15697 : _GEN_14865; // @[sequencer-master.scala 168:32]
  wire  _GEN_15706 = _T_1596 ? _GEN_15698 : _GEN_14866; // @[sequencer-master.scala 168:32]
  wire  _GEN_15707 = _T_1596 ? _GEN_15699 : _GEN_14867; // @[sequencer-master.scala 168:32]
  wire  _GEN_15708 = _T_1596 ? _GEN_15700 : _GEN_14868; // @[sequencer-master.scala 168:32]
  wire  _GEN_15709 = _T_1596 ? _GEN_15701 : _GEN_14869; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_15710 = 3'h0 == tail ? _T_1615[1:0] : _GEN_14588; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15711 = 3'h1 == tail ? _T_1615[1:0] : _GEN_14589; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15712 = 3'h2 == tail ? _T_1615[1:0] : _GEN_14590; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15713 = 3'h3 == tail ? _T_1615[1:0] : _GEN_14591; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15714 = 3'h4 == tail ? _T_1615[1:0] : _GEN_14592; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15715 = 3'h5 == tail ? _T_1615[1:0] : _GEN_14593; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15716 = 3'h6 == tail ? _T_1615[1:0] : _GEN_14594; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_15717 = 3'h7 == tail ? _T_1615[1:0] : _GEN_14595; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_15718 = 3'h0 == tail ? 4'h0 : _GEN_14596; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15719 = 3'h1 == tail ? 4'h0 : _GEN_14597; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15720 = 3'h2 == tail ? 4'h0 : _GEN_14598; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15721 = 3'h3 == tail ? 4'h0 : _GEN_14599; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15722 = 3'h4 == tail ? 4'h0 : _GEN_14600; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15723 = 3'h5 == tail ? 4'h0 : _GEN_14601; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15724 = 3'h6 == tail ? 4'h0 : _GEN_14602; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_15725 = 3'h7 == tail ? 4'h0 : _GEN_14603; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_15726 = 3'h0 == tail ? 3'h0 : _GEN_14604; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15727 = 3'h1 == tail ? 3'h0 : _GEN_14605; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15728 = 3'h2 == tail ? 3'h0 : _GEN_14606; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15729 = 3'h3 == tail ? 3'h0 : _GEN_14607; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15730 = 3'h4 == tail ? 3'h0 : _GEN_14608; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15731 = 3'h5 == tail ? 3'h0 : _GEN_14609; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15732 = 3'h6 == tail ? 3'h0 : _GEN_14610; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_15733 = 3'h7 == tail ? 3'h0 : _GEN_14611; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [3:0] _T_2177 = _T_1789[3:0] + 4'h3; // @[sequencer-master.scala 247:56]
  wire [3:0] _GEN_15734 = 3'h0 == tail ? _T_2177 : _GEN_15718; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15735 = 3'h1 == tail ? _T_2177 : _GEN_15719; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15736 = 3'h2 == tail ? _T_2177 : _GEN_15720; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15737 = 3'h3 == tail ? _T_2177 : _GEN_15721; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15738 = 3'h4 == tail ? _T_2177 : _GEN_15722; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15739 = 3'h5 == tail ? _T_2177 : _GEN_15723; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15740 = 3'h6 == tail ? _T_2177 : _GEN_15724; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15741 = 3'h7 == tail ? _T_2177 : _GEN_15725; // @[sequencer-master.scala 235:65 sequencer-master.scala 235:65]
  wire [3:0] _GEN_15742 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15734 : _GEN_15718; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15743 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15735 : _GEN_15719; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15744 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15736 : _GEN_15720; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15745 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15737 : _GEN_15721; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15746 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15738 : _GEN_15722; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15747 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15739 : _GEN_15723; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15748 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15740 : _GEN_15724; // @[sequencer-master.scala 235:47]
  wire [3:0] _GEN_15749 = ~(io_op_bits_base_vd_pred | io_op_bits_base_vd_scalar) ? _GEN_15741 : _GEN_15725; // @[sequencer-master.scala 235:47]
  wire [2:0] _GEN_15750 = 3'h0 == tail ? _T_2177[2:0] : _GEN_15726; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15751 = 3'h1 == tail ? _T_2177[2:0] : _GEN_15727; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15752 = 3'h2 == tail ? _T_2177[2:0] : _GEN_15728; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15753 = 3'h3 == tail ? _T_2177[2:0] : _GEN_15729; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15754 = 3'h4 == tail ? _T_2177[2:0] : _GEN_15730; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15755 = 3'h5 == tail ? _T_2177[2:0] : _GEN_15731; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15756 = 3'h6 == tail ? _T_2177[2:0] : _GEN_15732; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15757 = 3'h7 == tail ? _T_2177[2:0] : _GEN_15733; // @[sequencer-master.scala 236:63 sequencer-master.scala 236:63]
  wire [2:0] _GEN_15758 = io_op_bits_base_vd_pred ? _GEN_15750 : _GEN_15726; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15759 = io_op_bits_base_vd_pred ? _GEN_15751 : _GEN_15727; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15760 = io_op_bits_base_vd_pred ? _GEN_15752 : _GEN_15728; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15761 = io_op_bits_base_vd_pred ? _GEN_15753 : _GEN_15729; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15762 = io_op_bits_base_vd_pred ? _GEN_15754 : _GEN_15730; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15763 = io_op_bits_base_vd_pred ? _GEN_15755 : _GEN_15731; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15764 = io_op_bits_base_vd_pred ? _GEN_15756 : _GEN_15732; // @[sequencer-master.scala 236:45]
  wire [2:0] _GEN_15765 = io_op_bits_base_vd_pred ? _GEN_15757 : _GEN_15733; // @[sequencer-master.scala 236:45]
  wire  _GEN_15766 = io_op_bits_active_vfconv ? _GEN_14614 : _GEN_14132; // @[sequencer-master.scala 647:41]
  wire  _GEN_15767 = io_op_bits_active_vfconv ? _GEN_14615 : _GEN_14133; // @[sequencer-master.scala 647:41]
  wire  _GEN_15768 = io_op_bits_active_vfconv ? _GEN_14616 : _GEN_14134; // @[sequencer-master.scala 647:41]
  wire  _GEN_15769 = io_op_bits_active_vfconv ? _GEN_14617 : _GEN_14135; // @[sequencer-master.scala 647:41]
  wire  _GEN_15770 = io_op_bits_active_vfconv ? _GEN_14618 : _GEN_14136; // @[sequencer-master.scala 647:41]
  wire  _GEN_15771 = io_op_bits_active_vfconv ? _GEN_14619 : _GEN_14137; // @[sequencer-master.scala 647:41]
  wire  _GEN_15772 = io_op_bits_active_vfconv ? _GEN_14620 : _GEN_14138; // @[sequencer-master.scala 647:41]
  wire  _GEN_15773 = io_op_bits_active_vfconv ? _GEN_14621 : _GEN_14139; // @[sequencer-master.scala 647:41]
  wire  _GEN_15782 = io_op_bits_active_vfconv ? _GEN_14950 : _GEN_14148; // @[sequencer-master.scala 647:41]
  wire  _GEN_15783 = io_op_bits_active_vfconv ? _GEN_14951 : _GEN_14149; // @[sequencer-master.scala 647:41]
  wire  _GEN_15784 = io_op_bits_active_vfconv ? _GEN_14952 : _GEN_14150; // @[sequencer-master.scala 647:41]
  wire  _GEN_15785 = io_op_bits_active_vfconv ? _GEN_14953 : _GEN_14151; // @[sequencer-master.scala 647:41]
  wire  _GEN_15786 = io_op_bits_active_vfconv ? _GEN_14954 : _GEN_14152; // @[sequencer-master.scala 647:41]
  wire  _GEN_15787 = io_op_bits_active_vfconv ? _GEN_14955 : _GEN_14153; // @[sequencer-master.scala 647:41]
  wire  _GEN_15788 = io_op_bits_active_vfconv ? _GEN_14956 : _GEN_14154; // @[sequencer-master.scala 647:41]
  wire  _GEN_15789 = io_op_bits_active_vfconv ? _GEN_14957 : _GEN_14155; // @[sequencer-master.scala 647:41]
  wire  _GEN_15790 = io_op_bits_active_vfconv ? _GEN_15182 : _GEN_14156; // @[sequencer-master.scala 647:41]
  wire  _GEN_15791 = io_op_bits_active_vfconv ? _GEN_15183 : _GEN_14157; // @[sequencer-master.scala 647:41]
  wire  _GEN_15792 = io_op_bits_active_vfconv ? _GEN_15184 : _GEN_14158; // @[sequencer-master.scala 647:41]
  wire  _GEN_15793 = io_op_bits_active_vfconv ? _GEN_15185 : _GEN_14159; // @[sequencer-master.scala 647:41]
  wire  _GEN_15794 = io_op_bits_active_vfconv ? _GEN_15186 : _GEN_14160; // @[sequencer-master.scala 647:41]
  wire  _GEN_15795 = io_op_bits_active_vfconv ? _GEN_15187 : _GEN_14161; // @[sequencer-master.scala 647:41]
  wire  _GEN_15796 = io_op_bits_active_vfconv ? _GEN_15188 : _GEN_14162; // @[sequencer-master.scala 647:41]
  wire  _GEN_15797 = io_op_bits_active_vfconv ? _GEN_15189 : _GEN_14163; // @[sequencer-master.scala 647:41]
  wire  _GEN_15798 = io_op_bits_active_vfconv ? _GEN_14646 : _GEN_14164; // @[sequencer-master.scala 647:41]
  wire  _GEN_15799 = io_op_bits_active_vfconv ? _GEN_14647 : _GEN_14165; // @[sequencer-master.scala 647:41]
  wire  _GEN_15800 = io_op_bits_active_vfconv ? _GEN_14648 : _GEN_14166; // @[sequencer-master.scala 647:41]
  wire  _GEN_15801 = io_op_bits_active_vfconv ? _GEN_14649 : _GEN_14167; // @[sequencer-master.scala 647:41]
  wire  _GEN_15802 = io_op_bits_active_vfconv ? _GEN_14650 : _GEN_14168; // @[sequencer-master.scala 647:41]
  wire  _GEN_15803 = io_op_bits_active_vfconv ? _GEN_14651 : _GEN_14169; // @[sequencer-master.scala 647:41]
  wire  _GEN_15804 = io_op_bits_active_vfconv ? _GEN_14652 : _GEN_14170; // @[sequencer-master.scala 647:41]
  wire  _GEN_15805 = io_op_bits_active_vfconv ? _GEN_14653 : _GEN_14171; // @[sequencer-master.scala 647:41]
  wire  _GEN_15806 = io_op_bits_active_vfconv ? _GEN_14654 : _GEN_14172; // @[sequencer-master.scala 647:41]
  wire  _GEN_15807 = io_op_bits_active_vfconv ? _GEN_14655 : _GEN_14173; // @[sequencer-master.scala 647:41]
  wire  _GEN_15808 = io_op_bits_active_vfconv ? _GEN_14656 : _GEN_14174; // @[sequencer-master.scala 647:41]
  wire  _GEN_15809 = io_op_bits_active_vfconv ? _GEN_14657 : _GEN_14175; // @[sequencer-master.scala 647:41]
  wire  _GEN_15810 = io_op_bits_active_vfconv ? _GEN_14658 : _GEN_14176; // @[sequencer-master.scala 647:41]
  wire  _GEN_15811 = io_op_bits_active_vfconv ? _GEN_14659 : _GEN_14177; // @[sequencer-master.scala 647:41]
  wire  _GEN_15812 = io_op_bits_active_vfconv ? _GEN_14660 : _GEN_14178; // @[sequencer-master.scala 647:41]
  wire  _GEN_15813 = io_op_bits_active_vfconv ? _GEN_14661 : _GEN_14179; // @[sequencer-master.scala 647:41]
  wire  _GEN_15814 = io_op_bits_active_vfconv ? _GEN_15414 : _GEN_14180; // @[sequencer-master.scala 647:41]
  wire  _GEN_15815 = io_op_bits_active_vfconv ? _GEN_15415 : _GEN_14181; // @[sequencer-master.scala 647:41]
  wire  _GEN_15816 = io_op_bits_active_vfconv ? _GEN_15416 : _GEN_14182; // @[sequencer-master.scala 647:41]
  wire  _GEN_15817 = io_op_bits_active_vfconv ? _GEN_15417 : _GEN_14183; // @[sequencer-master.scala 647:41]
  wire  _GEN_15818 = io_op_bits_active_vfconv ? _GEN_15418 : _GEN_14184; // @[sequencer-master.scala 647:41]
  wire  _GEN_15819 = io_op_bits_active_vfconv ? _GEN_15419 : _GEN_14185; // @[sequencer-master.scala 647:41]
  wire  _GEN_15820 = io_op_bits_active_vfconv ? _GEN_15420 : _GEN_14186; // @[sequencer-master.scala 647:41]
  wire  _GEN_15821 = io_op_bits_active_vfconv ? _GEN_15421 : _GEN_14187; // @[sequencer-master.scala 647:41]
  wire  _GEN_15822 = io_op_bits_active_vfconv ? _GEN_14670 : _GEN_14188; // @[sequencer-master.scala 647:41]
  wire  _GEN_15823 = io_op_bits_active_vfconv ? _GEN_14671 : _GEN_14189; // @[sequencer-master.scala 647:41]
  wire  _GEN_15824 = io_op_bits_active_vfconv ? _GEN_14672 : _GEN_14190; // @[sequencer-master.scala 647:41]
  wire  _GEN_15825 = io_op_bits_active_vfconv ? _GEN_14673 : _GEN_14191; // @[sequencer-master.scala 647:41]
  wire  _GEN_15826 = io_op_bits_active_vfconv ? _GEN_14674 : _GEN_14192; // @[sequencer-master.scala 647:41]
  wire  _GEN_15827 = io_op_bits_active_vfconv ? _GEN_14675 : _GEN_14193; // @[sequencer-master.scala 647:41]
  wire  _GEN_15828 = io_op_bits_active_vfconv ? _GEN_14676 : _GEN_14194; // @[sequencer-master.scala 647:41]
  wire  _GEN_15829 = io_op_bits_active_vfconv ? _GEN_14677 : _GEN_14195; // @[sequencer-master.scala 647:41]
  wire  _GEN_15830 = io_op_bits_active_vfconv ? _GEN_15238 : _GEN_14196; // @[sequencer-master.scala 647:41]
  wire  _GEN_15831 = io_op_bits_active_vfconv ? _GEN_15239 : _GEN_14197; // @[sequencer-master.scala 647:41]
  wire  _GEN_15832 = io_op_bits_active_vfconv ? _GEN_15240 : _GEN_14198; // @[sequencer-master.scala 647:41]
  wire  _GEN_15833 = io_op_bits_active_vfconv ? _GEN_15241 : _GEN_14199; // @[sequencer-master.scala 647:41]
  wire  _GEN_15834 = io_op_bits_active_vfconv ? _GEN_15242 : _GEN_14200; // @[sequencer-master.scala 647:41]
  wire  _GEN_15835 = io_op_bits_active_vfconv ? _GEN_15243 : _GEN_14201; // @[sequencer-master.scala 647:41]
  wire  _GEN_15836 = io_op_bits_active_vfconv ? _GEN_15244 : _GEN_14202; // @[sequencer-master.scala 647:41]
  wire  _GEN_15837 = io_op_bits_active_vfconv ? _GEN_15245 : _GEN_14203; // @[sequencer-master.scala 647:41]
  wire  _GEN_15838 = io_op_bits_active_vfconv ? _GEN_15462 : _GEN_14204; // @[sequencer-master.scala 647:41]
  wire  _GEN_15839 = io_op_bits_active_vfconv ? _GEN_15463 : _GEN_14205; // @[sequencer-master.scala 647:41]
  wire  _GEN_15840 = io_op_bits_active_vfconv ? _GEN_15464 : _GEN_14206; // @[sequencer-master.scala 647:41]
  wire  _GEN_15841 = io_op_bits_active_vfconv ? _GEN_15465 : _GEN_14207; // @[sequencer-master.scala 647:41]
  wire  _GEN_15842 = io_op_bits_active_vfconv ? _GEN_15466 : _GEN_14208; // @[sequencer-master.scala 647:41]
  wire  _GEN_15843 = io_op_bits_active_vfconv ? _GEN_15467 : _GEN_14209; // @[sequencer-master.scala 647:41]
  wire  _GEN_15844 = io_op_bits_active_vfconv ? _GEN_15468 : _GEN_14210; // @[sequencer-master.scala 647:41]
  wire  _GEN_15845 = io_op_bits_active_vfconv ? _GEN_15469 : _GEN_14211; // @[sequencer-master.scala 647:41]
  wire  _GEN_15846 = io_op_bits_active_vfconv ? _GEN_15590 : _GEN_14212; // @[sequencer-master.scala 647:41]
  wire  _GEN_15847 = io_op_bits_active_vfconv ? _GEN_15591 : _GEN_14213; // @[sequencer-master.scala 647:41]
  wire  _GEN_15848 = io_op_bits_active_vfconv ? _GEN_15592 : _GEN_14214; // @[sequencer-master.scala 647:41]
  wire  _GEN_15849 = io_op_bits_active_vfconv ? _GEN_15593 : _GEN_14215; // @[sequencer-master.scala 647:41]
  wire  _GEN_15850 = io_op_bits_active_vfconv ? _GEN_15594 : _GEN_14216; // @[sequencer-master.scala 647:41]
  wire  _GEN_15851 = io_op_bits_active_vfconv ? _GEN_15595 : _GEN_14217; // @[sequencer-master.scala 647:41]
  wire  _GEN_15852 = io_op_bits_active_vfconv ? _GEN_15596 : _GEN_14218; // @[sequencer-master.scala 647:41]
  wire  _GEN_15853 = io_op_bits_active_vfconv ? _GEN_15597 : _GEN_14219; // @[sequencer-master.scala 647:41]
  wire  _GEN_15854 = io_op_bits_active_vfconv ? _GEN_15254 : _GEN_14220; // @[sequencer-master.scala 647:41]
  wire  _GEN_15855 = io_op_bits_active_vfconv ? _GEN_15255 : _GEN_14221; // @[sequencer-master.scala 647:41]
  wire  _GEN_15856 = io_op_bits_active_vfconv ? _GEN_15256 : _GEN_14222; // @[sequencer-master.scala 647:41]
  wire  _GEN_15857 = io_op_bits_active_vfconv ? _GEN_15257 : _GEN_14223; // @[sequencer-master.scala 647:41]
  wire  _GEN_15858 = io_op_bits_active_vfconv ? _GEN_15258 : _GEN_14224; // @[sequencer-master.scala 647:41]
  wire  _GEN_15859 = io_op_bits_active_vfconv ? _GEN_15259 : _GEN_14225; // @[sequencer-master.scala 647:41]
  wire  _GEN_15860 = io_op_bits_active_vfconv ? _GEN_15260 : _GEN_14226; // @[sequencer-master.scala 647:41]
  wire  _GEN_15861 = io_op_bits_active_vfconv ? _GEN_15261 : _GEN_14227; // @[sequencer-master.scala 647:41]
  wire  _GEN_15862 = io_op_bits_active_vfconv ? _GEN_15478 : _GEN_14228; // @[sequencer-master.scala 647:41]
  wire  _GEN_15863 = io_op_bits_active_vfconv ? _GEN_15479 : _GEN_14229; // @[sequencer-master.scala 647:41]
  wire  _GEN_15864 = io_op_bits_active_vfconv ? _GEN_15480 : _GEN_14230; // @[sequencer-master.scala 647:41]
  wire  _GEN_15865 = io_op_bits_active_vfconv ? _GEN_15481 : _GEN_14231; // @[sequencer-master.scala 647:41]
  wire  _GEN_15866 = io_op_bits_active_vfconv ? _GEN_15482 : _GEN_14232; // @[sequencer-master.scala 647:41]
  wire  _GEN_15867 = io_op_bits_active_vfconv ? _GEN_15483 : _GEN_14233; // @[sequencer-master.scala 647:41]
  wire  _GEN_15868 = io_op_bits_active_vfconv ? _GEN_15484 : _GEN_14234; // @[sequencer-master.scala 647:41]
  wire  _GEN_15869 = io_op_bits_active_vfconv ? _GEN_15485 : _GEN_14235; // @[sequencer-master.scala 647:41]
  wire  _GEN_15870 = io_op_bits_active_vfconv ? _GEN_15606 : _GEN_14236; // @[sequencer-master.scala 647:41]
  wire  _GEN_15871 = io_op_bits_active_vfconv ? _GEN_15607 : _GEN_14237; // @[sequencer-master.scala 647:41]
  wire  _GEN_15872 = io_op_bits_active_vfconv ? _GEN_15608 : _GEN_14238; // @[sequencer-master.scala 647:41]
  wire  _GEN_15873 = io_op_bits_active_vfconv ? _GEN_15609 : _GEN_14239; // @[sequencer-master.scala 647:41]
  wire  _GEN_15874 = io_op_bits_active_vfconv ? _GEN_15610 : _GEN_14240; // @[sequencer-master.scala 647:41]
  wire  _GEN_15875 = io_op_bits_active_vfconv ? _GEN_15611 : _GEN_14241; // @[sequencer-master.scala 647:41]
  wire  _GEN_15876 = io_op_bits_active_vfconv ? _GEN_15612 : _GEN_14242; // @[sequencer-master.scala 647:41]
  wire  _GEN_15877 = io_op_bits_active_vfconv ? _GEN_15613 : _GEN_14243; // @[sequencer-master.scala 647:41]
  wire  _GEN_15878 = io_op_bits_active_vfconv ? _GEN_15270 : _GEN_14244; // @[sequencer-master.scala 647:41]
  wire  _GEN_15879 = io_op_bits_active_vfconv ? _GEN_15271 : _GEN_14245; // @[sequencer-master.scala 647:41]
  wire  _GEN_15880 = io_op_bits_active_vfconv ? _GEN_15272 : _GEN_14246; // @[sequencer-master.scala 647:41]
  wire  _GEN_15881 = io_op_bits_active_vfconv ? _GEN_15273 : _GEN_14247; // @[sequencer-master.scala 647:41]
  wire  _GEN_15882 = io_op_bits_active_vfconv ? _GEN_15274 : _GEN_14248; // @[sequencer-master.scala 647:41]
  wire  _GEN_15883 = io_op_bits_active_vfconv ? _GEN_15275 : _GEN_14249; // @[sequencer-master.scala 647:41]
  wire  _GEN_15884 = io_op_bits_active_vfconv ? _GEN_15276 : _GEN_14250; // @[sequencer-master.scala 647:41]
  wire  _GEN_15885 = io_op_bits_active_vfconv ? _GEN_15277 : _GEN_14251; // @[sequencer-master.scala 647:41]
  wire  _GEN_15886 = io_op_bits_active_vfconv ? _GEN_15494 : _GEN_14252; // @[sequencer-master.scala 647:41]
  wire  _GEN_15887 = io_op_bits_active_vfconv ? _GEN_15495 : _GEN_14253; // @[sequencer-master.scala 647:41]
  wire  _GEN_15888 = io_op_bits_active_vfconv ? _GEN_15496 : _GEN_14254; // @[sequencer-master.scala 647:41]
  wire  _GEN_15889 = io_op_bits_active_vfconv ? _GEN_15497 : _GEN_14255; // @[sequencer-master.scala 647:41]
  wire  _GEN_15890 = io_op_bits_active_vfconv ? _GEN_15498 : _GEN_14256; // @[sequencer-master.scala 647:41]
  wire  _GEN_15891 = io_op_bits_active_vfconv ? _GEN_15499 : _GEN_14257; // @[sequencer-master.scala 647:41]
  wire  _GEN_15892 = io_op_bits_active_vfconv ? _GEN_15500 : _GEN_14258; // @[sequencer-master.scala 647:41]
  wire  _GEN_15893 = io_op_bits_active_vfconv ? _GEN_15501 : _GEN_14259; // @[sequencer-master.scala 647:41]
  wire  _GEN_15894 = io_op_bits_active_vfconv ? _GEN_15622 : _GEN_14260; // @[sequencer-master.scala 647:41]
  wire  _GEN_15895 = io_op_bits_active_vfconv ? _GEN_15623 : _GEN_14261; // @[sequencer-master.scala 647:41]
  wire  _GEN_15896 = io_op_bits_active_vfconv ? _GEN_15624 : _GEN_14262; // @[sequencer-master.scala 647:41]
  wire  _GEN_15897 = io_op_bits_active_vfconv ? _GEN_15625 : _GEN_14263; // @[sequencer-master.scala 647:41]
  wire  _GEN_15898 = io_op_bits_active_vfconv ? _GEN_15626 : _GEN_14264; // @[sequencer-master.scala 647:41]
  wire  _GEN_15899 = io_op_bits_active_vfconv ? _GEN_15627 : _GEN_14265; // @[sequencer-master.scala 647:41]
  wire  _GEN_15900 = io_op_bits_active_vfconv ? _GEN_15628 : _GEN_14266; // @[sequencer-master.scala 647:41]
  wire  _GEN_15901 = io_op_bits_active_vfconv ? _GEN_15629 : _GEN_14267; // @[sequencer-master.scala 647:41]
  wire  _GEN_15902 = io_op_bits_active_vfconv ? _GEN_15286 : _GEN_14268; // @[sequencer-master.scala 647:41]
  wire  _GEN_15903 = io_op_bits_active_vfconv ? _GEN_15287 : _GEN_14269; // @[sequencer-master.scala 647:41]
  wire  _GEN_15904 = io_op_bits_active_vfconv ? _GEN_15288 : _GEN_14270; // @[sequencer-master.scala 647:41]
  wire  _GEN_15905 = io_op_bits_active_vfconv ? _GEN_15289 : _GEN_14271; // @[sequencer-master.scala 647:41]
  wire  _GEN_15906 = io_op_bits_active_vfconv ? _GEN_15290 : _GEN_14272; // @[sequencer-master.scala 647:41]
  wire  _GEN_15907 = io_op_bits_active_vfconv ? _GEN_15291 : _GEN_14273; // @[sequencer-master.scala 647:41]
  wire  _GEN_15908 = io_op_bits_active_vfconv ? _GEN_15292 : _GEN_14274; // @[sequencer-master.scala 647:41]
  wire  _GEN_15909 = io_op_bits_active_vfconv ? _GEN_15293 : _GEN_14275; // @[sequencer-master.scala 647:41]
  wire  _GEN_15910 = io_op_bits_active_vfconv ? _GEN_15510 : _GEN_14276; // @[sequencer-master.scala 647:41]
  wire  _GEN_15911 = io_op_bits_active_vfconv ? _GEN_15511 : _GEN_14277; // @[sequencer-master.scala 647:41]
  wire  _GEN_15912 = io_op_bits_active_vfconv ? _GEN_15512 : _GEN_14278; // @[sequencer-master.scala 647:41]
  wire  _GEN_15913 = io_op_bits_active_vfconv ? _GEN_15513 : _GEN_14279; // @[sequencer-master.scala 647:41]
  wire  _GEN_15914 = io_op_bits_active_vfconv ? _GEN_15514 : _GEN_14280; // @[sequencer-master.scala 647:41]
  wire  _GEN_15915 = io_op_bits_active_vfconv ? _GEN_15515 : _GEN_14281; // @[sequencer-master.scala 647:41]
  wire  _GEN_15916 = io_op_bits_active_vfconv ? _GEN_15516 : _GEN_14282; // @[sequencer-master.scala 647:41]
  wire  _GEN_15917 = io_op_bits_active_vfconv ? _GEN_15517 : _GEN_14283; // @[sequencer-master.scala 647:41]
  wire  _GEN_15918 = io_op_bits_active_vfconv ? _GEN_15638 : _GEN_14284; // @[sequencer-master.scala 647:41]
  wire  _GEN_15919 = io_op_bits_active_vfconv ? _GEN_15639 : _GEN_14285; // @[sequencer-master.scala 647:41]
  wire  _GEN_15920 = io_op_bits_active_vfconv ? _GEN_15640 : _GEN_14286; // @[sequencer-master.scala 647:41]
  wire  _GEN_15921 = io_op_bits_active_vfconv ? _GEN_15641 : _GEN_14287; // @[sequencer-master.scala 647:41]
  wire  _GEN_15922 = io_op_bits_active_vfconv ? _GEN_15642 : _GEN_14288; // @[sequencer-master.scala 647:41]
  wire  _GEN_15923 = io_op_bits_active_vfconv ? _GEN_15643 : _GEN_14289; // @[sequencer-master.scala 647:41]
  wire  _GEN_15924 = io_op_bits_active_vfconv ? _GEN_15644 : _GEN_14290; // @[sequencer-master.scala 647:41]
  wire  _GEN_15925 = io_op_bits_active_vfconv ? _GEN_15645 : _GEN_14291; // @[sequencer-master.scala 647:41]
  wire  _GEN_15926 = io_op_bits_active_vfconv ? _GEN_15302 : _GEN_14292; // @[sequencer-master.scala 647:41]
  wire  _GEN_15927 = io_op_bits_active_vfconv ? _GEN_15303 : _GEN_14293; // @[sequencer-master.scala 647:41]
  wire  _GEN_15928 = io_op_bits_active_vfconv ? _GEN_15304 : _GEN_14294; // @[sequencer-master.scala 647:41]
  wire  _GEN_15929 = io_op_bits_active_vfconv ? _GEN_15305 : _GEN_14295; // @[sequencer-master.scala 647:41]
  wire  _GEN_15930 = io_op_bits_active_vfconv ? _GEN_15306 : _GEN_14296; // @[sequencer-master.scala 647:41]
  wire  _GEN_15931 = io_op_bits_active_vfconv ? _GEN_15307 : _GEN_14297; // @[sequencer-master.scala 647:41]
  wire  _GEN_15932 = io_op_bits_active_vfconv ? _GEN_15308 : _GEN_14298; // @[sequencer-master.scala 647:41]
  wire  _GEN_15933 = io_op_bits_active_vfconv ? _GEN_15309 : _GEN_14299; // @[sequencer-master.scala 647:41]
  wire  _GEN_15934 = io_op_bits_active_vfconv ? _GEN_15526 : _GEN_14300; // @[sequencer-master.scala 647:41]
  wire  _GEN_15935 = io_op_bits_active_vfconv ? _GEN_15527 : _GEN_14301; // @[sequencer-master.scala 647:41]
  wire  _GEN_15936 = io_op_bits_active_vfconv ? _GEN_15528 : _GEN_14302; // @[sequencer-master.scala 647:41]
  wire  _GEN_15937 = io_op_bits_active_vfconv ? _GEN_15529 : _GEN_14303; // @[sequencer-master.scala 647:41]
  wire  _GEN_15938 = io_op_bits_active_vfconv ? _GEN_15530 : _GEN_14304; // @[sequencer-master.scala 647:41]
  wire  _GEN_15939 = io_op_bits_active_vfconv ? _GEN_15531 : _GEN_14305; // @[sequencer-master.scala 647:41]
  wire  _GEN_15940 = io_op_bits_active_vfconv ? _GEN_15532 : _GEN_14306; // @[sequencer-master.scala 647:41]
  wire  _GEN_15941 = io_op_bits_active_vfconv ? _GEN_15533 : _GEN_14307; // @[sequencer-master.scala 647:41]
  wire  _GEN_15942 = io_op_bits_active_vfconv ? _GEN_15654 : _GEN_14308; // @[sequencer-master.scala 647:41]
  wire  _GEN_15943 = io_op_bits_active_vfconv ? _GEN_15655 : _GEN_14309; // @[sequencer-master.scala 647:41]
  wire  _GEN_15944 = io_op_bits_active_vfconv ? _GEN_15656 : _GEN_14310; // @[sequencer-master.scala 647:41]
  wire  _GEN_15945 = io_op_bits_active_vfconv ? _GEN_15657 : _GEN_14311; // @[sequencer-master.scala 647:41]
  wire  _GEN_15946 = io_op_bits_active_vfconv ? _GEN_15658 : _GEN_14312; // @[sequencer-master.scala 647:41]
  wire  _GEN_15947 = io_op_bits_active_vfconv ? _GEN_15659 : _GEN_14313; // @[sequencer-master.scala 647:41]
  wire  _GEN_15948 = io_op_bits_active_vfconv ? _GEN_15660 : _GEN_14314; // @[sequencer-master.scala 647:41]
  wire  _GEN_15949 = io_op_bits_active_vfconv ? _GEN_15661 : _GEN_14315; // @[sequencer-master.scala 647:41]
  wire  _GEN_15950 = io_op_bits_active_vfconv ? _GEN_15318 : _GEN_14316; // @[sequencer-master.scala 647:41]
  wire  _GEN_15951 = io_op_bits_active_vfconv ? _GEN_15319 : _GEN_14317; // @[sequencer-master.scala 647:41]
  wire  _GEN_15952 = io_op_bits_active_vfconv ? _GEN_15320 : _GEN_14318; // @[sequencer-master.scala 647:41]
  wire  _GEN_15953 = io_op_bits_active_vfconv ? _GEN_15321 : _GEN_14319; // @[sequencer-master.scala 647:41]
  wire  _GEN_15954 = io_op_bits_active_vfconv ? _GEN_15322 : _GEN_14320; // @[sequencer-master.scala 647:41]
  wire  _GEN_15955 = io_op_bits_active_vfconv ? _GEN_15323 : _GEN_14321; // @[sequencer-master.scala 647:41]
  wire  _GEN_15956 = io_op_bits_active_vfconv ? _GEN_15324 : _GEN_14322; // @[sequencer-master.scala 647:41]
  wire  _GEN_15957 = io_op_bits_active_vfconv ? _GEN_15325 : _GEN_14323; // @[sequencer-master.scala 647:41]
  wire  _GEN_15958 = io_op_bits_active_vfconv ? _GEN_15542 : _GEN_14324; // @[sequencer-master.scala 647:41]
  wire  _GEN_15959 = io_op_bits_active_vfconv ? _GEN_15543 : _GEN_14325; // @[sequencer-master.scala 647:41]
  wire  _GEN_15960 = io_op_bits_active_vfconv ? _GEN_15544 : _GEN_14326; // @[sequencer-master.scala 647:41]
  wire  _GEN_15961 = io_op_bits_active_vfconv ? _GEN_15545 : _GEN_14327; // @[sequencer-master.scala 647:41]
  wire  _GEN_15962 = io_op_bits_active_vfconv ? _GEN_15546 : _GEN_14328; // @[sequencer-master.scala 647:41]
  wire  _GEN_15963 = io_op_bits_active_vfconv ? _GEN_15547 : _GEN_14329; // @[sequencer-master.scala 647:41]
  wire  _GEN_15964 = io_op_bits_active_vfconv ? _GEN_15548 : _GEN_14330; // @[sequencer-master.scala 647:41]
  wire  _GEN_15965 = io_op_bits_active_vfconv ? _GEN_15549 : _GEN_14331; // @[sequencer-master.scala 647:41]
  wire  _GEN_15966 = io_op_bits_active_vfconv ? _GEN_15670 : _GEN_14332; // @[sequencer-master.scala 647:41]
  wire  _GEN_15967 = io_op_bits_active_vfconv ? _GEN_15671 : _GEN_14333; // @[sequencer-master.scala 647:41]
  wire  _GEN_15968 = io_op_bits_active_vfconv ? _GEN_15672 : _GEN_14334; // @[sequencer-master.scala 647:41]
  wire  _GEN_15969 = io_op_bits_active_vfconv ? _GEN_15673 : _GEN_14335; // @[sequencer-master.scala 647:41]
  wire  _GEN_15970 = io_op_bits_active_vfconv ? _GEN_15674 : _GEN_14336; // @[sequencer-master.scala 647:41]
  wire  _GEN_15971 = io_op_bits_active_vfconv ? _GEN_15675 : _GEN_14337; // @[sequencer-master.scala 647:41]
  wire  _GEN_15972 = io_op_bits_active_vfconv ? _GEN_15676 : _GEN_14338; // @[sequencer-master.scala 647:41]
  wire  _GEN_15973 = io_op_bits_active_vfconv ? _GEN_15677 : _GEN_14339; // @[sequencer-master.scala 647:41]
  wire  _GEN_15974 = io_op_bits_active_vfconv ? _GEN_15334 : _GEN_14340; // @[sequencer-master.scala 647:41]
  wire  _GEN_15975 = io_op_bits_active_vfconv ? _GEN_15335 : _GEN_14341; // @[sequencer-master.scala 647:41]
  wire  _GEN_15976 = io_op_bits_active_vfconv ? _GEN_15336 : _GEN_14342; // @[sequencer-master.scala 647:41]
  wire  _GEN_15977 = io_op_bits_active_vfconv ? _GEN_15337 : _GEN_14343; // @[sequencer-master.scala 647:41]
  wire  _GEN_15978 = io_op_bits_active_vfconv ? _GEN_15338 : _GEN_14344; // @[sequencer-master.scala 647:41]
  wire  _GEN_15979 = io_op_bits_active_vfconv ? _GEN_15339 : _GEN_14345; // @[sequencer-master.scala 647:41]
  wire  _GEN_15980 = io_op_bits_active_vfconv ? _GEN_15340 : _GEN_14346; // @[sequencer-master.scala 647:41]
  wire  _GEN_15981 = io_op_bits_active_vfconv ? _GEN_15341 : _GEN_14347; // @[sequencer-master.scala 647:41]
  wire  _GEN_15982 = io_op_bits_active_vfconv ? _GEN_15558 : _GEN_14348; // @[sequencer-master.scala 647:41]
  wire  _GEN_15983 = io_op_bits_active_vfconv ? _GEN_15559 : _GEN_14349; // @[sequencer-master.scala 647:41]
  wire  _GEN_15984 = io_op_bits_active_vfconv ? _GEN_15560 : _GEN_14350; // @[sequencer-master.scala 647:41]
  wire  _GEN_15985 = io_op_bits_active_vfconv ? _GEN_15561 : _GEN_14351; // @[sequencer-master.scala 647:41]
  wire  _GEN_15986 = io_op_bits_active_vfconv ? _GEN_15562 : _GEN_14352; // @[sequencer-master.scala 647:41]
  wire  _GEN_15987 = io_op_bits_active_vfconv ? _GEN_15563 : _GEN_14353; // @[sequencer-master.scala 647:41]
  wire  _GEN_15988 = io_op_bits_active_vfconv ? _GEN_15564 : _GEN_14354; // @[sequencer-master.scala 647:41]
  wire  _GEN_15989 = io_op_bits_active_vfconv ? _GEN_15565 : _GEN_14355; // @[sequencer-master.scala 647:41]
  wire  _GEN_15990 = io_op_bits_active_vfconv ? _GEN_15686 : _GEN_14356; // @[sequencer-master.scala 647:41]
  wire  _GEN_15991 = io_op_bits_active_vfconv ? _GEN_15687 : _GEN_14357; // @[sequencer-master.scala 647:41]
  wire  _GEN_15992 = io_op_bits_active_vfconv ? _GEN_15688 : _GEN_14358; // @[sequencer-master.scala 647:41]
  wire  _GEN_15993 = io_op_bits_active_vfconv ? _GEN_15689 : _GEN_14359; // @[sequencer-master.scala 647:41]
  wire  _GEN_15994 = io_op_bits_active_vfconv ? _GEN_15690 : _GEN_14360; // @[sequencer-master.scala 647:41]
  wire  _GEN_15995 = io_op_bits_active_vfconv ? _GEN_15691 : _GEN_14361; // @[sequencer-master.scala 647:41]
  wire  _GEN_15996 = io_op_bits_active_vfconv ? _GEN_15692 : _GEN_14362; // @[sequencer-master.scala 647:41]
  wire  _GEN_15997 = io_op_bits_active_vfconv ? _GEN_15693 : _GEN_14363; // @[sequencer-master.scala 647:41]
  wire  _GEN_15998 = io_op_bits_active_vfconv ? _GEN_15350 : _GEN_14364; // @[sequencer-master.scala 647:41]
  wire  _GEN_15999 = io_op_bits_active_vfconv ? _GEN_15351 : _GEN_14365; // @[sequencer-master.scala 647:41]
  wire  _GEN_16000 = io_op_bits_active_vfconv ? _GEN_15352 : _GEN_14366; // @[sequencer-master.scala 647:41]
  wire  _GEN_16001 = io_op_bits_active_vfconv ? _GEN_15353 : _GEN_14367; // @[sequencer-master.scala 647:41]
  wire  _GEN_16002 = io_op_bits_active_vfconv ? _GEN_15354 : _GEN_14368; // @[sequencer-master.scala 647:41]
  wire  _GEN_16003 = io_op_bits_active_vfconv ? _GEN_15355 : _GEN_14369; // @[sequencer-master.scala 647:41]
  wire  _GEN_16004 = io_op_bits_active_vfconv ? _GEN_15356 : _GEN_14370; // @[sequencer-master.scala 647:41]
  wire  _GEN_16005 = io_op_bits_active_vfconv ? _GEN_15357 : _GEN_14371; // @[sequencer-master.scala 647:41]
  wire  _GEN_16006 = io_op_bits_active_vfconv ? _GEN_15574 : _GEN_14372; // @[sequencer-master.scala 647:41]
  wire  _GEN_16007 = io_op_bits_active_vfconv ? _GEN_15575 : _GEN_14373; // @[sequencer-master.scala 647:41]
  wire  _GEN_16008 = io_op_bits_active_vfconv ? _GEN_15576 : _GEN_14374; // @[sequencer-master.scala 647:41]
  wire  _GEN_16009 = io_op_bits_active_vfconv ? _GEN_15577 : _GEN_14375; // @[sequencer-master.scala 647:41]
  wire  _GEN_16010 = io_op_bits_active_vfconv ? _GEN_15578 : _GEN_14376; // @[sequencer-master.scala 647:41]
  wire  _GEN_16011 = io_op_bits_active_vfconv ? _GEN_15579 : _GEN_14377; // @[sequencer-master.scala 647:41]
  wire  _GEN_16012 = io_op_bits_active_vfconv ? _GEN_15580 : _GEN_14378; // @[sequencer-master.scala 647:41]
  wire  _GEN_16013 = io_op_bits_active_vfconv ? _GEN_15581 : _GEN_14379; // @[sequencer-master.scala 647:41]
  wire  _GEN_16014 = io_op_bits_active_vfconv ? _GEN_15702 : _GEN_14380; // @[sequencer-master.scala 647:41]
  wire  _GEN_16015 = io_op_bits_active_vfconv ? _GEN_15703 : _GEN_14381; // @[sequencer-master.scala 647:41]
  wire  _GEN_16016 = io_op_bits_active_vfconv ? _GEN_15704 : _GEN_14382; // @[sequencer-master.scala 647:41]
  wire  _GEN_16017 = io_op_bits_active_vfconv ? _GEN_15705 : _GEN_14383; // @[sequencer-master.scala 647:41]
  wire  _GEN_16018 = io_op_bits_active_vfconv ? _GEN_15706 : _GEN_14384; // @[sequencer-master.scala 647:41]
  wire  _GEN_16019 = io_op_bits_active_vfconv ? _GEN_15707 : _GEN_14385; // @[sequencer-master.scala 647:41]
  wire  _GEN_16020 = io_op_bits_active_vfconv ? _GEN_15708 : _GEN_14386; // @[sequencer-master.scala 647:41]
  wire  _GEN_16021 = io_op_bits_active_vfconv ? _GEN_15709 : _GEN_14387; // @[sequencer-master.scala 647:41]
  wire  _GEN_16022 = io_op_bits_active_vfconv ? _GEN_14870 : _GEN_14388; // @[sequencer-master.scala 647:41]
  wire  _GEN_16023 = io_op_bits_active_vfconv ? _GEN_14871 : _GEN_14389; // @[sequencer-master.scala 647:41]
  wire  _GEN_16024 = io_op_bits_active_vfconv ? _GEN_14872 : _GEN_14390; // @[sequencer-master.scala 647:41]
  wire  _GEN_16025 = io_op_bits_active_vfconv ? _GEN_14873 : _GEN_14391; // @[sequencer-master.scala 647:41]
  wire  _GEN_16026 = io_op_bits_active_vfconv ? _GEN_14874 : _GEN_14392; // @[sequencer-master.scala 647:41]
  wire  _GEN_16027 = io_op_bits_active_vfconv ? _GEN_14875 : _GEN_14393; // @[sequencer-master.scala 647:41]
  wire  _GEN_16028 = io_op_bits_active_vfconv ? _GEN_14876 : _GEN_14394; // @[sequencer-master.scala 647:41]
  wire  _GEN_16029 = io_op_bits_active_vfconv ? _GEN_14877 : _GEN_14395; // @[sequencer-master.scala 647:41]
  wire  _GEN_16038 = io_op_bits_active_vfconv ? _GEN_14886 : e_0_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16039 = io_op_bits_active_vfconv ? _GEN_14887 : e_1_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16040 = io_op_bits_active_vfconv ? _GEN_14888 : e_2_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16041 = io_op_bits_active_vfconv ? _GEN_14889 : e_3_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16042 = io_op_bits_active_vfconv ? _GEN_14890 : e_4_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16043 = io_op_bits_active_vfconv ? _GEN_14891 : e_5_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16044 = io_op_bits_active_vfconv ? _GEN_14892 : e_6_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire  _GEN_16045 = io_op_bits_active_vfconv ? _GEN_14893 : e_7_active_vfvu; // @[sequencer-master.scala 647:41 sequencer-master.scala 109:14]
  wire [9:0] _GEN_16046 = io_op_bits_active_vfconv ? _GEN_14894 : _GEN_14412; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16047 = io_op_bits_active_vfconv ? _GEN_14895 : _GEN_14413; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16048 = io_op_bits_active_vfconv ? _GEN_14896 : _GEN_14414; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16049 = io_op_bits_active_vfconv ? _GEN_14897 : _GEN_14415; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16050 = io_op_bits_active_vfconv ? _GEN_14898 : _GEN_14416; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16051 = io_op_bits_active_vfconv ? _GEN_14899 : _GEN_14417; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16052 = io_op_bits_active_vfconv ? _GEN_14900 : _GEN_14418; // @[sequencer-master.scala 647:41]
  wire [9:0] _GEN_16053 = io_op_bits_active_vfconv ? _GEN_14901 : _GEN_14419; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16054 = io_op_bits_active_vfconv ? _GEN_14942 : _GEN_14420; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16055 = io_op_bits_active_vfconv ? _GEN_14943 : _GEN_14421; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16056 = io_op_bits_active_vfconv ? _GEN_14944 : _GEN_14422; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16057 = io_op_bits_active_vfconv ? _GEN_14945 : _GEN_14423; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16058 = io_op_bits_active_vfconv ? _GEN_14946 : _GEN_14424; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16059 = io_op_bits_active_vfconv ? _GEN_14947 : _GEN_14425; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16060 = io_op_bits_active_vfconv ? _GEN_14948 : _GEN_14426; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16061 = io_op_bits_active_vfconv ? _GEN_14949 : _GEN_14427; // @[sequencer-master.scala 647:41]
  wire  _GEN_16062 = io_op_bits_active_vfconv ? _GEN_14958 : _GEN_14428; // @[sequencer-master.scala 647:41]
  wire  _GEN_16063 = io_op_bits_active_vfconv ? _GEN_14959 : _GEN_14429; // @[sequencer-master.scala 647:41]
  wire  _GEN_16064 = io_op_bits_active_vfconv ? _GEN_14960 : _GEN_14430; // @[sequencer-master.scala 647:41]
  wire  _GEN_16065 = io_op_bits_active_vfconv ? _GEN_14961 : _GEN_14431; // @[sequencer-master.scala 647:41]
  wire  _GEN_16066 = io_op_bits_active_vfconv ? _GEN_14962 : _GEN_14432; // @[sequencer-master.scala 647:41]
  wire  _GEN_16067 = io_op_bits_active_vfconv ? _GEN_14963 : _GEN_14433; // @[sequencer-master.scala 647:41]
  wire  _GEN_16068 = io_op_bits_active_vfconv ? _GEN_14964 : _GEN_14434; // @[sequencer-master.scala 647:41]
  wire  _GEN_16069 = io_op_bits_active_vfconv ? _GEN_14965 : _GEN_14435; // @[sequencer-master.scala 647:41]
  wire  _GEN_16070 = io_op_bits_active_vfconv ? _GEN_14966 : _GEN_14436; // @[sequencer-master.scala 647:41]
  wire  _GEN_16071 = io_op_bits_active_vfconv ? _GEN_14967 : _GEN_14437; // @[sequencer-master.scala 647:41]
  wire  _GEN_16072 = io_op_bits_active_vfconv ? _GEN_14968 : _GEN_14438; // @[sequencer-master.scala 647:41]
  wire  _GEN_16073 = io_op_bits_active_vfconv ? _GEN_14969 : _GEN_14439; // @[sequencer-master.scala 647:41]
  wire  _GEN_16074 = io_op_bits_active_vfconv ? _GEN_14970 : _GEN_14440; // @[sequencer-master.scala 647:41]
  wire  _GEN_16075 = io_op_bits_active_vfconv ? _GEN_14971 : _GEN_14441; // @[sequencer-master.scala 647:41]
  wire  _GEN_16076 = io_op_bits_active_vfconv ? _GEN_14972 : _GEN_14442; // @[sequencer-master.scala 647:41]
  wire  _GEN_16077 = io_op_bits_active_vfconv ? _GEN_14973 : _GEN_14443; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16078 = io_op_bits_active_vfconv ? _GEN_14974 : _GEN_14444; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16079 = io_op_bits_active_vfconv ? _GEN_14975 : _GEN_14445; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16080 = io_op_bits_active_vfconv ? _GEN_14976 : _GEN_14446; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16081 = io_op_bits_active_vfconv ? _GEN_14977 : _GEN_14447; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16082 = io_op_bits_active_vfconv ? _GEN_14978 : _GEN_14448; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16083 = io_op_bits_active_vfconv ? _GEN_14979 : _GEN_14449; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16084 = io_op_bits_active_vfconv ? _GEN_14980 : _GEN_14450; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16085 = io_op_bits_active_vfconv ? _GEN_14981 : _GEN_14451; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16086 = io_op_bits_active_vfconv ? _GEN_15174 : _GEN_14452; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16087 = io_op_bits_active_vfconv ? _GEN_15175 : _GEN_14453; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16088 = io_op_bits_active_vfconv ? _GEN_15176 : _GEN_14454; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16089 = io_op_bits_active_vfconv ? _GEN_15177 : _GEN_14455; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16090 = io_op_bits_active_vfconv ? _GEN_15178 : _GEN_14456; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16091 = io_op_bits_active_vfconv ? _GEN_15179 : _GEN_14457; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16092 = io_op_bits_active_vfconv ? _GEN_15180 : _GEN_14458; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16093 = io_op_bits_active_vfconv ? _GEN_15181 : _GEN_14459; // @[sequencer-master.scala 647:41]
  wire  _GEN_16094 = io_op_bits_active_vfconv ? _GEN_15190 : _GEN_14460; // @[sequencer-master.scala 647:41]
  wire  _GEN_16095 = io_op_bits_active_vfconv ? _GEN_15191 : _GEN_14461; // @[sequencer-master.scala 647:41]
  wire  _GEN_16096 = io_op_bits_active_vfconv ? _GEN_15192 : _GEN_14462; // @[sequencer-master.scala 647:41]
  wire  _GEN_16097 = io_op_bits_active_vfconv ? _GEN_15193 : _GEN_14463; // @[sequencer-master.scala 647:41]
  wire  _GEN_16098 = io_op_bits_active_vfconv ? _GEN_15194 : _GEN_14464; // @[sequencer-master.scala 647:41]
  wire  _GEN_16099 = io_op_bits_active_vfconv ? _GEN_15195 : _GEN_14465; // @[sequencer-master.scala 647:41]
  wire  _GEN_16100 = io_op_bits_active_vfconv ? _GEN_15196 : _GEN_14466; // @[sequencer-master.scala 647:41]
  wire  _GEN_16101 = io_op_bits_active_vfconv ? _GEN_15197 : _GEN_14467; // @[sequencer-master.scala 647:41]
  wire  _GEN_16102 = io_op_bits_active_vfconv ? _GEN_15198 : _GEN_14468; // @[sequencer-master.scala 647:41]
  wire  _GEN_16103 = io_op_bits_active_vfconv ? _GEN_15199 : _GEN_14469; // @[sequencer-master.scala 647:41]
  wire  _GEN_16104 = io_op_bits_active_vfconv ? _GEN_15200 : _GEN_14470; // @[sequencer-master.scala 647:41]
  wire  _GEN_16105 = io_op_bits_active_vfconv ? _GEN_15201 : _GEN_14471; // @[sequencer-master.scala 647:41]
  wire  _GEN_16106 = io_op_bits_active_vfconv ? _GEN_15202 : _GEN_14472; // @[sequencer-master.scala 647:41]
  wire  _GEN_16107 = io_op_bits_active_vfconv ? _GEN_15203 : _GEN_14473; // @[sequencer-master.scala 647:41]
  wire  _GEN_16108 = io_op_bits_active_vfconv ? _GEN_15204 : _GEN_14474; // @[sequencer-master.scala 647:41]
  wire  _GEN_16109 = io_op_bits_active_vfconv ? _GEN_15205 : _GEN_14475; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16110 = io_op_bits_active_vfconv ? _GEN_15206 : _GEN_14476; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16111 = io_op_bits_active_vfconv ? _GEN_15207 : _GEN_14477; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16112 = io_op_bits_active_vfconv ? _GEN_15208 : _GEN_14478; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16113 = io_op_bits_active_vfconv ? _GEN_15209 : _GEN_14479; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16114 = io_op_bits_active_vfconv ? _GEN_15210 : _GEN_14480; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16115 = io_op_bits_active_vfconv ? _GEN_15211 : _GEN_14481; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16116 = io_op_bits_active_vfconv ? _GEN_15212 : _GEN_14482; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16117 = io_op_bits_active_vfconv ? _GEN_15213 : _GEN_14483; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16118 = io_op_bits_active_vfconv ? _GEN_15214 : _GEN_14484; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16119 = io_op_bits_active_vfconv ? _GEN_15215 : _GEN_14485; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16120 = io_op_bits_active_vfconv ? _GEN_15216 : _GEN_14486; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16121 = io_op_bits_active_vfconv ? _GEN_15217 : _GEN_14487; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16122 = io_op_bits_active_vfconv ? _GEN_15218 : _GEN_14488; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16123 = io_op_bits_active_vfconv ? _GEN_15219 : _GEN_14489; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16124 = io_op_bits_active_vfconv ? _GEN_15220 : _GEN_14490; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16125 = io_op_bits_active_vfconv ? _GEN_15221 : _GEN_14491; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16126 = io_op_bits_active_vfconv ? _GEN_15222 : _GEN_14492; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16127 = io_op_bits_active_vfconv ? _GEN_15223 : _GEN_14493; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16128 = io_op_bits_active_vfconv ? _GEN_15224 : _GEN_14494; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16129 = io_op_bits_active_vfconv ? _GEN_15225 : _GEN_14495; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16130 = io_op_bits_active_vfconv ? _GEN_15226 : _GEN_14496; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16131 = io_op_bits_active_vfconv ? _GEN_15227 : _GEN_14497; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16132 = io_op_bits_active_vfconv ? _GEN_15228 : _GEN_14498; // @[sequencer-master.scala 647:41]
  wire [63:0] _GEN_16133 = io_op_bits_active_vfconv ? _GEN_15229 : _GEN_14499; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16134 = io_op_bits_active_vfconv ? _GEN_15406 : _GEN_14548; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16135 = io_op_bits_active_vfconv ? _GEN_15407 : _GEN_14549; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16136 = io_op_bits_active_vfconv ? _GEN_15408 : _GEN_14550; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16137 = io_op_bits_active_vfconv ? _GEN_15409 : _GEN_14551; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16138 = io_op_bits_active_vfconv ? _GEN_15410 : _GEN_14552; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16139 = io_op_bits_active_vfconv ? _GEN_15411 : _GEN_14553; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16140 = io_op_bits_active_vfconv ? _GEN_15412 : _GEN_14554; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16141 = io_op_bits_active_vfconv ? _GEN_15413 : _GEN_14555; // @[sequencer-master.scala 647:41]
  wire  _GEN_16142 = io_op_bits_active_vfconv ? _GEN_15422 : _GEN_14556; // @[sequencer-master.scala 647:41]
  wire  _GEN_16143 = io_op_bits_active_vfconv ? _GEN_15423 : _GEN_14557; // @[sequencer-master.scala 647:41]
  wire  _GEN_16144 = io_op_bits_active_vfconv ? _GEN_15424 : _GEN_14558; // @[sequencer-master.scala 647:41]
  wire  _GEN_16145 = io_op_bits_active_vfconv ? _GEN_15425 : _GEN_14559; // @[sequencer-master.scala 647:41]
  wire  _GEN_16146 = io_op_bits_active_vfconv ? _GEN_15426 : _GEN_14560; // @[sequencer-master.scala 647:41]
  wire  _GEN_16147 = io_op_bits_active_vfconv ? _GEN_15427 : _GEN_14561; // @[sequencer-master.scala 647:41]
  wire  _GEN_16148 = io_op_bits_active_vfconv ? _GEN_15428 : _GEN_14562; // @[sequencer-master.scala 647:41]
  wire  _GEN_16149 = io_op_bits_active_vfconv ? _GEN_15429 : _GEN_14563; // @[sequencer-master.scala 647:41]
  wire  _GEN_16150 = io_op_bits_active_vfconv ? _GEN_15430 : _GEN_14564; // @[sequencer-master.scala 647:41]
  wire  _GEN_16151 = io_op_bits_active_vfconv ? _GEN_15431 : _GEN_14565; // @[sequencer-master.scala 647:41]
  wire  _GEN_16152 = io_op_bits_active_vfconv ? _GEN_15432 : _GEN_14566; // @[sequencer-master.scala 647:41]
  wire  _GEN_16153 = io_op_bits_active_vfconv ? _GEN_15433 : _GEN_14567; // @[sequencer-master.scala 647:41]
  wire  _GEN_16154 = io_op_bits_active_vfconv ? _GEN_15434 : _GEN_14568; // @[sequencer-master.scala 647:41]
  wire  _GEN_16155 = io_op_bits_active_vfconv ? _GEN_15435 : _GEN_14569; // @[sequencer-master.scala 647:41]
  wire  _GEN_16156 = io_op_bits_active_vfconv ? _GEN_15436 : _GEN_14570; // @[sequencer-master.scala 647:41]
  wire  _GEN_16157 = io_op_bits_active_vfconv ? _GEN_15437 : _GEN_14571; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16158 = io_op_bits_active_vfconv ? _GEN_15438 : _GEN_14572; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16159 = io_op_bits_active_vfconv ? _GEN_15439 : _GEN_14573; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16160 = io_op_bits_active_vfconv ? _GEN_15440 : _GEN_14574; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16161 = io_op_bits_active_vfconv ? _GEN_15441 : _GEN_14575; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16162 = io_op_bits_active_vfconv ? _GEN_15442 : _GEN_14576; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16163 = io_op_bits_active_vfconv ? _GEN_15443 : _GEN_14577; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16164 = io_op_bits_active_vfconv ? _GEN_15444 : _GEN_14578; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16165 = io_op_bits_active_vfconv ? _GEN_15445 : _GEN_14579; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16166 = io_op_bits_active_vfconv ? _GEN_15446 : _GEN_14580; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16167 = io_op_bits_active_vfconv ? _GEN_15447 : _GEN_14581; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16168 = io_op_bits_active_vfconv ? _GEN_15448 : _GEN_14582; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16169 = io_op_bits_active_vfconv ? _GEN_15449 : _GEN_14583; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16170 = io_op_bits_active_vfconv ? _GEN_15450 : _GEN_14584; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16171 = io_op_bits_active_vfconv ? _GEN_15451 : _GEN_14585; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16172 = io_op_bits_active_vfconv ? _GEN_15452 : _GEN_14586; // @[sequencer-master.scala 647:41]
  wire [7:0] _GEN_16173 = io_op_bits_active_vfconv ? _GEN_15453 : _GEN_14587; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16174 = io_op_bits_active_vfconv ? _GEN_15710 : _GEN_14588; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16175 = io_op_bits_active_vfconv ? _GEN_15711 : _GEN_14589; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16176 = io_op_bits_active_vfconv ? _GEN_15712 : _GEN_14590; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16177 = io_op_bits_active_vfconv ? _GEN_15713 : _GEN_14591; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16178 = io_op_bits_active_vfconv ? _GEN_15714 : _GEN_14592; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16179 = io_op_bits_active_vfconv ? _GEN_15715 : _GEN_14593; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16180 = io_op_bits_active_vfconv ? _GEN_15716 : _GEN_14594; // @[sequencer-master.scala 647:41]
  wire [1:0] _GEN_16181 = io_op_bits_active_vfconv ? _GEN_15717 : _GEN_14595; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16182 = io_op_bits_active_vfconv ? _GEN_15742 : _GEN_14596; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16183 = io_op_bits_active_vfconv ? _GEN_15743 : _GEN_14597; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16184 = io_op_bits_active_vfconv ? _GEN_15744 : _GEN_14598; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16185 = io_op_bits_active_vfconv ? _GEN_15745 : _GEN_14599; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16186 = io_op_bits_active_vfconv ? _GEN_15746 : _GEN_14600; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16187 = io_op_bits_active_vfconv ? _GEN_15747 : _GEN_14601; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16188 = io_op_bits_active_vfconv ? _GEN_15748 : _GEN_14602; // @[sequencer-master.scala 647:41]
  wire [3:0] _GEN_16189 = io_op_bits_active_vfconv ? _GEN_15749 : _GEN_14603; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16190 = io_op_bits_active_vfconv ? _GEN_15758 : _GEN_14604; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16191 = io_op_bits_active_vfconv ? _GEN_15759 : _GEN_14605; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16192 = io_op_bits_active_vfconv ? _GEN_15760 : _GEN_14606; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16193 = io_op_bits_active_vfconv ? _GEN_15761 : _GEN_14607; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16194 = io_op_bits_active_vfconv ? _GEN_15762 : _GEN_14608; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16195 = io_op_bits_active_vfconv ? _GEN_15763 : _GEN_14609; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16196 = io_op_bits_active_vfconv ? _GEN_15764 : _GEN_14610; // @[sequencer-master.scala 647:41]
  wire [2:0] _GEN_16197 = io_op_bits_active_vfconv ? _GEN_15765 : _GEN_14611; // @[sequencer-master.scala 647:41]
  wire  _GEN_16198 = io_op_bits_active_vfconv | _GEN_14612; // @[sequencer-master.scala 647:41 sequencer-master.scala 265:41]
  wire [2:0] _GEN_16199 = io_op_bits_active_vfconv ? _T_1645 : _GEN_14613; // @[sequencer-master.scala 647:41 sequencer-master.scala 265:66]
  wire  _GEN_16200 = _GEN_32729 | _GEN_15766; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16201 = _GEN_32730 | _GEN_15767; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16202 = _GEN_32731 | _GEN_15768; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16203 = _GEN_32732 | _GEN_15769; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16204 = _GEN_32733 | _GEN_15770; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16205 = _GEN_32734 | _GEN_15771; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16206 = _GEN_32735 | _GEN_15772; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16207 = _GEN_32736 | _GEN_15773; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_16216 = 3'h0 == tail ? 1'h0 : _GEN_15782; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16217 = 3'h1 == tail ? 1'h0 : _GEN_15783; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16218 = 3'h2 == tail ? 1'h0 : _GEN_15784; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16219 = 3'h3 == tail ? 1'h0 : _GEN_15785; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16220 = 3'h4 == tail ? 1'h0 : _GEN_15786; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16221 = 3'h5 == tail ? 1'h0 : _GEN_15787; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16222 = 3'h6 == tail ? 1'h0 : _GEN_15788; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16223 = 3'h7 == tail ? 1'h0 : _GEN_15789; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_16224 = 3'h0 == tail ? 1'h0 : _GEN_15790; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16225 = 3'h1 == tail ? 1'h0 : _GEN_15791; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16226 = 3'h2 == tail ? 1'h0 : _GEN_15792; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16227 = 3'h3 == tail ? 1'h0 : _GEN_15793; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16228 = 3'h4 == tail ? 1'h0 : _GEN_15794; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16229 = 3'h5 == tail ? 1'h0 : _GEN_15795; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16230 = 3'h6 == tail ? 1'h0 : _GEN_15796; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16231 = 3'h7 == tail ? 1'h0 : _GEN_15797; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_16232 = 3'h0 == tail ? 1'h0 : _GEN_15798; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16233 = 3'h1 == tail ? 1'h0 : _GEN_15799; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16234 = 3'h2 == tail ? 1'h0 : _GEN_15800; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16235 = 3'h3 == tail ? 1'h0 : _GEN_15801; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16236 = 3'h4 == tail ? 1'h0 : _GEN_15802; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16237 = 3'h5 == tail ? 1'h0 : _GEN_15803; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16238 = 3'h6 == tail ? 1'h0 : _GEN_15804; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16239 = 3'h7 == tail ? 1'h0 : _GEN_15805; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_16240 = 3'h0 == tail ? 1'h0 : _GEN_15806; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16241 = 3'h1 == tail ? 1'h0 : _GEN_15807; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16242 = 3'h2 == tail ? 1'h0 : _GEN_15808; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16243 = 3'h3 == tail ? 1'h0 : _GEN_15809; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16244 = 3'h4 == tail ? 1'h0 : _GEN_15810; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16245 = 3'h5 == tail ? 1'h0 : _GEN_15811; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16246 = 3'h6 == tail ? 1'h0 : _GEN_15812; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16247 = 3'h7 == tail ? 1'h0 : _GEN_15813; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_16248 = 3'h0 == tail ? 1'h0 : _GEN_15814; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16249 = 3'h1 == tail ? 1'h0 : _GEN_15815; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16250 = 3'h2 == tail ? 1'h0 : _GEN_15816; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16251 = 3'h3 == tail ? 1'h0 : _GEN_15817; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16252 = 3'h4 == tail ? 1'h0 : _GEN_15818; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16253 = 3'h5 == tail ? 1'h0 : _GEN_15819; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16254 = 3'h6 == tail ? 1'h0 : _GEN_15820; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16255 = 3'h7 == tail ? 1'h0 : _GEN_15821; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_16256 = _GEN_32729 | _GEN_15822; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16257 = _GEN_32730 | _GEN_15823; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16258 = _GEN_32731 | _GEN_15824; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16259 = _GEN_32732 | _GEN_15825; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16260 = _GEN_32733 | _GEN_15826; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16261 = _GEN_32734 | _GEN_15827; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16262 = _GEN_32735 | _GEN_15828; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16263 = _GEN_32736 | _GEN_15829; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_16264 = 3'h0 == tail ? 1'h0 : _GEN_15830; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16265 = 3'h1 == tail ? 1'h0 : _GEN_15831; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16266 = 3'h2 == tail ? 1'h0 : _GEN_15832; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16267 = 3'h3 == tail ? 1'h0 : _GEN_15833; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16268 = 3'h4 == tail ? 1'h0 : _GEN_15834; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16269 = 3'h5 == tail ? 1'h0 : _GEN_15835; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16270 = 3'h6 == tail ? 1'h0 : _GEN_15836; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16271 = 3'h7 == tail ? 1'h0 : _GEN_15837; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16272 = 3'h0 == tail ? 1'h0 : _GEN_15838; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16273 = 3'h1 == tail ? 1'h0 : _GEN_15839; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16274 = 3'h2 == tail ? 1'h0 : _GEN_15840; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16275 = 3'h3 == tail ? 1'h0 : _GEN_15841; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16276 = 3'h4 == tail ? 1'h0 : _GEN_15842; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16277 = 3'h5 == tail ? 1'h0 : _GEN_15843; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16278 = 3'h6 == tail ? 1'h0 : _GEN_15844; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16279 = 3'h7 == tail ? 1'h0 : _GEN_15845; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16280 = 3'h0 == tail ? 1'h0 : _GEN_15846; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16281 = 3'h1 == tail ? 1'h0 : _GEN_15847; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16282 = 3'h2 == tail ? 1'h0 : _GEN_15848; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16283 = 3'h3 == tail ? 1'h0 : _GEN_15849; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16284 = 3'h4 == tail ? 1'h0 : _GEN_15850; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16285 = 3'h5 == tail ? 1'h0 : _GEN_15851; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16286 = 3'h6 == tail ? 1'h0 : _GEN_15852; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16287 = 3'h7 == tail ? 1'h0 : _GEN_15853; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16288 = 3'h0 == tail ? 1'h0 : _GEN_15854; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16289 = 3'h1 == tail ? 1'h0 : _GEN_15855; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16290 = 3'h2 == tail ? 1'h0 : _GEN_15856; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16291 = 3'h3 == tail ? 1'h0 : _GEN_15857; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16292 = 3'h4 == tail ? 1'h0 : _GEN_15858; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16293 = 3'h5 == tail ? 1'h0 : _GEN_15859; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16294 = 3'h6 == tail ? 1'h0 : _GEN_15860; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16295 = 3'h7 == tail ? 1'h0 : _GEN_15861; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16296 = 3'h0 == tail ? 1'h0 : _GEN_15862; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16297 = 3'h1 == tail ? 1'h0 : _GEN_15863; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16298 = 3'h2 == tail ? 1'h0 : _GEN_15864; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16299 = 3'h3 == tail ? 1'h0 : _GEN_15865; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16300 = 3'h4 == tail ? 1'h0 : _GEN_15866; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16301 = 3'h5 == tail ? 1'h0 : _GEN_15867; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16302 = 3'h6 == tail ? 1'h0 : _GEN_15868; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16303 = 3'h7 == tail ? 1'h0 : _GEN_15869; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16304 = 3'h0 == tail ? 1'h0 : _GEN_15870; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16305 = 3'h1 == tail ? 1'h0 : _GEN_15871; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16306 = 3'h2 == tail ? 1'h0 : _GEN_15872; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16307 = 3'h3 == tail ? 1'h0 : _GEN_15873; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16308 = 3'h4 == tail ? 1'h0 : _GEN_15874; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16309 = 3'h5 == tail ? 1'h0 : _GEN_15875; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16310 = 3'h6 == tail ? 1'h0 : _GEN_15876; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16311 = 3'h7 == tail ? 1'h0 : _GEN_15877; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16312 = 3'h0 == tail ? 1'h0 : _GEN_15878; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16313 = 3'h1 == tail ? 1'h0 : _GEN_15879; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16314 = 3'h2 == tail ? 1'h0 : _GEN_15880; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16315 = 3'h3 == tail ? 1'h0 : _GEN_15881; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16316 = 3'h4 == tail ? 1'h0 : _GEN_15882; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16317 = 3'h5 == tail ? 1'h0 : _GEN_15883; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16318 = 3'h6 == tail ? 1'h0 : _GEN_15884; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16319 = 3'h7 == tail ? 1'h0 : _GEN_15885; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16320 = 3'h0 == tail ? 1'h0 : _GEN_15886; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16321 = 3'h1 == tail ? 1'h0 : _GEN_15887; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16322 = 3'h2 == tail ? 1'h0 : _GEN_15888; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16323 = 3'h3 == tail ? 1'h0 : _GEN_15889; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16324 = 3'h4 == tail ? 1'h0 : _GEN_15890; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16325 = 3'h5 == tail ? 1'h0 : _GEN_15891; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16326 = 3'h6 == tail ? 1'h0 : _GEN_15892; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16327 = 3'h7 == tail ? 1'h0 : _GEN_15893; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16328 = 3'h0 == tail ? 1'h0 : _GEN_15894; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16329 = 3'h1 == tail ? 1'h0 : _GEN_15895; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16330 = 3'h2 == tail ? 1'h0 : _GEN_15896; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16331 = 3'h3 == tail ? 1'h0 : _GEN_15897; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16332 = 3'h4 == tail ? 1'h0 : _GEN_15898; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16333 = 3'h5 == tail ? 1'h0 : _GEN_15899; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16334 = 3'h6 == tail ? 1'h0 : _GEN_15900; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16335 = 3'h7 == tail ? 1'h0 : _GEN_15901; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16336 = 3'h0 == tail ? 1'h0 : _GEN_15902; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16337 = 3'h1 == tail ? 1'h0 : _GEN_15903; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16338 = 3'h2 == tail ? 1'h0 : _GEN_15904; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16339 = 3'h3 == tail ? 1'h0 : _GEN_15905; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16340 = 3'h4 == tail ? 1'h0 : _GEN_15906; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16341 = 3'h5 == tail ? 1'h0 : _GEN_15907; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16342 = 3'h6 == tail ? 1'h0 : _GEN_15908; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16343 = 3'h7 == tail ? 1'h0 : _GEN_15909; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16344 = 3'h0 == tail ? 1'h0 : _GEN_15910; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16345 = 3'h1 == tail ? 1'h0 : _GEN_15911; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16346 = 3'h2 == tail ? 1'h0 : _GEN_15912; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16347 = 3'h3 == tail ? 1'h0 : _GEN_15913; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16348 = 3'h4 == tail ? 1'h0 : _GEN_15914; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16349 = 3'h5 == tail ? 1'h0 : _GEN_15915; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16350 = 3'h6 == tail ? 1'h0 : _GEN_15916; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16351 = 3'h7 == tail ? 1'h0 : _GEN_15917; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16352 = 3'h0 == tail ? 1'h0 : _GEN_15918; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16353 = 3'h1 == tail ? 1'h0 : _GEN_15919; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16354 = 3'h2 == tail ? 1'h0 : _GEN_15920; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16355 = 3'h3 == tail ? 1'h0 : _GEN_15921; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16356 = 3'h4 == tail ? 1'h0 : _GEN_15922; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16357 = 3'h5 == tail ? 1'h0 : _GEN_15923; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16358 = 3'h6 == tail ? 1'h0 : _GEN_15924; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16359 = 3'h7 == tail ? 1'h0 : _GEN_15925; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16360 = 3'h0 == tail ? 1'h0 : _GEN_15926; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16361 = 3'h1 == tail ? 1'h0 : _GEN_15927; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16362 = 3'h2 == tail ? 1'h0 : _GEN_15928; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16363 = 3'h3 == tail ? 1'h0 : _GEN_15929; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16364 = 3'h4 == tail ? 1'h0 : _GEN_15930; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16365 = 3'h5 == tail ? 1'h0 : _GEN_15931; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16366 = 3'h6 == tail ? 1'h0 : _GEN_15932; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16367 = 3'h7 == tail ? 1'h0 : _GEN_15933; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16368 = 3'h0 == tail ? 1'h0 : _GEN_15934; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16369 = 3'h1 == tail ? 1'h0 : _GEN_15935; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16370 = 3'h2 == tail ? 1'h0 : _GEN_15936; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16371 = 3'h3 == tail ? 1'h0 : _GEN_15937; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16372 = 3'h4 == tail ? 1'h0 : _GEN_15938; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16373 = 3'h5 == tail ? 1'h0 : _GEN_15939; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16374 = 3'h6 == tail ? 1'h0 : _GEN_15940; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16375 = 3'h7 == tail ? 1'h0 : _GEN_15941; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16376 = 3'h0 == tail ? 1'h0 : _GEN_15942; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16377 = 3'h1 == tail ? 1'h0 : _GEN_15943; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16378 = 3'h2 == tail ? 1'h0 : _GEN_15944; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16379 = 3'h3 == tail ? 1'h0 : _GEN_15945; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16380 = 3'h4 == tail ? 1'h0 : _GEN_15946; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16381 = 3'h5 == tail ? 1'h0 : _GEN_15947; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16382 = 3'h6 == tail ? 1'h0 : _GEN_15948; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16383 = 3'h7 == tail ? 1'h0 : _GEN_15949; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16384 = 3'h0 == tail ? 1'h0 : _GEN_15950; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16385 = 3'h1 == tail ? 1'h0 : _GEN_15951; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16386 = 3'h2 == tail ? 1'h0 : _GEN_15952; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16387 = 3'h3 == tail ? 1'h0 : _GEN_15953; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16388 = 3'h4 == tail ? 1'h0 : _GEN_15954; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16389 = 3'h5 == tail ? 1'h0 : _GEN_15955; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16390 = 3'h6 == tail ? 1'h0 : _GEN_15956; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16391 = 3'h7 == tail ? 1'h0 : _GEN_15957; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16392 = 3'h0 == tail ? 1'h0 : _GEN_15958; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16393 = 3'h1 == tail ? 1'h0 : _GEN_15959; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16394 = 3'h2 == tail ? 1'h0 : _GEN_15960; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16395 = 3'h3 == tail ? 1'h0 : _GEN_15961; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16396 = 3'h4 == tail ? 1'h0 : _GEN_15962; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16397 = 3'h5 == tail ? 1'h0 : _GEN_15963; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16398 = 3'h6 == tail ? 1'h0 : _GEN_15964; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16399 = 3'h7 == tail ? 1'h0 : _GEN_15965; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16400 = 3'h0 == tail ? 1'h0 : _GEN_15966; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16401 = 3'h1 == tail ? 1'h0 : _GEN_15967; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16402 = 3'h2 == tail ? 1'h0 : _GEN_15968; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16403 = 3'h3 == tail ? 1'h0 : _GEN_15969; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16404 = 3'h4 == tail ? 1'h0 : _GEN_15970; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16405 = 3'h5 == tail ? 1'h0 : _GEN_15971; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16406 = 3'h6 == tail ? 1'h0 : _GEN_15972; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16407 = 3'h7 == tail ? 1'h0 : _GEN_15973; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16408 = 3'h0 == tail ? 1'h0 : _GEN_15974; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16409 = 3'h1 == tail ? 1'h0 : _GEN_15975; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16410 = 3'h2 == tail ? 1'h0 : _GEN_15976; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16411 = 3'h3 == tail ? 1'h0 : _GEN_15977; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16412 = 3'h4 == tail ? 1'h0 : _GEN_15978; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16413 = 3'h5 == tail ? 1'h0 : _GEN_15979; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16414 = 3'h6 == tail ? 1'h0 : _GEN_15980; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16415 = 3'h7 == tail ? 1'h0 : _GEN_15981; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16416 = 3'h0 == tail ? 1'h0 : _GEN_15982; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16417 = 3'h1 == tail ? 1'h0 : _GEN_15983; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16418 = 3'h2 == tail ? 1'h0 : _GEN_15984; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16419 = 3'h3 == tail ? 1'h0 : _GEN_15985; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16420 = 3'h4 == tail ? 1'h0 : _GEN_15986; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16421 = 3'h5 == tail ? 1'h0 : _GEN_15987; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16422 = 3'h6 == tail ? 1'h0 : _GEN_15988; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16423 = 3'h7 == tail ? 1'h0 : _GEN_15989; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16424 = 3'h0 == tail ? 1'h0 : _GEN_15990; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16425 = 3'h1 == tail ? 1'h0 : _GEN_15991; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16426 = 3'h2 == tail ? 1'h0 : _GEN_15992; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16427 = 3'h3 == tail ? 1'h0 : _GEN_15993; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16428 = 3'h4 == tail ? 1'h0 : _GEN_15994; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16429 = 3'h5 == tail ? 1'h0 : _GEN_15995; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16430 = 3'h6 == tail ? 1'h0 : _GEN_15996; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16431 = 3'h7 == tail ? 1'h0 : _GEN_15997; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16432 = 3'h0 == tail ? 1'h0 : _GEN_15998; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16433 = 3'h1 == tail ? 1'h0 : _GEN_15999; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16434 = 3'h2 == tail ? 1'h0 : _GEN_16000; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16435 = 3'h3 == tail ? 1'h0 : _GEN_16001; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16436 = 3'h4 == tail ? 1'h0 : _GEN_16002; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16437 = 3'h5 == tail ? 1'h0 : _GEN_16003; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16438 = 3'h6 == tail ? 1'h0 : _GEN_16004; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16439 = 3'h7 == tail ? 1'h0 : _GEN_16005; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_16440 = 3'h0 == tail ? 1'h0 : _GEN_16006; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16441 = 3'h1 == tail ? 1'h0 : _GEN_16007; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16442 = 3'h2 == tail ? 1'h0 : _GEN_16008; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16443 = 3'h3 == tail ? 1'h0 : _GEN_16009; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16444 = 3'h4 == tail ? 1'h0 : _GEN_16010; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16445 = 3'h5 == tail ? 1'h0 : _GEN_16011; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16446 = 3'h6 == tail ? 1'h0 : _GEN_16012; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16447 = 3'h7 == tail ? 1'h0 : _GEN_16013; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_16448 = 3'h0 == tail ? 1'h0 : _GEN_16014; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16449 = 3'h1 == tail ? 1'h0 : _GEN_16015; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16450 = 3'h2 == tail ? 1'h0 : _GEN_16016; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16451 = 3'h3 == tail ? 1'h0 : _GEN_16017; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16452 = 3'h4 == tail ? 1'h0 : _GEN_16018; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16453 = 3'h5 == tail ? 1'h0 : _GEN_16019; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16454 = 3'h6 == tail ? 1'h0 : _GEN_16020; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16455 = 3'h7 == tail ? 1'h0 : _GEN_16021; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_16456 = 3'h0 == tail ? 1'h0 : _GEN_16022; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16457 = 3'h1 == tail ? 1'h0 : _GEN_16023; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16458 = 3'h2 == tail ? 1'h0 : _GEN_16024; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16459 = 3'h3 == tail ? 1'h0 : _GEN_16025; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16460 = 3'h4 == tail ? 1'h0 : _GEN_16026; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16461 = 3'h5 == tail ? 1'h0 : _GEN_16027; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16462 = 3'h6 == tail ? 1'h0 : _GEN_16028; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16463 = 3'h7 == tail ? 1'h0 : _GEN_16029; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_16472 = _GEN_32729 | _GEN_12514; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16473 = _GEN_32730 | _GEN_12515; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16474 = _GEN_32731 | _GEN_12516; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16475 = _GEN_32732 | _GEN_12517; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16476 = _GEN_32733 | _GEN_12518; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16477 = _GEN_32734 | _GEN_12519; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16478 = _GEN_32735 | _GEN_12520; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_16479 = _GEN_32736 | _GEN_12521; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_16480 = 3'h0 == tail ? _e_tail_fn_union_2 : _GEN_16046; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16481 = 3'h1 == tail ? _e_tail_fn_union_2 : _GEN_16047; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16482 = 3'h2 == tail ? _e_tail_fn_union_2 : _GEN_16048; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16483 = 3'h3 == tail ? _e_tail_fn_union_2 : _GEN_16049; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16484 = 3'h4 == tail ? _e_tail_fn_union_2 : _GEN_16050; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16485 = 3'h5 == tail ? _e_tail_fn_union_2 : _GEN_16051; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16486 = 3'h6 == tail ? _e_tail_fn_union_2 : _GEN_16052; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_16487 = 3'h7 == tail ? _e_tail_fn_union_2 : _GEN_16053; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_16488 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_16054; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16489 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_16055; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16490 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_16056; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16491 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_16057; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16492 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_16058; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16493 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_16059; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16494 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_16060; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_16495 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_16061; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16496 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_16216; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16497 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_16217; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16498 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_16218; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16499 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_16219; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16500 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_16220; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16501 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_16221; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16502 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_16222; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16503 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_16223; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16504 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_16062; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16505 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_16063; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16506 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_16064; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16507 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_16065; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16508 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_16066; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16509 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_16067; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16510 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_16068; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16511 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_16069; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16512 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_16070; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16513 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_16071; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16514 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_16072; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16515 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_16073; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16516 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_16074; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16517 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_16075; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16518 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_16076; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_16519 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_16077; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_16520 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_16078; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16521 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_16079; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16522 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_16080; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16523 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_16081; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16524 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_16082; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16525 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_16083; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16526 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_16084; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_16527 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_16085; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_16528 = io_op_bits_base_vp_valid ? _GEN_16488 : _GEN_16054; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16529 = io_op_bits_base_vp_valid ? _GEN_16489 : _GEN_16055; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16530 = io_op_bits_base_vp_valid ? _GEN_16490 : _GEN_16056; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16531 = io_op_bits_base_vp_valid ? _GEN_16491 : _GEN_16057; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16532 = io_op_bits_base_vp_valid ? _GEN_16492 : _GEN_16058; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16533 = io_op_bits_base_vp_valid ? _GEN_16493 : _GEN_16059; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16534 = io_op_bits_base_vp_valid ? _GEN_16494 : _GEN_16060; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_16535 = io_op_bits_base_vp_valid ? _GEN_16495 : _GEN_16061; // @[sequencer-master.scala 320:41]
  wire  _GEN_16536 = io_op_bits_base_vp_valid ? _GEN_16496 : _GEN_16216; // @[sequencer-master.scala 320:41]
  wire  _GEN_16537 = io_op_bits_base_vp_valid ? _GEN_16497 : _GEN_16217; // @[sequencer-master.scala 320:41]
  wire  _GEN_16538 = io_op_bits_base_vp_valid ? _GEN_16498 : _GEN_16218; // @[sequencer-master.scala 320:41]
  wire  _GEN_16539 = io_op_bits_base_vp_valid ? _GEN_16499 : _GEN_16219; // @[sequencer-master.scala 320:41]
  wire  _GEN_16540 = io_op_bits_base_vp_valid ? _GEN_16500 : _GEN_16220; // @[sequencer-master.scala 320:41]
  wire  _GEN_16541 = io_op_bits_base_vp_valid ? _GEN_16501 : _GEN_16221; // @[sequencer-master.scala 320:41]
  wire  _GEN_16542 = io_op_bits_base_vp_valid ? _GEN_16502 : _GEN_16222; // @[sequencer-master.scala 320:41]
  wire  _GEN_16543 = io_op_bits_base_vp_valid ? _GEN_16503 : _GEN_16223; // @[sequencer-master.scala 320:41]
  wire  _GEN_16544 = io_op_bits_base_vp_valid ? _GEN_16504 : _GEN_16062; // @[sequencer-master.scala 320:41]
  wire  _GEN_16545 = io_op_bits_base_vp_valid ? _GEN_16505 : _GEN_16063; // @[sequencer-master.scala 320:41]
  wire  _GEN_16546 = io_op_bits_base_vp_valid ? _GEN_16506 : _GEN_16064; // @[sequencer-master.scala 320:41]
  wire  _GEN_16547 = io_op_bits_base_vp_valid ? _GEN_16507 : _GEN_16065; // @[sequencer-master.scala 320:41]
  wire  _GEN_16548 = io_op_bits_base_vp_valid ? _GEN_16508 : _GEN_16066; // @[sequencer-master.scala 320:41]
  wire  _GEN_16549 = io_op_bits_base_vp_valid ? _GEN_16509 : _GEN_16067; // @[sequencer-master.scala 320:41]
  wire  _GEN_16550 = io_op_bits_base_vp_valid ? _GEN_16510 : _GEN_16068; // @[sequencer-master.scala 320:41]
  wire  _GEN_16551 = io_op_bits_base_vp_valid ? _GEN_16511 : _GEN_16069; // @[sequencer-master.scala 320:41]
  wire  _GEN_16552 = io_op_bits_base_vp_valid ? _GEN_16512 : _GEN_16070; // @[sequencer-master.scala 320:41]
  wire  _GEN_16553 = io_op_bits_base_vp_valid ? _GEN_16513 : _GEN_16071; // @[sequencer-master.scala 320:41]
  wire  _GEN_16554 = io_op_bits_base_vp_valid ? _GEN_16514 : _GEN_16072; // @[sequencer-master.scala 320:41]
  wire  _GEN_16555 = io_op_bits_base_vp_valid ? _GEN_16515 : _GEN_16073; // @[sequencer-master.scala 320:41]
  wire  _GEN_16556 = io_op_bits_base_vp_valid ? _GEN_16516 : _GEN_16074; // @[sequencer-master.scala 320:41]
  wire  _GEN_16557 = io_op_bits_base_vp_valid ? _GEN_16517 : _GEN_16075; // @[sequencer-master.scala 320:41]
  wire  _GEN_16558 = io_op_bits_base_vp_valid ? _GEN_16518 : _GEN_16076; // @[sequencer-master.scala 320:41]
  wire  _GEN_16559 = io_op_bits_base_vp_valid ? _GEN_16519 : _GEN_16077; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16560 = io_op_bits_base_vp_valid ? _GEN_16520 : _GEN_16078; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16561 = io_op_bits_base_vp_valid ? _GEN_16521 : _GEN_16079; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16562 = io_op_bits_base_vp_valid ? _GEN_16522 : _GEN_16080; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16563 = io_op_bits_base_vp_valid ? _GEN_16523 : _GEN_16081; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16564 = io_op_bits_base_vp_valid ? _GEN_16524 : _GEN_16082; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16565 = io_op_bits_base_vp_valid ? _GEN_16525 : _GEN_16083; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16566 = io_op_bits_base_vp_valid ? _GEN_16526 : _GEN_16084; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_16567 = io_op_bits_base_vp_valid ? _GEN_16527 : _GEN_16085; // @[sequencer-master.scala 320:41]
  wire  _GEN_16568 = _GEN_32729 | _GEN_16264; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16569 = _GEN_32730 | _GEN_16265; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16570 = _GEN_32731 | _GEN_16266; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16571 = _GEN_32732 | _GEN_16267; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16572 = _GEN_32733 | _GEN_16268; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16573 = _GEN_32734 | _GEN_16269; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16574 = _GEN_32735 | _GEN_16270; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16575 = _GEN_32736 | _GEN_16271; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16576 = _T_26 ? _GEN_16568 : _GEN_16264; // @[sequencer-master.scala 154:24]
  wire  _GEN_16577 = _T_26 ? _GEN_16569 : _GEN_16265; // @[sequencer-master.scala 154:24]
  wire  _GEN_16578 = _T_26 ? _GEN_16570 : _GEN_16266; // @[sequencer-master.scala 154:24]
  wire  _GEN_16579 = _T_26 ? _GEN_16571 : _GEN_16267; // @[sequencer-master.scala 154:24]
  wire  _GEN_16580 = _T_26 ? _GEN_16572 : _GEN_16268; // @[sequencer-master.scala 154:24]
  wire  _GEN_16581 = _T_26 ? _GEN_16573 : _GEN_16269; // @[sequencer-master.scala 154:24]
  wire  _GEN_16582 = _T_26 ? _GEN_16574 : _GEN_16270; // @[sequencer-master.scala 154:24]
  wire  _GEN_16583 = _T_26 ? _GEN_16575 : _GEN_16271; // @[sequencer-master.scala 154:24]
  wire  _GEN_16584 = _GEN_32729 | _GEN_16288; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16585 = _GEN_32730 | _GEN_16289; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16586 = _GEN_32731 | _GEN_16290; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16587 = _GEN_32732 | _GEN_16291; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16588 = _GEN_32733 | _GEN_16292; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16589 = _GEN_32734 | _GEN_16293; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16590 = _GEN_32735 | _GEN_16294; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16591 = _GEN_32736 | _GEN_16295; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16592 = _T_48 ? _GEN_16584 : _GEN_16288; // @[sequencer-master.scala 154:24]
  wire  _GEN_16593 = _T_48 ? _GEN_16585 : _GEN_16289; // @[sequencer-master.scala 154:24]
  wire  _GEN_16594 = _T_48 ? _GEN_16586 : _GEN_16290; // @[sequencer-master.scala 154:24]
  wire  _GEN_16595 = _T_48 ? _GEN_16587 : _GEN_16291; // @[sequencer-master.scala 154:24]
  wire  _GEN_16596 = _T_48 ? _GEN_16588 : _GEN_16292; // @[sequencer-master.scala 154:24]
  wire  _GEN_16597 = _T_48 ? _GEN_16589 : _GEN_16293; // @[sequencer-master.scala 154:24]
  wire  _GEN_16598 = _T_48 ? _GEN_16590 : _GEN_16294; // @[sequencer-master.scala 154:24]
  wire  _GEN_16599 = _T_48 ? _GEN_16591 : _GEN_16295; // @[sequencer-master.scala 154:24]
  wire  _GEN_16600 = _GEN_32729 | _GEN_16312; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16601 = _GEN_32730 | _GEN_16313; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16602 = _GEN_32731 | _GEN_16314; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16603 = _GEN_32732 | _GEN_16315; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16604 = _GEN_32733 | _GEN_16316; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16605 = _GEN_32734 | _GEN_16317; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16606 = _GEN_32735 | _GEN_16318; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16607 = _GEN_32736 | _GEN_16319; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16608 = _T_70 ? _GEN_16600 : _GEN_16312; // @[sequencer-master.scala 154:24]
  wire  _GEN_16609 = _T_70 ? _GEN_16601 : _GEN_16313; // @[sequencer-master.scala 154:24]
  wire  _GEN_16610 = _T_70 ? _GEN_16602 : _GEN_16314; // @[sequencer-master.scala 154:24]
  wire  _GEN_16611 = _T_70 ? _GEN_16603 : _GEN_16315; // @[sequencer-master.scala 154:24]
  wire  _GEN_16612 = _T_70 ? _GEN_16604 : _GEN_16316; // @[sequencer-master.scala 154:24]
  wire  _GEN_16613 = _T_70 ? _GEN_16605 : _GEN_16317; // @[sequencer-master.scala 154:24]
  wire  _GEN_16614 = _T_70 ? _GEN_16606 : _GEN_16318; // @[sequencer-master.scala 154:24]
  wire  _GEN_16615 = _T_70 ? _GEN_16607 : _GEN_16319; // @[sequencer-master.scala 154:24]
  wire  _GEN_16616 = _GEN_32729 | _GEN_16336; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16617 = _GEN_32730 | _GEN_16337; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16618 = _GEN_32731 | _GEN_16338; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16619 = _GEN_32732 | _GEN_16339; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16620 = _GEN_32733 | _GEN_16340; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16621 = _GEN_32734 | _GEN_16341; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16622 = _GEN_32735 | _GEN_16342; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16623 = _GEN_32736 | _GEN_16343; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16624 = _T_92 ? _GEN_16616 : _GEN_16336; // @[sequencer-master.scala 154:24]
  wire  _GEN_16625 = _T_92 ? _GEN_16617 : _GEN_16337; // @[sequencer-master.scala 154:24]
  wire  _GEN_16626 = _T_92 ? _GEN_16618 : _GEN_16338; // @[sequencer-master.scala 154:24]
  wire  _GEN_16627 = _T_92 ? _GEN_16619 : _GEN_16339; // @[sequencer-master.scala 154:24]
  wire  _GEN_16628 = _T_92 ? _GEN_16620 : _GEN_16340; // @[sequencer-master.scala 154:24]
  wire  _GEN_16629 = _T_92 ? _GEN_16621 : _GEN_16341; // @[sequencer-master.scala 154:24]
  wire  _GEN_16630 = _T_92 ? _GEN_16622 : _GEN_16342; // @[sequencer-master.scala 154:24]
  wire  _GEN_16631 = _T_92 ? _GEN_16623 : _GEN_16343; // @[sequencer-master.scala 154:24]
  wire  _GEN_16632 = _GEN_32729 | _GEN_16360; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16633 = _GEN_32730 | _GEN_16361; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16634 = _GEN_32731 | _GEN_16362; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16635 = _GEN_32732 | _GEN_16363; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16636 = _GEN_32733 | _GEN_16364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16637 = _GEN_32734 | _GEN_16365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16638 = _GEN_32735 | _GEN_16366; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16639 = _GEN_32736 | _GEN_16367; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16640 = _T_114 ? _GEN_16632 : _GEN_16360; // @[sequencer-master.scala 154:24]
  wire  _GEN_16641 = _T_114 ? _GEN_16633 : _GEN_16361; // @[sequencer-master.scala 154:24]
  wire  _GEN_16642 = _T_114 ? _GEN_16634 : _GEN_16362; // @[sequencer-master.scala 154:24]
  wire  _GEN_16643 = _T_114 ? _GEN_16635 : _GEN_16363; // @[sequencer-master.scala 154:24]
  wire  _GEN_16644 = _T_114 ? _GEN_16636 : _GEN_16364; // @[sequencer-master.scala 154:24]
  wire  _GEN_16645 = _T_114 ? _GEN_16637 : _GEN_16365; // @[sequencer-master.scala 154:24]
  wire  _GEN_16646 = _T_114 ? _GEN_16638 : _GEN_16366; // @[sequencer-master.scala 154:24]
  wire  _GEN_16647 = _T_114 ? _GEN_16639 : _GEN_16367; // @[sequencer-master.scala 154:24]
  wire  _GEN_16648 = _GEN_32729 | _GEN_16384; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16649 = _GEN_32730 | _GEN_16385; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16650 = _GEN_32731 | _GEN_16386; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16651 = _GEN_32732 | _GEN_16387; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16652 = _GEN_32733 | _GEN_16388; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16653 = _GEN_32734 | _GEN_16389; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16654 = _GEN_32735 | _GEN_16390; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16655 = _GEN_32736 | _GEN_16391; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16656 = _T_136 ? _GEN_16648 : _GEN_16384; // @[sequencer-master.scala 154:24]
  wire  _GEN_16657 = _T_136 ? _GEN_16649 : _GEN_16385; // @[sequencer-master.scala 154:24]
  wire  _GEN_16658 = _T_136 ? _GEN_16650 : _GEN_16386; // @[sequencer-master.scala 154:24]
  wire  _GEN_16659 = _T_136 ? _GEN_16651 : _GEN_16387; // @[sequencer-master.scala 154:24]
  wire  _GEN_16660 = _T_136 ? _GEN_16652 : _GEN_16388; // @[sequencer-master.scala 154:24]
  wire  _GEN_16661 = _T_136 ? _GEN_16653 : _GEN_16389; // @[sequencer-master.scala 154:24]
  wire  _GEN_16662 = _T_136 ? _GEN_16654 : _GEN_16390; // @[sequencer-master.scala 154:24]
  wire  _GEN_16663 = _T_136 ? _GEN_16655 : _GEN_16391; // @[sequencer-master.scala 154:24]
  wire  _GEN_16664 = _GEN_32729 | _GEN_16408; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16665 = _GEN_32730 | _GEN_16409; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16666 = _GEN_32731 | _GEN_16410; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16667 = _GEN_32732 | _GEN_16411; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16668 = _GEN_32733 | _GEN_16412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16669 = _GEN_32734 | _GEN_16413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16670 = _GEN_32735 | _GEN_16414; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16671 = _GEN_32736 | _GEN_16415; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16672 = _T_158 ? _GEN_16664 : _GEN_16408; // @[sequencer-master.scala 154:24]
  wire  _GEN_16673 = _T_158 ? _GEN_16665 : _GEN_16409; // @[sequencer-master.scala 154:24]
  wire  _GEN_16674 = _T_158 ? _GEN_16666 : _GEN_16410; // @[sequencer-master.scala 154:24]
  wire  _GEN_16675 = _T_158 ? _GEN_16667 : _GEN_16411; // @[sequencer-master.scala 154:24]
  wire  _GEN_16676 = _T_158 ? _GEN_16668 : _GEN_16412; // @[sequencer-master.scala 154:24]
  wire  _GEN_16677 = _T_158 ? _GEN_16669 : _GEN_16413; // @[sequencer-master.scala 154:24]
  wire  _GEN_16678 = _T_158 ? _GEN_16670 : _GEN_16414; // @[sequencer-master.scala 154:24]
  wire  _GEN_16679 = _T_158 ? _GEN_16671 : _GEN_16415; // @[sequencer-master.scala 154:24]
  wire  _GEN_16680 = _GEN_32729 | _GEN_16432; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16681 = _GEN_32730 | _GEN_16433; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16682 = _GEN_32731 | _GEN_16434; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16683 = _GEN_32732 | _GEN_16435; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16684 = _GEN_32733 | _GEN_16436; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16685 = _GEN_32734 | _GEN_16437; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16686 = _GEN_32735 | _GEN_16438; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16687 = _GEN_32736 | _GEN_16439; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_16688 = _T_180 ? _GEN_16680 : _GEN_16432; // @[sequencer-master.scala 154:24]
  wire  _GEN_16689 = _T_180 ? _GEN_16681 : _GEN_16433; // @[sequencer-master.scala 154:24]
  wire  _GEN_16690 = _T_180 ? _GEN_16682 : _GEN_16434; // @[sequencer-master.scala 154:24]
  wire  _GEN_16691 = _T_180 ? _GEN_16683 : _GEN_16435; // @[sequencer-master.scala 154:24]
  wire  _GEN_16692 = _T_180 ? _GEN_16684 : _GEN_16436; // @[sequencer-master.scala 154:24]
  wire  _GEN_16693 = _T_180 ? _GEN_16685 : _GEN_16437; // @[sequencer-master.scala 154:24]
  wire  _GEN_16694 = _T_180 ? _GEN_16686 : _GEN_16438; // @[sequencer-master.scala 154:24]
  wire  _GEN_16695 = _T_180 ? _GEN_16687 : _GEN_16439; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_16696 = 3'h0 == tail ? _T_1615[1:0] : _GEN_16174; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16697 = 3'h1 == tail ? _T_1615[1:0] : _GEN_16175; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16698 = 3'h2 == tail ? _T_1615[1:0] : _GEN_16176; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16699 = 3'h3 == tail ? _T_1615[1:0] : _GEN_16177; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16700 = 3'h4 == tail ? _T_1615[1:0] : _GEN_16178; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16701 = 3'h5 == tail ? _T_1615[1:0] : _GEN_16179; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16702 = 3'h6 == tail ? _T_1615[1:0] : _GEN_16180; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_16703 = 3'h7 == tail ? _T_1615[1:0] : _GEN_16181; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_16704 = 3'h0 == tail ? 4'h0 : _GEN_16182; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16705 = 3'h1 == tail ? 4'h0 : _GEN_16183; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16706 = 3'h2 == tail ? 4'h0 : _GEN_16184; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16707 = 3'h3 == tail ? 4'h0 : _GEN_16185; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16708 = 3'h4 == tail ? 4'h0 : _GEN_16186; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16709 = 3'h5 == tail ? 4'h0 : _GEN_16187; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16710 = 3'h6 == tail ? 4'h0 : _GEN_16188; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_16711 = 3'h7 == tail ? 4'h0 : _GEN_16189; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_16712 = 3'h0 == tail ? 3'h0 : _GEN_16190; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16713 = 3'h1 == tail ? 3'h0 : _GEN_16191; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16714 = 3'h2 == tail ? 3'h0 : _GEN_16192; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16715 = 3'h3 == tail ? 3'h0 : _GEN_16193; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16716 = 3'h4 == tail ? 3'h0 : _GEN_16194; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16717 = 3'h5 == tail ? 3'h0 : _GEN_16195; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16718 = 3'h6 == tail ? 3'h0 : _GEN_16196; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_16719 = 3'h7 == tail ? 3'h0 : _GEN_16197; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_16720 = io_op_bits_active_vrpred ? _GEN_16200 : _GEN_15766; // @[sequencer-master.scala 648:41]
  wire  _GEN_16721 = io_op_bits_active_vrpred ? _GEN_16201 : _GEN_15767; // @[sequencer-master.scala 648:41]
  wire  _GEN_16722 = io_op_bits_active_vrpred ? _GEN_16202 : _GEN_15768; // @[sequencer-master.scala 648:41]
  wire  _GEN_16723 = io_op_bits_active_vrpred ? _GEN_16203 : _GEN_15769; // @[sequencer-master.scala 648:41]
  wire  _GEN_16724 = io_op_bits_active_vrpred ? _GEN_16204 : _GEN_15770; // @[sequencer-master.scala 648:41]
  wire  _GEN_16725 = io_op_bits_active_vrpred ? _GEN_16205 : _GEN_15771; // @[sequencer-master.scala 648:41]
  wire  _GEN_16726 = io_op_bits_active_vrpred ? _GEN_16206 : _GEN_15772; // @[sequencer-master.scala 648:41]
  wire  _GEN_16727 = io_op_bits_active_vrpred ? _GEN_16207 : _GEN_15773; // @[sequencer-master.scala 648:41]
  wire  _GEN_16736 = io_op_bits_active_vrpred ? _GEN_16536 : _GEN_15782; // @[sequencer-master.scala 648:41]
  wire  _GEN_16737 = io_op_bits_active_vrpred ? _GEN_16537 : _GEN_15783; // @[sequencer-master.scala 648:41]
  wire  _GEN_16738 = io_op_bits_active_vrpred ? _GEN_16538 : _GEN_15784; // @[sequencer-master.scala 648:41]
  wire  _GEN_16739 = io_op_bits_active_vrpred ? _GEN_16539 : _GEN_15785; // @[sequencer-master.scala 648:41]
  wire  _GEN_16740 = io_op_bits_active_vrpred ? _GEN_16540 : _GEN_15786; // @[sequencer-master.scala 648:41]
  wire  _GEN_16741 = io_op_bits_active_vrpred ? _GEN_16541 : _GEN_15787; // @[sequencer-master.scala 648:41]
  wire  _GEN_16742 = io_op_bits_active_vrpred ? _GEN_16542 : _GEN_15788; // @[sequencer-master.scala 648:41]
  wire  _GEN_16743 = io_op_bits_active_vrpred ? _GEN_16543 : _GEN_15789; // @[sequencer-master.scala 648:41]
  wire  _GEN_16744 = io_op_bits_active_vrpred ? _GEN_16224 : _GEN_15790; // @[sequencer-master.scala 648:41]
  wire  _GEN_16745 = io_op_bits_active_vrpred ? _GEN_16225 : _GEN_15791; // @[sequencer-master.scala 648:41]
  wire  _GEN_16746 = io_op_bits_active_vrpred ? _GEN_16226 : _GEN_15792; // @[sequencer-master.scala 648:41]
  wire  _GEN_16747 = io_op_bits_active_vrpred ? _GEN_16227 : _GEN_15793; // @[sequencer-master.scala 648:41]
  wire  _GEN_16748 = io_op_bits_active_vrpred ? _GEN_16228 : _GEN_15794; // @[sequencer-master.scala 648:41]
  wire  _GEN_16749 = io_op_bits_active_vrpred ? _GEN_16229 : _GEN_15795; // @[sequencer-master.scala 648:41]
  wire  _GEN_16750 = io_op_bits_active_vrpred ? _GEN_16230 : _GEN_15796; // @[sequencer-master.scala 648:41]
  wire  _GEN_16751 = io_op_bits_active_vrpred ? _GEN_16231 : _GEN_15797; // @[sequencer-master.scala 648:41]
  wire  _GEN_16752 = io_op_bits_active_vrpred ? _GEN_16232 : _GEN_15798; // @[sequencer-master.scala 648:41]
  wire  _GEN_16753 = io_op_bits_active_vrpred ? _GEN_16233 : _GEN_15799; // @[sequencer-master.scala 648:41]
  wire  _GEN_16754 = io_op_bits_active_vrpred ? _GEN_16234 : _GEN_15800; // @[sequencer-master.scala 648:41]
  wire  _GEN_16755 = io_op_bits_active_vrpred ? _GEN_16235 : _GEN_15801; // @[sequencer-master.scala 648:41]
  wire  _GEN_16756 = io_op_bits_active_vrpred ? _GEN_16236 : _GEN_15802; // @[sequencer-master.scala 648:41]
  wire  _GEN_16757 = io_op_bits_active_vrpred ? _GEN_16237 : _GEN_15803; // @[sequencer-master.scala 648:41]
  wire  _GEN_16758 = io_op_bits_active_vrpred ? _GEN_16238 : _GEN_15804; // @[sequencer-master.scala 648:41]
  wire  _GEN_16759 = io_op_bits_active_vrpred ? _GEN_16239 : _GEN_15805; // @[sequencer-master.scala 648:41]
  wire  _GEN_16760 = io_op_bits_active_vrpred ? _GEN_16240 : _GEN_15806; // @[sequencer-master.scala 648:41]
  wire  _GEN_16761 = io_op_bits_active_vrpred ? _GEN_16241 : _GEN_15807; // @[sequencer-master.scala 648:41]
  wire  _GEN_16762 = io_op_bits_active_vrpred ? _GEN_16242 : _GEN_15808; // @[sequencer-master.scala 648:41]
  wire  _GEN_16763 = io_op_bits_active_vrpred ? _GEN_16243 : _GEN_15809; // @[sequencer-master.scala 648:41]
  wire  _GEN_16764 = io_op_bits_active_vrpred ? _GEN_16244 : _GEN_15810; // @[sequencer-master.scala 648:41]
  wire  _GEN_16765 = io_op_bits_active_vrpred ? _GEN_16245 : _GEN_15811; // @[sequencer-master.scala 648:41]
  wire  _GEN_16766 = io_op_bits_active_vrpred ? _GEN_16246 : _GEN_15812; // @[sequencer-master.scala 648:41]
  wire  _GEN_16767 = io_op_bits_active_vrpred ? _GEN_16247 : _GEN_15813; // @[sequencer-master.scala 648:41]
  wire  _GEN_16768 = io_op_bits_active_vrpred ? _GEN_16248 : _GEN_15814; // @[sequencer-master.scala 648:41]
  wire  _GEN_16769 = io_op_bits_active_vrpred ? _GEN_16249 : _GEN_15815; // @[sequencer-master.scala 648:41]
  wire  _GEN_16770 = io_op_bits_active_vrpred ? _GEN_16250 : _GEN_15816; // @[sequencer-master.scala 648:41]
  wire  _GEN_16771 = io_op_bits_active_vrpred ? _GEN_16251 : _GEN_15817; // @[sequencer-master.scala 648:41]
  wire  _GEN_16772 = io_op_bits_active_vrpred ? _GEN_16252 : _GEN_15818; // @[sequencer-master.scala 648:41]
  wire  _GEN_16773 = io_op_bits_active_vrpred ? _GEN_16253 : _GEN_15819; // @[sequencer-master.scala 648:41]
  wire  _GEN_16774 = io_op_bits_active_vrpred ? _GEN_16254 : _GEN_15820; // @[sequencer-master.scala 648:41]
  wire  _GEN_16775 = io_op_bits_active_vrpred ? _GEN_16255 : _GEN_15821; // @[sequencer-master.scala 648:41]
  wire  _GEN_16776 = io_op_bits_active_vrpred ? _GEN_16256 : _GEN_15822; // @[sequencer-master.scala 648:41]
  wire  _GEN_16777 = io_op_bits_active_vrpred ? _GEN_16257 : _GEN_15823; // @[sequencer-master.scala 648:41]
  wire  _GEN_16778 = io_op_bits_active_vrpred ? _GEN_16258 : _GEN_15824; // @[sequencer-master.scala 648:41]
  wire  _GEN_16779 = io_op_bits_active_vrpred ? _GEN_16259 : _GEN_15825; // @[sequencer-master.scala 648:41]
  wire  _GEN_16780 = io_op_bits_active_vrpred ? _GEN_16260 : _GEN_15826; // @[sequencer-master.scala 648:41]
  wire  _GEN_16781 = io_op_bits_active_vrpred ? _GEN_16261 : _GEN_15827; // @[sequencer-master.scala 648:41]
  wire  _GEN_16782 = io_op_bits_active_vrpred ? _GEN_16262 : _GEN_15828; // @[sequencer-master.scala 648:41]
  wire  _GEN_16783 = io_op_bits_active_vrpred ? _GEN_16263 : _GEN_15829; // @[sequencer-master.scala 648:41]
  wire  _GEN_16784 = io_op_bits_active_vrpred ? _GEN_16576 : _GEN_15830; // @[sequencer-master.scala 648:41]
  wire  _GEN_16785 = io_op_bits_active_vrpred ? _GEN_16577 : _GEN_15831; // @[sequencer-master.scala 648:41]
  wire  _GEN_16786 = io_op_bits_active_vrpred ? _GEN_16578 : _GEN_15832; // @[sequencer-master.scala 648:41]
  wire  _GEN_16787 = io_op_bits_active_vrpred ? _GEN_16579 : _GEN_15833; // @[sequencer-master.scala 648:41]
  wire  _GEN_16788 = io_op_bits_active_vrpred ? _GEN_16580 : _GEN_15834; // @[sequencer-master.scala 648:41]
  wire  _GEN_16789 = io_op_bits_active_vrpred ? _GEN_16581 : _GEN_15835; // @[sequencer-master.scala 648:41]
  wire  _GEN_16790 = io_op_bits_active_vrpred ? _GEN_16582 : _GEN_15836; // @[sequencer-master.scala 648:41]
  wire  _GEN_16791 = io_op_bits_active_vrpred ? _GEN_16583 : _GEN_15837; // @[sequencer-master.scala 648:41]
  wire  _GEN_16792 = io_op_bits_active_vrpred ? _GEN_16272 : _GEN_15838; // @[sequencer-master.scala 648:41]
  wire  _GEN_16793 = io_op_bits_active_vrpred ? _GEN_16273 : _GEN_15839; // @[sequencer-master.scala 648:41]
  wire  _GEN_16794 = io_op_bits_active_vrpred ? _GEN_16274 : _GEN_15840; // @[sequencer-master.scala 648:41]
  wire  _GEN_16795 = io_op_bits_active_vrpred ? _GEN_16275 : _GEN_15841; // @[sequencer-master.scala 648:41]
  wire  _GEN_16796 = io_op_bits_active_vrpred ? _GEN_16276 : _GEN_15842; // @[sequencer-master.scala 648:41]
  wire  _GEN_16797 = io_op_bits_active_vrpred ? _GEN_16277 : _GEN_15843; // @[sequencer-master.scala 648:41]
  wire  _GEN_16798 = io_op_bits_active_vrpred ? _GEN_16278 : _GEN_15844; // @[sequencer-master.scala 648:41]
  wire  _GEN_16799 = io_op_bits_active_vrpred ? _GEN_16279 : _GEN_15845; // @[sequencer-master.scala 648:41]
  wire  _GEN_16800 = io_op_bits_active_vrpred ? _GEN_16280 : _GEN_15846; // @[sequencer-master.scala 648:41]
  wire  _GEN_16801 = io_op_bits_active_vrpred ? _GEN_16281 : _GEN_15847; // @[sequencer-master.scala 648:41]
  wire  _GEN_16802 = io_op_bits_active_vrpred ? _GEN_16282 : _GEN_15848; // @[sequencer-master.scala 648:41]
  wire  _GEN_16803 = io_op_bits_active_vrpred ? _GEN_16283 : _GEN_15849; // @[sequencer-master.scala 648:41]
  wire  _GEN_16804 = io_op_bits_active_vrpred ? _GEN_16284 : _GEN_15850; // @[sequencer-master.scala 648:41]
  wire  _GEN_16805 = io_op_bits_active_vrpred ? _GEN_16285 : _GEN_15851; // @[sequencer-master.scala 648:41]
  wire  _GEN_16806 = io_op_bits_active_vrpred ? _GEN_16286 : _GEN_15852; // @[sequencer-master.scala 648:41]
  wire  _GEN_16807 = io_op_bits_active_vrpred ? _GEN_16287 : _GEN_15853; // @[sequencer-master.scala 648:41]
  wire  _GEN_16808 = io_op_bits_active_vrpred ? _GEN_16592 : _GEN_15854; // @[sequencer-master.scala 648:41]
  wire  _GEN_16809 = io_op_bits_active_vrpred ? _GEN_16593 : _GEN_15855; // @[sequencer-master.scala 648:41]
  wire  _GEN_16810 = io_op_bits_active_vrpred ? _GEN_16594 : _GEN_15856; // @[sequencer-master.scala 648:41]
  wire  _GEN_16811 = io_op_bits_active_vrpred ? _GEN_16595 : _GEN_15857; // @[sequencer-master.scala 648:41]
  wire  _GEN_16812 = io_op_bits_active_vrpred ? _GEN_16596 : _GEN_15858; // @[sequencer-master.scala 648:41]
  wire  _GEN_16813 = io_op_bits_active_vrpred ? _GEN_16597 : _GEN_15859; // @[sequencer-master.scala 648:41]
  wire  _GEN_16814 = io_op_bits_active_vrpred ? _GEN_16598 : _GEN_15860; // @[sequencer-master.scala 648:41]
  wire  _GEN_16815 = io_op_bits_active_vrpred ? _GEN_16599 : _GEN_15861; // @[sequencer-master.scala 648:41]
  wire  _GEN_16816 = io_op_bits_active_vrpred ? _GEN_16296 : _GEN_15862; // @[sequencer-master.scala 648:41]
  wire  _GEN_16817 = io_op_bits_active_vrpred ? _GEN_16297 : _GEN_15863; // @[sequencer-master.scala 648:41]
  wire  _GEN_16818 = io_op_bits_active_vrpred ? _GEN_16298 : _GEN_15864; // @[sequencer-master.scala 648:41]
  wire  _GEN_16819 = io_op_bits_active_vrpred ? _GEN_16299 : _GEN_15865; // @[sequencer-master.scala 648:41]
  wire  _GEN_16820 = io_op_bits_active_vrpred ? _GEN_16300 : _GEN_15866; // @[sequencer-master.scala 648:41]
  wire  _GEN_16821 = io_op_bits_active_vrpred ? _GEN_16301 : _GEN_15867; // @[sequencer-master.scala 648:41]
  wire  _GEN_16822 = io_op_bits_active_vrpred ? _GEN_16302 : _GEN_15868; // @[sequencer-master.scala 648:41]
  wire  _GEN_16823 = io_op_bits_active_vrpred ? _GEN_16303 : _GEN_15869; // @[sequencer-master.scala 648:41]
  wire  _GEN_16824 = io_op_bits_active_vrpred ? _GEN_16304 : _GEN_15870; // @[sequencer-master.scala 648:41]
  wire  _GEN_16825 = io_op_bits_active_vrpred ? _GEN_16305 : _GEN_15871; // @[sequencer-master.scala 648:41]
  wire  _GEN_16826 = io_op_bits_active_vrpred ? _GEN_16306 : _GEN_15872; // @[sequencer-master.scala 648:41]
  wire  _GEN_16827 = io_op_bits_active_vrpred ? _GEN_16307 : _GEN_15873; // @[sequencer-master.scala 648:41]
  wire  _GEN_16828 = io_op_bits_active_vrpred ? _GEN_16308 : _GEN_15874; // @[sequencer-master.scala 648:41]
  wire  _GEN_16829 = io_op_bits_active_vrpred ? _GEN_16309 : _GEN_15875; // @[sequencer-master.scala 648:41]
  wire  _GEN_16830 = io_op_bits_active_vrpred ? _GEN_16310 : _GEN_15876; // @[sequencer-master.scala 648:41]
  wire  _GEN_16831 = io_op_bits_active_vrpred ? _GEN_16311 : _GEN_15877; // @[sequencer-master.scala 648:41]
  wire  _GEN_16832 = io_op_bits_active_vrpred ? _GEN_16608 : _GEN_15878; // @[sequencer-master.scala 648:41]
  wire  _GEN_16833 = io_op_bits_active_vrpred ? _GEN_16609 : _GEN_15879; // @[sequencer-master.scala 648:41]
  wire  _GEN_16834 = io_op_bits_active_vrpred ? _GEN_16610 : _GEN_15880; // @[sequencer-master.scala 648:41]
  wire  _GEN_16835 = io_op_bits_active_vrpred ? _GEN_16611 : _GEN_15881; // @[sequencer-master.scala 648:41]
  wire  _GEN_16836 = io_op_bits_active_vrpred ? _GEN_16612 : _GEN_15882; // @[sequencer-master.scala 648:41]
  wire  _GEN_16837 = io_op_bits_active_vrpred ? _GEN_16613 : _GEN_15883; // @[sequencer-master.scala 648:41]
  wire  _GEN_16838 = io_op_bits_active_vrpred ? _GEN_16614 : _GEN_15884; // @[sequencer-master.scala 648:41]
  wire  _GEN_16839 = io_op_bits_active_vrpred ? _GEN_16615 : _GEN_15885; // @[sequencer-master.scala 648:41]
  wire  _GEN_16840 = io_op_bits_active_vrpred ? _GEN_16320 : _GEN_15886; // @[sequencer-master.scala 648:41]
  wire  _GEN_16841 = io_op_bits_active_vrpred ? _GEN_16321 : _GEN_15887; // @[sequencer-master.scala 648:41]
  wire  _GEN_16842 = io_op_bits_active_vrpred ? _GEN_16322 : _GEN_15888; // @[sequencer-master.scala 648:41]
  wire  _GEN_16843 = io_op_bits_active_vrpred ? _GEN_16323 : _GEN_15889; // @[sequencer-master.scala 648:41]
  wire  _GEN_16844 = io_op_bits_active_vrpred ? _GEN_16324 : _GEN_15890; // @[sequencer-master.scala 648:41]
  wire  _GEN_16845 = io_op_bits_active_vrpred ? _GEN_16325 : _GEN_15891; // @[sequencer-master.scala 648:41]
  wire  _GEN_16846 = io_op_bits_active_vrpred ? _GEN_16326 : _GEN_15892; // @[sequencer-master.scala 648:41]
  wire  _GEN_16847 = io_op_bits_active_vrpred ? _GEN_16327 : _GEN_15893; // @[sequencer-master.scala 648:41]
  wire  _GEN_16848 = io_op_bits_active_vrpred ? _GEN_16328 : _GEN_15894; // @[sequencer-master.scala 648:41]
  wire  _GEN_16849 = io_op_bits_active_vrpred ? _GEN_16329 : _GEN_15895; // @[sequencer-master.scala 648:41]
  wire  _GEN_16850 = io_op_bits_active_vrpred ? _GEN_16330 : _GEN_15896; // @[sequencer-master.scala 648:41]
  wire  _GEN_16851 = io_op_bits_active_vrpred ? _GEN_16331 : _GEN_15897; // @[sequencer-master.scala 648:41]
  wire  _GEN_16852 = io_op_bits_active_vrpred ? _GEN_16332 : _GEN_15898; // @[sequencer-master.scala 648:41]
  wire  _GEN_16853 = io_op_bits_active_vrpred ? _GEN_16333 : _GEN_15899; // @[sequencer-master.scala 648:41]
  wire  _GEN_16854 = io_op_bits_active_vrpred ? _GEN_16334 : _GEN_15900; // @[sequencer-master.scala 648:41]
  wire  _GEN_16855 = io_op_bits_active_vrpred ? _GEN_16335 : _GEN_15901; // @[sequencer-master.scala 648:41]
  wire  _GEN_16856 = io_op_bits_active_vrpred ? _GEN_16624 : _GEN_15902; // @[sequencer-master.scala 648:41]
  wire  _GEN_16857 = io_op_bits_active_vrpred ? _GEN_16625 : _GEN_15903; // @[sequencer-master.scala 648:41]
  wire  _GEN_16858 = io_op_bits_active_vrpred ? _GEN_16626 : _GEN_15904; // @[sequencer-master.scala 648:41]
  wire  _GEN_16859 = io_op_bits_active_vrpred ? _GEN_16627 : _GEN_15905; // @[sequencer-master.scala 648:41]
  wire  _GEN_16860 = io_op_bits_active_vrpred ? _GEN_16628 : _GEN_15906; // @[sequencer-master.scala 648:41]
  wire  _GEN_16861 = io_op_bits_active_vrpred ? _GEN_16629 : _GEN_15907; // @[sequencer-master.scala 648:41]
  wire  _GEN_16862 = io_op_bits_active_vrpred ? _GEN_16630 : _GEN_15908; // @[sequencer-master.scala 648:41]
  wire  _GEN_16863 = io_op_bits_active_vrpred ? _GEN_16631 : _GEN_15909; // @[sequencer-master.scala 648:41]
  wire  _GEN_16864 = io_op_bits_active_vrpred ? _GEN_16344 : _GEN_15910; // @[sequencer-master.scala 648:41]
  wire  _GEN_16865 = io_op_bits_active_vrpred ? _GEN_16345 : _GEN_15911; // @[sequencer-master.scala 648:41]
  wire  _GEN_16866 = io_op_bits_active_vrpred ? _GEN_16346 : _GEN_15912; // @[sequencer-master.scala 648:41]
  wire  _GEN_16867 = io_op_bits_active_vrpred ? _GEN_16347 : _GEN_15913; // @[sequencer-master.scala 648:41]
  wire  _GEN_16868 = io_op_bits_active_vrpred ? _GEN_16348 : _GEN_15914; // @[sequencer-master.scala 648:41]
  wire  _GEN_16869 = io_op_bits_active_vrpred ? _GEN_16349 : _GEN_15915; // @[sequencer-master.scala 648:41]
  wire  _GEN_16870 = io_op_bits_active_vrpred ? _GEN_16350 : _GEN_15916; // @[sequencer-master.scala 648:41]
  wire  _GEN_16871 = io_op_bits_active_vrpred ? _GEN_16351 : _GEN_15917; // @[sequencer-master.scala 648:41]
  wire  _GEN_16872 = io_op_bits_active_vrpred ? _GEN_16352 : _GEN_15918; // @[sequencer-master.scala 648:41]
  wire  _GEN_16873 = io_op_bits_active_vrpred ? _GEN_16353 : _GEN_15919; // @[sequencer-master.scala 648:41]
  wire  _GEN_16874 = io_op_bits_active_vrpred ? _GEN_16354 : _GEN_15920; // @[sequencer-master.scala 648:41]
  wire  _GEN_16875 = io_op_bits_active_vrpred ? _GEN_16355 : _GEN_15921; // @[sequencer-master.scala 648:41]
  wire  _GEN_16876 = io_op_bits_active_vrpred ? _GEN_16356 : _GEN_15922; // @[sequencer-master.scala 648:41]
  wire  _GEN_16877 = io_op_bits_active_vrpred ? _GEN_16357 : _GEN_15923; // @[sequencer-master.scala 648:41]
  wire  _GEN_16878 = io_op_bits_active_vrpred ? _GEN_16358 : _GEN_15924; // @[sequencer-master.scala 648:41]
  wire  _GEN_16879 = io_op_bits_active_vrpred ? _GEN_16359 : _GEN_15925; // @[sequencer-master.scala 648:41]
  wire  _GEN_16880 = io_op_bits_active_vrpred ? _GEN_16640 : _GEN_15926; // @[sequencer-master.scala 648:41]
  wire  _GEN_16881 = io_op_bits_active_vrpred ? _GEN_16641 : _GEN_15927; // @[sequencer-master.scala 648:41]
  wire  _GEN_16882 = io_op_bits_active_vrpred ? _GEN_16642 : _GEN_15928; // @[sequencer-master.scala 648:41]
  wire  _GEN_16883 = io_op_bits_active_vrpred ? _GEN_16643 : _GEN_15929; // @[sequencer-master.scala 648:41]
  wire  _GEN_16884 = io_op_bits_active_vrpred ? _GEN_16644 : _GEN_15930; // @[sequencer-master.scala 648:41]
  wire  _GEN_16885 = io_op_bits_active_vrpred ? _GEN_16645 : _GEN_15931; // @[sequencer-master.scala 648:41]
  wire  _GEN_16886 = io_op_bits_active_vrpred ? _GEN_16646 : _GEN_15932; // @[sequencer-master.scala 648:41]
  wire  _GEN_16887 = io_op_bits_active_vrpred ? _GEN_16647 : _GEN_15933; // @[sequencer-master.scala 648:41]
  wire  _GEN_16888 = io_op_bits_active_vrpred ? _GEN_16368 : _GEN_15934; // @[sequencer-master.scala 648:41]
  wire  _GEN_16889 = io_op_bits_active_vrpred ? _GEN_16369 : _GEN_15935; // @[sequencer-master.scala 648:41]
  wire  _GEN_16890 = io_op_bits_active_vrpred ? _GEN_16370 : _GEN_15936; // @[sequencer-master.scala 648:41]
  wire  _GEN_16891 = io_op_bits_active_vrpred ? _GEN_16371 : _GEN_15937; // @[sequencer-master.scala 648:41]
  wire  _GEN_16892 = io_op_bits_active_vrpred ? _GEN_16372 : _GEN_15938; // @[sequencer-master.scala 648:41]
  wire  _GEN_16893 = io_op_bits_active_vrpred ? _GEN_16373 : _GEN_15939; // @[sequencer-master.scala 648:41]
  wire  _GEN_16894 = io_op_bits_active_vrpred ? _GEN_16374 : _GEN_15940; // @[sequencer-master.scala 648:41]
  wire  _GEN_16895 = io_op_bits_active_vrpred ? _GEN_16375 : _GEN_15941; // @[sequencer-master.scala 648:41]
  wire  _GEN_16896 = io_op_bits_active_vrpred ? _GEN_16376 : _GEN_15942; // @[sequencer-master.scala 648:41]
  wire  _GEN_16897 = io_op_bits_active_vrpred ? _GEN_16377 : _GEN_15943; // @[sequencer-master.scala 648:41]
  wire  _GEN_16898 = io_op_bits_active_vrpred ? _GEN_16378 : _GEN_15944; // @[sequencer-master.scala 648:41]
  wire  _GEN_16899 = io_op_bits_active_vrpred ? _GEN_16379 : _GEN_15945; // @[sequencer-master.scala 648:41]
  wire  _GEN_16900 = io_op_bits_active_vrpred ? _GEN_16380 : _GEN_15946; // @[sequencer-master.scala 648:41]
  wire  _GEN_16901 = io_op_bits_active_vrpred ? _GEN_16381 : _GEN_15947; // @[sequencer-master.scala 648:41]
  wire  _GEN_16902 = io_op_bits_active_vrpred ? _GEN_16382 : _GEN_15948; // @[sequencer-master.scala 648:41]
  wire  _GEN_16903 = io_op_bits_active_vrpred ? _GEN_16383 : _GEN_15949; // @[sequencer-master.scala 648:41]
  wire  _GEN_16904 = io_op_bits_active_vrpred ? _GEN_16656 : _GEN_15950; // @[sequencer-master.scala 648:41]
  wire  _GEN_16905 = io_op_bits_active_vrpred ? _GEN_16657 : _GEN_15951; // @[sequencer-master.scala 648:41]
  wire  _GEN_16906 = io_op_bits_active_vrpred ? _GEN_16658 : _GEN_15952; // @[sequencer-master.scala 648:41]
  wire  _GEN_16907 = io_op_bits_active_vrpred ? _GEN_16659 : _GEN_15953; // @[sequencer-master.scala 648:41]
  wire  _GEN_16908 = io_op_bits_active_vrpred ? _GEN_16660 : _GEN_15954; // @[sequencer-master.scala 648:41]
  wire  _GEN_16909 = io_op_bits_active_vrpred ? _GEN_16661 : _GEN_15955; // @[sequencer-master.scala 648:41]
  wire  _GEN_16910 = io_op_bits_active_vrpred ? _GEN_16662 : _GEN_15956; // @[sequencer-master.scala 648:41]
  wire  _GEN_16911 = io_op_bits_active_vrpred ? _GEN_16663 : _GEN_15957; // @[sequencer-master.scala 648:41]
  wire  _GEN_16912 = io_op_bits_active_vrpred ? _GEN_16392 : _GEN_15958; // @[sequencer-master.scala 648:41]
  wire  _GEN_16913 = io_op_bits_active_vrpred ? _GEN_16393 : _GEN_15959; // @[sequencer-master.scala 648:41]
  wire  _GEN_16914 = io_op_bits_active_vrpred ? _GEN_16394 : _GEN_15960; // @[sequencer-master.scala 648:41]
  wire  _GEN_16915 = io_op_bits_active_vrpred ? _GEN_16395 : _GEN_15961; // @[sequencer-master.scala 648:41]
  wire  _GEN_16916 = io_op_bits_active_vrpred ? _GEN_16396 : _GEN_15962; // @[sequencer-master.scala 648:41]
  wire  _GEN_16917 = io_op_bits_active_vrpred ? _GEN_16397 : _GEN_15963; // @[sequencer-master.scala 648:41]
  wire  _GEN_16918 = io_op_bits_active_vrpred ? _GEN_16398 : _GEN_15964; // @[sequencer-master.scala 648:41]
  wire  _GEN_16919 = io_op_bits_active_vrpred ? _GEN_16399 : _GEN_15965; // @[sequencer-master.scala 648:41]
  wire  _GEN_16920 = io_op_bits_active_vrpred ? _GEN_16400 : _GEN_15966; // @[sequencer-master.scala 648:41]
  wire  _GEN_16921 = io_op_bits_active_vrpred ? _GEN_16401 : _GEN_15967; // @[sequencer-master.scala 648:41]
  wire  _GEN_16922 = io_op_bits_active_vrpred ? _GEN_16402 : _GEN_15968; // @[sequencer-master.scala 648:41]
  wire  _GEN_16923 = io_op_bits_active_vrpred ? _GEN_16403 : _GEN_15969; // @[sequencer-master.scala 648:41]
  wire  _GEN_16924 = io_op_bits_active_vrpred ? _GEN_16404 : _GEN_15970; // @[sequencer-master.scala 648:41]
  wire  _GEN_16925 = io_op_bits_active_vrpred ? _GEN_16405 : _GEN_15971; // @[sequencer-master.scala 648:41]
  wire  _GEN_16926 = io_op_bits_active_vrpred ? _GEN_16406 : _GEN_15972; // @[sequencer-master.scala 648:41]
  wire  _GEN_16927 = io_op_bits_active_vrpred ? _GEN_16407 : _GEN_15973; // @[sequencer-master.scala 648:41]
  wire  _GEN_16928 = io_op_bits_active_vrpred ? _GEN_16672 : _GEN_15974; // @[sequencer-master.scala 648:41]
  wire  _GEN_16929 = io_op_bits_active_vrpred ? _GEN_16673 : _GEN_15975; // @[sequencer-master.scala 648:41]
  wire  _GEN_16930 = io_op_bits_active_vrpred ? _GEN_16674 : _GEN_15976; // @[sequencer-master.scala 648:41]
  wire  _GEN_16931 = io_op_bits_active_vrpred ? _GEN_16675 : _GEN_15977; // @[sequencer-master.scala 648:41]
  wire  _GEN_16932 = io_op_bits_active_vrpred ? _GEN_16676 : _GEN_15978; // @[sequencer-master.scala 648:41]
  wire  _GEN_16933 = io_op_bits_active_vrpred ? _GEN_16677 : _GEN_15979; // @[sequencer-master.scala 648:41]
  wire  _GEN_16934 = io_op_bits_active_vrpred ? _GEN_16678 : _GEN_15980; // @[sequencer-master.scala 648:41]
  wire  _GEN_16935 = io_op_bits_active_vrpred ? _GEN_16679 : _GEN_15981; // @[sequencer-master.scala 648:41]
  wire  _GEN_16936 = io_op_bits_active_vrpred ? _GEN_16416 : _GEN_15982; // @[sequencer-master.scala 648:41]
  wire  _GEN_16937 = io_op_bits_active_vrpred ? _GEN_16417 : _GEN_15983; // @[sequencer-master.scala 648:41]
  wire  _GEN_16938 = io_op_bits_active_vrpred ? _GEN_16418 : _GEN_15984; // @[sequencer-master.scala 648:41]
  wire  _GEN_16939 = io_op_bits_active_vrpred ? _GEN_16419 : _GEN_15985; // @[sequencer-master.scala 648:41]
  wire  _GEN_16940 = io_op_bits_active_vrpred ? _GEN_16420 : _GEN_15986; // @[sequencer-master.scala 648:41]
  wire  _GEN_16941 = io_op_bits_active_vrpred ? _GEN_16421 : _GEN_15987; // @[sequencer-master.scala 648:41]
  wire  _GEN_16942 = io_op_bits_active_vrpred ? _GEN_16422 : _GEN_15988; // @[sequencer-master.scala 648:41]
  wire  _GEN_16943 = io_op_bits_active_vrpred ? _GEN_16423 : _GEN_15989; // @[sequencer-master.scala 648:41]
  wire  _GEN_16944 = io_op_bits_active_vrpred ? _GEN_16424 : _GEN_15990; // @[sequencer-master.scala 648:41]
  wire  _GEN_16945 = io_op_bits_active_vrpred ? _GEN_16425 : _GEN_15991; // @[sequencer-master.scala 648:41]
  wire  _GEN_16946 = io_op_bits_active_vrpred ? _GEN_16426 : _GEN_15992; // @[sequencer-master.scala 648:41]
  wire  _GEN_16947 = io_op_bits_active_vrpred ? _GEN_16427 : _GEN_15993; // @[sequencer-master.scala 648:41]
  wire  _GEN_16948 = io_op_bits_active_vrpred ? _GEN_16428 : _GEN_15994; // @[sequencer-master.scala 648:41]
  wire  _GEN_16949 = io_op_bits_active_vrpred ? _GEN_16429 : _GEN_15995; // @[sequencer-master.scala 648:41]
  wire  _GEN_16950 = io_op_bits_active_vrpred ? _GEN_16430 : _GEN_15996; // @[sequencer-master.scala 648:41]
  wire  _GEN_16951 = io_op_bits_active_vrpred ? _GEN_16431 : _GEN_15997; // @[sequencer-master.scala 648:41]
  wire  _GEN_16952 = io_op_bits_active_vrpred ? _GEN_16688 : _GEN_15998; // @[sequencer-master.scala 648:41]
  wire  _GEN_16953 = io_op_bits_active_vrpred ? _GEN_16689 : _GEN_15999; // @[sequencer-master.scala 648:41]
  wire  _GEN_16954 = io_op_bits_active_vrpred ? _GEN_16690 : _GEN_16000; // @[sequencer-master.scala 648:41]
  wire  _GEN_16955 = io_op_bits_active_vrpred ? _GEN_16691 : _GEN_16001; // @[sequencer-master.scala 648:41]
  wire  _GEN_16956 = io_op_bits_active_vrpred ? _GEN_16692 : _GEN_16002; // @[sequencer-master.scala 648:41]
  wire  _GEN_16957 = io_op_bits_active_vrpred ? _GEN_16693 : _GEN_16003; // @[sequencer-master.scala 648:41]
  wire  _GEN_16958 = io_op_bits_active_vrpred ? _GEN_16694 : _GEN_16004; // @[sequencer-master.scala 648:41]
  wire  _GEN_16959 = io_op_bits_active_vrpred ? _GEN_16695 : _GEN_16005; // @[sequencer-master.scala 648:41]
  wire  _GEN_16960 = io_op_bits_active_vrpred ? _GEN_16440 : _GEN_16006; // @[sequencer-master.scala 648:41]
  wire  _GEN_16961 = io_op_bits_active_vrpred ? _GEN_16441 : _GEN_16007; // @[sequencer-master.scala 648:41]
  wire  _GEN_16962 = io_op_bits_active_vrpred ? _GEN_16442 : _GEN_16008; // @[sequencer-master.scala 648:41]
  wire  _GEN_16963 = io_op_bits_active_vrpred ? _GEN_16443 : _GEN_16009; // @[sequencer-master.scala 648:41]
  wire  _GEN_16964 = io_op_bits_active_vrpred ? _GEN_16444 : _GEN_16010; // @[sequencer-master.scala 648:41]
  wire  _GEN_16965 = io_op_bits_active_vrpred ? _GEN_16445 : _GEN_16011; // @[sequencer-master.scala 648:41]
  wire  _GEN_16966 = io_op_bits_active_vrpred ? _GEN_16446 : _GEN_16012; // @[sequencer-master.scala 648:41]
  wire  _GEN_16967 = io_op_bits_active_vrpred ? _GEN_16447 : _GEN_16013; // @[sequencer-master.scala 648:41]
  wire  _GEN_16968 = io_op_bits_active_vrpred ? _GEN_16448 : _GEN_16014; // @[sequencer-master.scala 648:41]
  wire  _GEN_16969 = io_op_bits_active_vrpred ? _GEN_16449 : _GEN_16015; // @[sequencer-master.scala 648:41]
  wire  _GEN_16970 = io_op_bits_active_vrpred ? _GEN_16450 : _GEN_16016; // @[sequencer-master.scala 648:41]
  wire  _GEN_16971 = io_op_bits_active_vrpred ? _GEN_16451 : _GEN_16017; // @[sequencer-master.scala 648:41]
  wire  _GEN_16972 = io_op_bits_active_vrpred ? _GEN_16452 : _GEN_16018; // @[sequencer-master.scala 648:41]
  wire  _GEN_16973 = io_op_bits_active_vrpred ? _GEN_16453 : _GEN_16019; // @[sequencer-master.scala 648:41]
  wire  _GEN_16974 = io_op_bits_active_vrpred ? _GEN_16454 : _GEN_16020; // @[sequencer-master.scala 648:41]
  wire  _GEN_16975 = io_op_bits_active_vrpred ? _GEN_16455 : _GEN_16021; // @[sequencer-master.scala 648:41]
  wire  _GEN_16976 = io_op_bits_active_vrpred ? _GEN_16456 : _GEN_16022; // @[sequencer-master.scala 648:41]
  wire  _GEN_16977 = io_op_bits_active_vrpred ? _GEN_16457 : _GEN_16023; // @[sequencer-master.scala 648:41]
  wire  _GEN_16978 = io_op_bits_active_vrpred ? _GEN_16458 : _GEN_16024; // @[sequencer-master.scala 648:41]
  wire  _GEN_16979 = io_op_bits_active_vrpred ? _GEN_16459 : _GEN_16025; // @[sequencer-master.scala 648:41]
  wire  _GEN_16980 = io_op_bits_active_vrpred ? _GEN_16460 : _GEN_16026; // @[sequencer-master.scala 648:41]
  wire  _GEN_16981 = io_op_bits_active_vrpred ? _GEN_16461 : _GEN_16027; // @[sequencer-master.scala 648:41]
  wire  _GEN_16982 = io_op_bits_active_vrpred ? _GEN_16462 : _GEN_16028; // @[sequencer-master.scala 648:41]
  wire  _GEN_16983 = io_op_bits_active_vrpred ? _GEN_16463 : _GEN_16029; // @[sequencer-master.scala 648:41]
  wire  _GEN_16992 = io_op_bits_active_vrpred ? _GEN_16472 : _GEN_12514; // @[sequencer-master.scala 648:41]
  wire  _GEN_16993 = io_op_bits_active_vrpred ? _GEN_16473 : _GEN_12515; // @[sequencer-master.scala 648:41]
  wire  _GEN_16994 = io_op_bits_active_vrpred ? _GEN_16474 : _GEN_12516; // @[sequencer-master.scala 648:41]
  wire  _GEN_16995 = io_op_bits_active_vrpred ? _GEN_16475 : _GEN_12517; // @[sequencer-master.scala 648:41]
  wire  _GEN_16996 = io_op_bits_active_vrpred ? _GEN_16476 : _GEN_12518; // @[sequencer-master.scala 648:41]
  wire  _GEN_16997 = io_op_bits_active_vrpred ? _GEN_16477 : _GEN_12519; // @[sequencer-master.scala 648:41]
  wire  _GEN_16998 = io_op_bits_active_vrpred ? _GEN_16478 : _GEN_12520; // @[sequencer-master.scala 648:41]
  wire  _GEN_16999 = io_op_bits_active_vrpred ? _GEN_16479 : _GEN_12521; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17000 = io_op_bits_active_vrpred ? _GEN_16480 : _GEN_16046; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17001 = io_op_bits_active_vrpred ? _GEN_16481 : _GEN_16047; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17002 = io_op_bits_active_vrpred ? _GEN_16482 : _GEN_16048; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17003 = io_op_bits_active_vrpred ? _GEN_16483 : _GEN_16049; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17004 = io_op_bits_active_vrpred ? _GEN_16484 : _GEN_16050; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17005 = io_op_bits_active_vrpred ? _GEN_16485 : _GEN_16051; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17006 = io_op_bits_active_vrpred ? _GEN_16486 : _GEN_16052; // @[sequencer-master.scala 648:41]
  wire [9:0] _GEN_17007 = io_op_bits_active_vrpred ? _GEN_16487 : _GEN_16053; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17008 = io_op_bits_active_vrpred ? _GEN_16528 : _GEN_16054; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17009 = io_op_bits_active_vrpred ? _GEN_16529 : _GEN_16055; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17010 = io_op_bits_active_vrpred ? _GEN_16530 : _GEN_16056; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17011 = io_op_bits_active_vrpred ? _GEN_16531 : _GEN_16057; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17012 = io_op_bits_active_vrpred ? _GEN_16532 : _GEN_16058; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17013 = io_op_bits_active_vrpred ? _GEN_16533 : _GEN_16059; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17014 = io_op_bits_active_vrpred ? _GEN_16534 : _GEN_16060; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17015 = io_op_bits_active_vrpred ? _GEN_16535 : _GEN_16061; // @[sequencer-master.scala 648:41]
  wire  _GEN_17016 = io_op_bits_active_vrpred ? _GEN_16544 : _GEN_16062; // @[sequencer-master.scala 648:41]
  wire  _GEN_17017 = io_op_bits_active_vrpred ? _GEN_16545 : _GEN_16063; // @[sequencer-master.scala 648:41]
  wire  _GEN_17018 = io_op_bits_active_vrpred ? _GEN_16546 : _GEN_16064; // @[sequencer-master.scala 648:41]
  wire  _GEN_17019 = io_op_bits_active_vrpred ? _GEN_16547 : _GEN_16065; // @[sequencer-master.scala 648:41]
  wire  _GEN_17020 = io_op_bits_active_vrpred ? _GEN_16548 : _GEN_16066; // @[sequencer-master.scala 648:41]
  wire  _GEN_17021 = io_op_bits_active_vrpred ? _GEN_16549 : _GEN_16067; // @[sequencer-master.scala 648:41]
  wire  _GEN_17022 = io_op_bits_active_vrpred ? _GEN_16550 : _GEN_16068; // @[sequencer-master.scala 648:41]
  wire  _GEN_17023 = io_op_bits_active_vrpred ? _GEN_16551 : _GEN_16069; // @[sequencer-master.scala 648:41]
  wire  _GEN_17024 = io_op_bits_active_vrpred ? _GEN_16552 : _GEN_16070; // @[sequencer-master.scala 648:41]
  wire  _GEN_17025 = io_op_bits_active_vrpred ? _GEN_16553 : _GEN_16071; // @[sequencer-master.scala 648:41]
  wire  _GEN_17026 = io_op_bits_active_vrpred ? _GEN_16554 : _GEN_16072; // @[sequencer-master.scala 648:41]
  wire  _GEN_17027 = io_op_bits_active_vrpred ? _GEN_16555 : _GEN_16073; // @[sequencer-master.scala 648:41]
  wire  _GEN_17028 = io_op_bits_active_vrpred ? _GEN_16556 : _GEN_16074; // @[sequencer-master.scala 648:41]
  wire  _GEN_17029 = io_op_bits_active_vrpred ? _GEN_16557 : _GEN_16075; // @[sequencer-master.scala 648:41]
  wire  _GEN_17030 = io_op_bits_active_vrpred ? _GEN_16558 : _GEN_16076; // @[sequencer-master.scala 648:41]
  wire  _GEN_17031 = io_op_bits_active_vrpred ? _GEN_16559 : _GEN_16077; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17032 = io_op_bits_active_vrpred ? _GEN_16560 : _GEN_16078; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17033 = io_op_bits_active_vrpred ? _GEN_16561 : _GEN_16079; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17034 = io_op_bits_active_vrpred ? _GEN_16562 : _GEN_16080; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17035 = io_op_bits_active_vrpred ? _GEN_16563 : _GEN_16081; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17036 = io_op_bits_active_vrpred ? _GEN_16564 : _GEN_16082; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17037 = io_op_bits_active_vrpred ? _GEN_16565 : _GEN_16083; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17038 = io_op_bits_active_vrpred ? _GEN_16566 : _GEN_16084; // @[sequencer-master.scala 648:41]
  wire [7:0] _GEN_17039 = io_op_bits_active_vrpred ? _GEN_16567 : _GEN_16085; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17040 = io_op_bits_active_vrpred ? _GEN_16696 : _GEN_16174; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17041 = io_op_bits_active_vrpred ? _GEN_16697 : _GEN_16175; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17042 = io_op_bits_active_vrpred ? _GEN_16698 : _GEN_16176; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17043 = io_op_bits_active_vrpred ? _GEN_16699 : _GEN_16177; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17044 = io_op_bits_active_vrpred ? _GEN_16700 : _GEN_16178; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17045 = io_op_bits_active_vrpred ? _GEN_16701 : _GEN_16179; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17046 = io_op_bits_active_vrpred ? _GEN_16702 : _GEN_16180; // @[sequencer-master.scala 648:41]
  wire [1:0] _GEN_17047 = io_op_bits_active_vrpred ? _GEN_16703 : _GEN_16181; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17048 = io_op_bits_active_vrpred ? _GEN_16704 : _GEN_16182; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17049 = io_op_bits_active_vrpred ? _GEN_16705 : _GEN_16183; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17050 = io_op_bits_active_vrpred ? _GEN_16706 : _GEN_16184; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17051 = io_op_bits_active_vrpred ? _GEN_16707 : _GEN_16185; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17052 = io_op_bits_active_vrpred ? _GEN_16708 : _GEN_16186; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17053 = io_op_bits_active_vrpred ? _GEN_16709 : _GEN_16187; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17054 = io_op_bits_active_vrpred ? _GEN_16710 : _GEN_16188; // @[sequencer-master.scala 648:41]
  wire [3:0] _GEN_17055 = io_op_bits_active_vrpred ? _GEN_16711 : _GEN_16189; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17056 = io_op_bits_active_vrpred ? _GEN_16712 : _GEN_16190; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17057 = io_op_bits_active_vrpred ? _GEN_16713 : _GEN_16191; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17058 = io_op_bits_active_vrpred ? _GEN_16714 : _GEN_16192; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17059 = io_op_bits_active_vrpred ? _GEN_16715 : _GEN_16193; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17060 = io_op_bits_active_vrpred ? _GEN_16716 : _GEN_16194; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17061 = io_op_bits_active_vrpred ? _GEN_16717 : _GEN_16195; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17062 = io_op_bits_active_vrpred ? _GEN_16718 : _GEN_16196; // @[sequencer-master.scala 648:41]
  wire [2:0] _GEN_17063 = io_op_bits_active_vrpred ? _GEN_16719 : _GEN_16197; // @[sequencer-master.scala 648:41]
  wire  _GEN_17064 = io_op_bits_active_vrpred | _GEN_16198; // @[sequencer-master.scala 648:41 sequencer-master.scala 265:41]
  wire [2:0] _GEN_17065 = io_op_bits_active_vrpred ? _T_1645 : _GEN_16199; // @[sequencer-master.scala 648:41 sequencer-master.scala 265:66]
  wire  _GEN_17066 = _GEN_32729 | _GEN_16720; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17067 = _GEN_32730 | _GEN_16721; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17068 = _GEN_32731 | _GEN_16722; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17069 = _GEN_32732 | _GEN_16723; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17070 = _GEN_32733 | _GEN_16724; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17071 = _GEN_32734 | _GEN_16725; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17072 = _GEN_32735 | _GEN_16726; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17073 = _GEN_32736 | _GEN_16727; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_17082 = 3'h0 == tail ? 1'h0 : _GEN_16736; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17083 = 3'h1 == tail ? 1'h0 : _GEN_16737; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17084 = 3'h2 == tail ? 1'h0 : _GEN_16738; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17085 = 3'h3 == tail ? 1'h0 : _GEN_16739; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17086 = 3'h4 == tail ? 1'h0 : _GEN_16740; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17087 = 3'h5 == tail ? 1'h0 : _GEN_16741; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17088 = 3'h6 == tail ? 1'h0 : _GEN_16742; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17089 = 3'h7 == tail ? 1'h0 : _GEN_16743; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_17090 = 3'h0 == tail ? 1'h0 : _GEN_16744; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17091 = 3'h1 == tail ? 1'h0 : _GEN_16745; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17092 = 3'h2 == tail ? 1'h0 : _GEN_16746; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17093 = 3'h3 == tail ? 1'h0 : _GEN_16747; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17094 = 3'h4 == tail ? 1'h0 : _GEN_16748; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17095 = 3'h5 == tail ? 1'h0 : _GEN_16749; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17096 = 3'h6 == tail ? 1'h0 : _GEN_16750; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17097 = 3'h7 == tail ? 1'h0 : _GEN_16751; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_17098 = 3'h0 == tail ? 1'h0 : _GEN_16752; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17099 = 3'h1 == tail ? 1'h0 : _GEN_16753; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17100 = 3'h2 == tail ? 1'h0 : _GEN_16754; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17101 = 3'h3 == tail ? 1'h0 : _GEN_16755; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17102 = 3'h4 == tail ? 1'h0 : _GEN_16756; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17103 = 3'h5 == tail ? 1'h0 : _GEN_16757; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17104 = 3'h6 == tail ? 1'h0 : _GEN_16758; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17105 = 3'h7 == tail ? 1'h0 : _GEN_16759; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_17106 = 3'h0 == tail ? 1'h0 : _GEN_16760; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17107 = 3'h1 == tail ? 1'h0 : _GEN_16761; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17108 = 3'h2 == tail ? 1'h0 : _GEN_16762; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17109 = 3'h3 == tail ? 1'h0 : _GEN_16763; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17110 = 3'h4 == tail ? 1'h0 : _GEN_16764; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17111 = 3'h5 == tail ? 1'h0 : _GEN_16765; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17112 = 3'h6 == tail ? 1'h0 : _GEN_16766; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17113 = 3'h7 == tail ? 1'h0 : _GEN_16767; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_17114 = 3'h0 == tail ? 1'h0 : _GEN_16768; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17115 = 3'h1 == tail ? 1'h0 : _GEN_16769; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17116 = 3'h2 == tail ? 1'h0 : _GEN_16770; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17117 = 3'h3 == tail ? 1'h0 : _GEN_16771; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17118 = 3'h4 == tail ? 1'h0 : _GEN_16772; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17119 = 3'h5 == tail ? 1'h0 : _GEN_16773; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17120 = 3'h6 == tail ? 1'h0 : _GEN_16774; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17121 = 3'h7 == tail ? 1'h0 : _GEN_16775; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_17122 = _GEN_32729 | _GEN_16776; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17123 = _GEN_32730 | _GEN_16777; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17124 = _GEN_32731 | _GEN_16778; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17125 = _GEN_32732 | _GEN_16779; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17126 = _GEN_32733 | _GEN_16780; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17127 = _GEN_32734 | _GEN_16781; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17128 = _GEN_32735 | _GEN_16782; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17129 = _GEN_32736 | _GEN_16783; // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_17130 = 3'h0 == tail ? 1'h0 : _GEN_16784; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17131 = 3'h1 == tail ? 1'h0 : _GEN_16785; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17132 = 3'h2 == tail ? 1'h0 : _GEN_16786; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17133 = 3'h3 == tail ? 1'h0 : _GEN_16787; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17134 = 3'h4 == tail ? 1'h0 : _GEN_16788; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17135 = 3'h5 == tail ? 1'h0 : _GEN_16789; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17136 = 3'h6 == tail ? 1'h0 : _GEN_16790; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17137 = 3'h7 == tail ? 1'h0 : _GEN_16791; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17138 = 3'h0 == tail ? 1'h0 : _GEN_16792; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17139 = 3'h1 == tail ? 1'h0 : _GEN_16793; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17140 = 3'h2 == tail ? 1'h0 : _GEN_16794; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17141 = 3'h3 == tail ? 1'h0 : _GEN_16795; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17142 = 3'h4 == tail ? 1'h0 : _GEN_16796; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17143 = 3'h5 == tail ? 1'h0 : _GEN_16797; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17144 = 3'h6 == tail ? 1'h0 : _GEN_16798; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17145 = 3'h7 == tail ? 1'h0 : _GEN_16799; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17146 = 3'h0 == tail ? 1'h0 : _GEN_16800; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17147 = 3'h1 == tail ? 1'h0 : _GEN_16801; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17148 = 3'h2 == tail ? 1'h0 : _GEN_16802; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17149 = 3'h3 == tail ? 1'h0 : _GEN_16803; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17150 = 3'h4 == tail ? 1'h0 : _GEN_16804; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17151 = 3'h5 == tail ? 1'h0 : _GEN_16805; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17152 = 3'h6 == tail ? 1'h0 : _GEN_16806; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17153 = 3'h7 == tail ? 1'h0 : _GEN_16807; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17154 = 3'h0 == tail ? 1'h0 : _GEN_16808; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17155 = 3'h1 == tail ? 1'h0 : _GEN_16809; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17156 = 3'h2 == tail ? 1'h0 : _GEN_16810; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17157 = 3'h3 == tail ? 1'h0 : _GEN_16811; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17158 = 3'h4 == tail ? 1'h0 : _GEN_16812; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17159 = 3'h5 == tail ? 1'h0 : _GEN_16813; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17160 = 3'h6 == tail ? 1'h0 : _GEN_16814; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17161 = 3'h7 == tail ? 1'h0 : _GEN_16815; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17162 = 3'h0 == tail ? 1'h0 : _GEN_16816; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17163 = 3'h1 == tail ? 1'h0 : _GEN_16817; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17164 = 3'h2 == tail ? 1'h0 : _GEN_16818; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17165 = 3'h3 == tail ? 1'h0 : _GEN_16819; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17166 = 3'h4 == tail ? 1'h0 : _GEN_16820; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17167 = 3'h5 == tail ? 1'h0 : _GEN_16821; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17168 = 3'h6 == tail ? 1'h0 : _GEN_16822; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17169 = 3'h7 == tail ? 1'h0 : _GEN_16823; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17170 = 3'h0 == tail ? 1'h0 : _GEN_16824; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17171 = 3'h1 == tail ? 1'h0 : _GEN_16825; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17172 = 3'h2 == tail ? 1'h0 : _GEN_16826; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17173 = 3'h3 == tail ? 1'h0 : _GEN_16827; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17174 = 3'h4 == tail ? 1'h0 : _GEN_16828; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17175 = 3'h5 == tail ? 1'h0 : _GEN_16829; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17176 = 3'h6 == tail ? 1'h0 : _GEN_16830; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17177 = 3'h7 == tail ? 1'h0 : _GEN_16831; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17178 = 3'h0 == tail ? 1'h0 : _GEN_16832; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17179 = 3'h1 == tail ? 1'h0 : _GEN_16833; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17180 = 3'h2 == tail ? 1'h0 : _GEN_16834; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17181 = 3'h3 == tail ? 1'h0 : _GEN_16835; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17182 = 3'h4 == tail ? 1'h0 : _GEN_16836; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17183 = 3'h5 == tail ? 1'h0 : _GEN_16837; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17184 = 3'h6 == tail ? 1'h0 : _GEN_16838; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17185 = 3'h7 == tail ? 1'h0 : _GEN_16839; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17186 = 3'h0 == tail ? 1'h0 : _GEN_16840; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17187 = 3'h1 == tail ? 1'h0 : _GEN_16841; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17188 = 3'h2 == tail ? 1'h0 : _GEN_16842; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17189 = 3'h3 == tail ? 1'h0 : _GEN_16843; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17190 = 3'h4 == tail ? 1'h0 : _GEN_16844; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17191 = 3'h5 == tail ? 1'h0 : _GEN_16845; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17192 = 3'h6 == tail ? 1'h0 : _GEN_16846; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17193 = 3'h7 == tail ? 1'h0 : _GEN_16847; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17194 = 3'h0 == tail ? 1'h0 : _GEN_16848; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17195 = 3'h1 == tail ? 1'h0 : _GEN_16849; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17196 = 3'h2 == tail ? 1'h0 : _GEN_16850; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17197 = 3'h3 == tail ? 1'h0 : _GEN_16851; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17198 = 3'h4 == tail ? 1'h0 : _GEN_16852; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17199 = 3'h5 == tail ? 1'h0 : _GEN_16853; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17200 = 3'h6 == tail ? 1'h0 : _GEN_16854; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17201 = 3'h7 == tail ? 1'h0 : _GEN_16855; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17202 = 3'h0 == tail ? 1'h0 : _GEN_16856; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17203 = 3'h1 == tail ? 1'h0 : _GEN_16857; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17204 = 3'h2 == tail ? 1'h0 : _GEN_16858; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17205 = 3'h3 == tail ? 1'h0 : _GEN_16859; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17206 = 3'h4 == tail ? 1'h0 : _GEN_16860; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17207 = 3'h5 == tail ? 1'h0 : _GEN_16861; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17208 = 3'h6 == tail ? 1'h0 : _GEN_16862; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17209 = 3'h7 == tail ? 1'h0 : _GEN_16863; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17210 = 3'h0 == tail ? 1'h0 : _GEN_16864; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17211 = 3'h1 == tail ? 1'h0 : _GEN_16865; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17212 = 3'h2 == tail ? 1'h0 : _GEN_16866; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17213 = 3'h3 == tail ? 1'h0 : _GEN_16867; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17214 = 3'h4 == tail ? 1'h0 : _GEN_16868; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17215 = 3'h5 == tail ? 1'h0 : _GEN_16869; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17216 = 3'h6 == tail ? 1'h0 : _GEN_16870; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17217 = 3'h7 == tail ? 1'h0 : _GEN_16871; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17218 = 3'h0 == tail ? 1'h0 : _GEN_16872; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17219 = 3'h1 == tail ? 1'h0 : _GEN_16873; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17220 = 3'h2 == tail ? 1'h0 : _GEN_16874; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17221 = 3'h3 == tail ? 1'h0 : _GEN_16875; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17222 = 3'h4 == tail ? 1'h0 : _GEN_16876; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17223 = 3'h5 == tail ? 1'h0 : _GEN_16877; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17224 = 3'h6 == tail ? 1'h0 : _GEN_16878; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17225 = 3'h7 == tail ? 1'h0 : _GEN_16879; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17226 = 3'h0 == tail ? 1'h0 : _GEN_16880; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17227 = 3'h1 == tail ? 1'h0 : _GEN_16881; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17228 = 3'h2 == tail ? 1'h0 : _GEN_16882; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17229 = 3'h3 == tail ? 1'h0 : _GEN_16883; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17230 = 3'h4 == tail ? 1'h0 : _GEN_16884; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17231 = 3'h5 == tail ? 1'h0 : _GEN_16885; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17232 = 3'h6 == tail ? 1'h0 : _GEN_16886; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17233 = 3'h7 == tail ? 1'h0 : _GEN_16887; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17234 = 3'h0 == tail ? 1'h0 : _GEN_16888; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17235 = 3'h1 == tail ? 1'h0 : _GEN_16889; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17236 = 3'h2 == tail ? 1'h0 : _GEN_16890; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17237 = 3'h3 == tail ? 1'h0 : _GEN_16891; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17238 = 3'h4 == tail ? 1'h0 : _GEN_16892; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17239 = 3'h5 == tail ? 1'h0 : _GEN_16893; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17240 = 3'h6 == tail ? 1'h0 : _GEN_16894; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17241 = 3'h7 == tail ? 1'h0 : _GEN_16895; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17242 = 3'h0 == tail ? 1'h0 : _GEN_16896; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17243 = 3'h1 == tail ? 1'h0 : _GEN_16897; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17244 = 3'h2 == tail ? 1'h0 : _GEN_16898; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17245 = 3'h3 == tail ? 1'h0 : _GEN_16899; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17246 = 3'h4 == tail ? 1'h0 : _GEN_16900; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17247 = 3'h5 == tail ? 1'h0 : _GEN_16901; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17248 = 3'h6 == tail ? 1'h0 : _GEN_16902; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17249 = 3'h7 == tail ? 1'h0 : _GEN_16903; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17250 = 3'h0 == tail ? 1'h0 : _GEN_16904; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17251 = 3'h1 == tail ? 1'h0 : _GEN_16905; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17252 = 3'h2 == tail ? 1'h0 : _GEN_16906; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17253 = 3'h3 == tail ? 1'h0 : _GEN_16907; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17254 = 3'h4 == tail ? 1'h0 : _GEN_16908; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17255 = 3'h5 == tail ? 1'h0 : _GEN_16909; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17256 = 3'h6 == tail ? 1'h0 : _GEN_16910; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17257 = 3'h7 == tail ? 1'h0 : _GEN_16911; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17258 = 3'h0 == tail ? 1'h0 : _GEN_16912; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17259 = 3'h1 == tail ? 1'h0 : _GEN_16913; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17260 = 3'h2 == tail ? 1'h0 : _GEN_16914; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17261 = 3'h3 == tail ? 1'h0 : _GEN_16915; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17262 = 3'h4 == tail ? 1'h0 : _GEN_16916; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17263 = 3'h5 == tail ? 1'h0 : _GEN_16917; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17264 = 3'h6 == tail ? 1'h0 : _GEN_16918; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17265 = 3'h7 == tail ? 1'h0 : _GEN_16919; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17266 = 3'h0 == tail ? 1'h0 : _GEN_16920; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17267 = 3'h1 == tail ? 1'h0 : _GEN_16921; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17268 = 3'h2 == tail ? 1'h0 : _GEN_16922; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17269 = 3'h3 == tail ? 1'h0 : _GEN_16923; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17270 = 3'h4 == tail ? 1'h0 : _GEN_16924; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17271 = 3'h5 == tail ? 1'h0 : _GEN_16925; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17272 = 3'h6 == tail ? 1'h0 : _GEN_16926; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17273 = 3'h7 == tail ? 1'h0 : _GEN_16927; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17274 = 3'h0 == tail ? 1'h0 : _GEN_16928; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17275 = 3'h1 == tail ? 1'h0 : _GEN_16929; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17276 = 3'h2 == tail ? 1'h0 : _GEN_16930; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17277 = 3'h3 == tail ? 1'h0 : _GEN_16931; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17278 = 3'h4 == tail ? 1'h0 : _GEN_16932; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17279 = 3'h5 == tail ? 1'h0 : _GEN_16933; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17280 = 3'h6 == tail ? 1'h0 : _GEN_16934; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17281 = 3'h7 == tail ? 1'h0 : _GEN_16935; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17282 = 3'h0 == tail ? 1'h0 : _GEN_16936; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17283 = 3'h1 == tail ? 1'h0 : _GEN_16937; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17284 = 3'h2 == tail ? 1'h0 : _GEN_16938; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17285 = 3'h3 == tail ? 1'h0 : _GEN_16939; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17286 = 3'h4 == tail ? 1'h0 : _GEN_16940; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17287 = 3'h5 == tail ? 1'h0 : _GEN_16941; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17288 = 3'h6 == tail ? 1'h0 : _GEN_16942; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17289 = 3'h7 == tail ? 1'h0 : _GEN_16943; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17290 = 3'h0 == tail ? 1'h0 : _GEN_16944; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17291 = 3'h1 == tail ? 1'h0 : _GEN_16945; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17292 = 3'h2 == tail ? 1'h0 : _GEN_16946; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17293 = 3'h3 == tail ? 1'h0 : _GEN_16947; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17294 = 3'h4 == tail ? 1'h0 : _GEN_16948; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17295 = 3'h5 == tail ? 1'h0 : _GEN_16949; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17296 = 3'h6 == tail ? 1'h0 : _GEN_16950; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17297 = 3'h7 == tail ? 1'h0 : _GEN_16951; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17298 = 3'h0 == tail ? 1'h0 : _GEN_16952; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17299 = 3'h1 == tail ? 1'h0 : _GEN_16953; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17300 = 3'h2 == tail ? 1'h0 : _GEN_16954; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17301 = 3'h3 == tail ? 1'h0 : _GEN_16955; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17302 = 3'h4 == tail ? 1'h0 : _GEN_16956; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17303 = 3'h5 == tail ? 1'h0 : _GEN_16957; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17304 = 3'h6 == tail ? 1'h0 : _GEN_16958; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17305 = 3'h7 == tail ? 1'h0 : _GEN_16959; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_17306 = 3'h0 == tail ? 1'h0 : _GEN_16960; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17307 = 3'h1 == tail ? 1'h0 : _GEN_16961; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17308 = 3'h2 == tail ? 1'h0 : _GEN_16962; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17309 = 3'h3 == tail ? 1'h0 : _GEN_16963; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17310 = 3'h4 == tail ? 1'h0 : _GEN_16964; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17311 = 3'h5 == tail ? 1'h0 : _GEN_16965; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17312 = 3'h6 == tail ? 1'h0 : _GEN_16966; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17313 = 3'h7 == tail ? 1'h0 : _GEN_16967; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_17314 = 3'h0 == tail ? 1'h0 : _GEN_16968; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17315 = 3'h1 == tail ? 1'h0 : _GEN_16969; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17316 = 3'h2 == tail ? 1'h0 : _GEN_16970; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17317 = 3'h3 == tail ? 1'h0 : _GEN_16971; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17318 = 3'h4 == tail ? 1'h0 : _GEN_16972; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17319 = 3'h5 == tail ? 1'h0 : _GEN_16973; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17320 = 3'h6 == tail ? 1'h0 : _GEN_16974; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17321 = 3'h7 == tail ? 1'h0 : _GEN_16975; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_17322 = 3'h0 == tail ? 1'h0 : _GEN_16976; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17323 = 3'h1 == tail ? 1'h0 : _GEN_16977; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17324 = 3'h2 == tail ? 1'h0 : _GEN_16978; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17325 = 3'h3 == tail ? 1'h0 : _GEN_16979; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17326 = 3'h4 == tail ? 1'h0 : _GEN_16980; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17327 = 3'h5 == tail ? 1'h0 : _GEN_16981; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17328 = 3'h6 == tail ? 1'h0 : _GEN_16982; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17329 = 3'h7 == tail ? 1'h0 : _GEN_16983; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_17338 = _GEN_32729 | _GEN_16992; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17339 = _GEN_32730 | _GEN_16993; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17340 = _GEN_32731 | _GEN_16994; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17341 = _GEN_32732 | _GEN_16995; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17342 = _GEN_32733 | _GEN_16996; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17343 = _GEN_32734 | _GEN_16997; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17344 = _GEN_32735 | _GEN_16998; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_17345 = _GEN_32736 | _GEN_16999; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_17346 = 3'h0 == tail ? _e_tail_fn_union_2 : _GEN_17000; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17347 = 3'h1 == tail ? _e_tail_fn_union_2 : _GEN_17001; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17348 = 3'h2 == tail ? _e_tail_fn_union_2 : _GEN_17002; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17349 = 3'h3 == tail ? _e_tail_fn_union_2 : _GEN_17003; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17350 = 3'h4 == tail ? _e_tail_fn_union_2 : _GEN_17004; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17351 = 3'h5 == tail ? _e_tail_fn_union_2 : _GEN_17005; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17352 = 3'h6 == tail ? _e_tail_fn_union_2 : _GEN_17006; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_17353 = 3'h7 == tail ? _e_tail_fn_union_2 : _GEN_17007; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_17354 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_17008; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17355 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_17009; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17356 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_17010; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17357 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_17011; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17358 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_17012; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17359 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_17013; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17360 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_17014; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_17361 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_17015; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17362 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_17082; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17363 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_17083; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17364 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_17084; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17365 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_17085; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17366 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_17086; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17367 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_17087; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17368 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_17088; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17369 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_17089; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17370 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_17016; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17371 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_17017; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17372 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_17018; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17373 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_17019; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17374 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_17020; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17375 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_17021; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17376 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_17022; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17377 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_17023; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17378 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_17024; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17379 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_17025; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17380 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_17026; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17381 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_17027; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17382 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_17028; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17383 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_17029; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17384 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_17030; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_17385 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_17031; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_17386 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_17032; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17387 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_17033; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17388 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_17034; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17389 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_17035; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17390 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_17036; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17391 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_17037; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17392 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_17038; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_17393 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_17039; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_17394 = io_op_bits_base_vp_valid ? _GEN_17354 : _GEN_17008; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17395 = io_op_bits_base_vp_valid ? _GEN_17355 : _GEN_17009; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17396 = io_op_bits_base_vp_valid ? _GEN_17356 : _GEN_17010; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17397 = io_op_bits_base_vp_valid ? _GEN_17357 : _GEN_17011; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17398 = io_op_bits_base_vp_valid ? _GEN_17358 : _GEN_17012; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17399 = io_op_bits_base_vp_valid ? _GEN_17359 : _GEN_17013; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17400 = io_op_bits_base_vp_valid ? _GEN_17360 : _GEN_17014; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_17401 = io_op_bits_base_vp_valid ? _GEN_17361 : _GEN_17015; // @[sequencer-master.scala 320:41]
  wire  _GEN_17402 = io_op_bits_base_vp_valid ? _GEN_17362 : _GEN_17082; // @[sequencer-master.scala 320:41]
  wire  _GEN_17403 = io_op_bits_base_vp_valid ? _GEN_17363 : _GEN_17083; // @[sequencer-master.scala 320:41]
  wire  _GEN_17404 = io_op_bits_base_vp_valid ? _GEN_17364 : _GEN_17084; // @[sequencer-master.scala 320:41]
  wire  _GEN_17405 = io_op_bits_base_vp_valid ? _GEN_17365 : _GEN_17085; // @[sequencer-master.scala 320:41]
  wire  _GEN_17406 = io_op_bits_base_vp_valid ? _GEN_17366 : _GEN_17086; // @[sequencer-master.scala 320:41]
  wire  _GEN_17407 = io_op_bits_base_vp_valid ? _GEN_17367 : _GEN_17087; // @[sequencer-master.scala 320:41]
  wire  _GEN_17408 = io_op_bits_base_vp_valid ? _GEN_17368 : _GEN_17088; // @[sequencer-master.scala 320:41]
  wire  _GEN_17409 = io_op_bits_base_vp_valid ? _GEN_17369 : _GEN_17089; // @[sequencer-master.scala 320:41]
  wire  _GEN_17410 = io_op_bits_base_vp_valid ? _GEN_17370 : _GEN_17016; // @[sequencer-master.scala 320:41]
  wire  _GEN_17411 = io_op_bits_base_vp_valid ? _GEN_17371 : _GEN_17017; // @[sequencer-master.scala 320:41]
  wire  _GEN_17412 = io_op_bits_base_vp_valid ? _GEN_17372 : _GEN_17018; // @[sequencer-master.scala 320:41]
  wire  _GEN_17413 = io_op_bits_base_vp_valid ? _GEN_17373 : _GEN_17019; // @[sequencer-master.scala 320:41]
  wire  _GEN_17414 = io_op_bits_base_vp_valid ? _GEN_17374 : _GEN_17020; // @[sequencer-master.scala 320:41]
  wire  _GEN_17415 = io_op_bits_base_vp_valid ? _GEN_17375 : _GEN_17021; // @[sequencer-master.scala 320:41]
  wire  _GEN_17416 = io_op_bits_base_vp_valid ? _GEN_17376 : _GEN_17022; // @[sequencer-master.scala 320:41]
  wire  _GEN_17417 = io_op_bits_base_vp_valid ? _GEN_17377 : _GEN_17023; // @[sequencer-master.scala 320:41]
  wire  _GEN_17418 = io_op_bits_base_vp_valid ? _GEN_17378 : _GEN_17024; // @[sequencer-master.scala 320:41]
  wire  _GEN_17419 = io_op_bits_base_vp_valid ? _GEN_17379 : _GEN_17025; // @[sequencer-master.scala 320:41]
  wire  _GEN_17420 = io_op_bits_base_vp_valid ? _GEN_17380 : _GEN_17026; // @[sequencer-master.scala 320:41]
  wire  _GEN_17421 = io_op_bits_base_vp_valid ? _GEN_17381 : _GEN_17027; // @[sequencer-master.scala 320:41]
  wire  _GEN_17422 = io_op_bits_base_vp_valid ? _GEN_17382 : _GEN_17028; // @[sequencer-master.scala 320:41]
  wire  _GEN_17423 = io_op_bits_base_vp_valid ? _GEN_17383 : _GEN_17029; // @[sequencer-master.scala 320:41]
  wire  _GEN_17424 = io_op_bits_base_vp_valid ? _GEN_17384 : _GEN_17030; // @[sequencer-master.scala 320:41]
  wire  _GEN_17425 = io_op_bits_base_vp_valid ? _GEN_17385 : _GEN_17031; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17426 = io_op_bits_base_vp_valid ? _GEN_17386 : _GEN_17032; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17427 = io_op_bits_base_vp_valid ? _GEN_17387 : _GEN_17033; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17428 = io_op_bits_base_vp_valid ? _GEN_17388 : _GEN_17034; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17429 = io_op_bits_base_vp_valid ? _GEN_17389 : _GEN_17035; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17430 = io_op_bits_base_vp_valid ? _GEN_17390 : _GEN_17036; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17431 = io_op_bits_base_vp_valid ? _GEN_17391 : _GEN_17037; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17432 = io_op_bits_base_vp_valid ? _GEN_17392 : _GEN_17038; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_17433 = io_op_bits_base_vp_valid ? _GEN_17393 : _GEN_17039; // @[sequencer-master.scala 320:41]
  wire  _GEN_17434 = _GEN_32729 | _GEN_17130; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17435 = _GEN_32730 | _GEN_17131; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17436 = _GEN_32731 | _GEN_17132; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17437 = _GEN_32732 | _GEN_17133; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17438 = _GEN_32733 | _GEN_17134; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17439 = _GEN_32734 | _GEN_17135; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17440 = _GEN_32735 | _GEN_17136; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17441 = _GEN_32736 | _GEN_17137; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17442 = _T_26 ? _GEN_17434 : _GEN_17130; // @[sequencer-master.scala 154:24]
  wire  _GEN_17443 = _T_26 ? _GEN_17435 : _GEN_17131; // @[sequencer-master.scala 154:24]
  wire  _GEN_17444 = _T_26 ? _GEN_17436 : _GEN_17132; // @[sequencer-master.scala 154:24]
  wire  _GEN_17445 = _T_26 ? _GEN_17437 : _GEN_17133; // @[sequencer-master.scala 154:24]
  wire  _GEN_17446 = _T_26 ? _GEN_17438 : _GEN_17134; // @[sequencer-master.scala 154:24]
  wire  _GEN_17447 = _T_26 ? _GEN_17439 : _GEN_17135; // @[sequencer-master.scala 154:24]
  wire  _GEN_17448 = _T_26 ? _GEN_17440 : _GEN_17136; // @[sequencer-master.scala 154:24]
  wire  _GEN_17449 = _T_26 ? _GEN_17441 : _GEN_17137; // @[sequencer-master.scala 154:24]
  wire  _GEN_17450 = _GEN_32729 | _GEN_17154; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17451 = _GEN_32730 | _GEN_17155; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17452 = _GEN_32731 | _GEN_17156; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17453 = _GEN_32732 | _GEN_17157; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17454 = _GEN_32733 | _GEN_17158; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17455 = _GEN_32734 | _GEN_17159; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17456 = _GEN_32735 | _GEN_17160; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17457 = _GEN_32736 | _GEN_17161; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17458 = _T_48 ? _GEN_17450 : _GEN_17154; // @[sequencer-master.scala 154:24]
  wire  _GEN_17459 = _T_48 ? _GEN_17451 : _GEN_17155; // @[sequencer-master.scala 154:24]
  wire  _GEN_17460 = _T_48 ? _GEN_17452 : _GEN_17156; // @[sequencer-master.scala 154:24]
  wire  _GEN_17461 = _T_48 ? _GEN_17453 : _GEN_17157; // @[sequencer-master.scala 154:24]
  wire  _GEN_17462 = _T_48 ? _GEN_17454 : _GEN_17158; // @[sequencer-master.scala 154:24]
  wire  _GEN_17463 = _T_48 ? _GEN_17455 : _GEN_17159; // @[sequencer-master.scala 154:24]
  wire  _GEN_17464 = _T_48 ? _GEN_17456 : _GEN_17160; // @[sequencer-master.scala 154:24]
  wire  _GEN_17465 = _T_48 ? _GEN_17457 : _GEN_17161; // @[sequencer-master.scala 154:24]
  wire  _GEN_17466 = _GEN_32729 | _GEN_17178; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17467 = _GEN_32730 | _GEN_17179; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17468 = _GEN_32731 | _GEN_17180; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17469 = _GEN_32732 | _GEN_17181; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17470 = _GEN_32733 | _GEN_17182; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17471 = _GEN_32734 | _GEN_17183; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17472 = _GEN_32735 | _GEN_17184; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17473 = _GEN_32736 | _GEN_17185; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17474 = _T_70 ? _GEN_17466 : _GEN_17178; // @[sequencer-master.scala 154:24]
  wire  _GEN_17475 = _T_70 ? _GEN_17467 : _GEN_17179; // @[sequencer-master.scala 154:24]
  wire  _GEN_17476 = _T_70 ? _GEN_17468 : _GEN_17180; // @[sequencer-master.scala 154:24]
  wire  _GEN_17477 = _T_70 ? _GEN_17469 : _GEN_17181; // @[sequencer-master.scala 154:24]
  wire  _GEN_17478 = _T_70 ? _GEN_17470 : _GEN_17182; // @[sequencer-master.scala 154:24]
  wire  _GEN_17479 = _T_70 ? _GEN_17471 : _GEN_17183; // @[sequencer-master.scala 154:24]
  wire  _GEN_17480 = _T_70 ? _GEN_17472 : _GEN_17184; // @[sequencer-master.scala 154:24]
  wire  _GEN_17481 = _T_70 ? _GEN_17473 : _GEN_17185; // @[sequencer-master.scala 154:24]
  wire  _GEN_17482 = _GEN_32729 | _GEN_17202; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17483 = _GEN_32730 | _GEN_17203; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17484 = _GEN_32731 | _GEN_17204; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17485 = _GEN_32732 | _GEN_17205; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17486 = _GEN_32733 | _GEN_17206; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17487 = _GEN_32734 | _GEN_17207; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17488 = _GEN_32735 | _GEN_17208; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17489 = _GEN_32736 | _GEN_17209; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17490 = _T_92 ? _GEN_17482 : _GEN_17202; // @[sequencer-master.scala 154:24]
  wire  _GEN_17491 = _T_92 ? _GEN_17483 : _GEN_17203; // @[sequencer-master.scala 154:24]
  wire  _GEN_17492 = _T_92 ? _GEN_17484 : _GEN_17204; // @[sequencer-master.scala 154:24]
  wire  _GEN_17493 = _T_92 ? _GEN_17485 : _GEN_17205; // @[sequencer-master.scala 154:24]
  wire  _GEN_17494 = _T_92 ? _GEN_17486 : _GEN_17206; // @[sequencer-master.scala 154:24]
  wire  _GEN_17495 = _T_92 ? _GEN_17487 : _GEN_17207; // @[sequencer-master.scala 154:24]
  wire  _GEN_17496 = _T_92 ? _GEN_17488 : _GEN_17208; // @[sequencer-master.scala 154:24]
  wire  _GEN_17497 = _T_92 ? _GEN_17489 : _GEN_17209; // @[sequencer-master.scala 154:24]
  wire  _GEN_17498 = _GEN_32729 | _GEN_17226; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17499 = _GEN_32730 | _GEN_17227; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17500 = _GEN_32731 | _GEN_17228; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17501 = _GEN_32732 | _GEN_17229; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17502 = _GEN_32733 | _GEN_17230; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17503 = _GEN_32734 | _GEN_17231; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17504 = _GEN_32735 | _GEN_17232; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17505 = _GEN_32736 | _GEN_17233; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17506 = _T_114 ? _GEN_17498 : _GEN_17226; // @[sequencer-master.scala 154:24]
  wire  _GEN_17507 = _T_114 ? _GEN_17499 : _GEN_17227; // @[sequencer-master.scala 154:24]
  wire  _GEN_17508 = _T_114 ? _GEN_17500 : _GEN_17228; // @[sequencer-master.scala 154:24]
  wire  _GEN_17509 = _T_114 ? _GEN_17501 : _GEN_17229; // @[sequencer-master.scala 154:24]
  wire  _GEN_17510 = _T_114 ? _GEN_17502 : _GEN_17230; // @[sequencer-master.scala 154:24]
  wire  _GEN_17511 = _T_114 ? _GEN_17503 : _GEN_17231; // @[sequencer-master.scala 154:24]
  wire  _GEN_17512 = _T_114 ? _GEN_17504 : _GEN_17232; // @[sequencer-master.scala 154:24]
  wire  _GEN_17513 = _T_114 ? _GEN_17505 : _GEN_17233; // @[sequencer-master.scala 154:24]
  wire  _GEN_17514 = _GEN_32729 | _GEN_17250; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17515 = _GEN_32730 | _GEN_17251; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17516 = _GEN_32731 | _GEN_17252; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17517 = _GEN_32732 | _GEN_17253; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17518 = _GEN_32733 | _GEN_17254; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17519 = _GEN_32734 | _GEN_17255; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17520 = _GEN_32735 | _GEN_17256; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17521 = _GEN_32736 | _GEN_17257; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17522 = _T_136 ? _GEN_17514 : _GEN_17250; // @[sequencer-master.scala 154:24]
  wire  _GEN_17523 = _T_136 ? _GEN_17515 : _GEN_17251; // @[sequencer-master.scala 154:24]
  wire  _GEN_17524 = _T_136 ? _GEN_17516 : _GEN_17252; // @[sequencer-master.scala 154:24]
  wire  _GEN_17525 = _T_136 ? _GEN_17517 : _GEN_17253; // @[sequencer-master.scala 154:24]
  wire  _GEN_17526 = _T_136 ? _GEN_17518 : _GEN_17254; // @[sequencer-master.scala 154:24]
  wire  _GEN_17527 = _T_136 ? _GEN_17519 : _GEN_17255; // @[sequencer-master.scala 154:24]
  wire  _GEN_17528 = _T_136 ? _GEN_17520 : _GEN_17256; // @[sequencer-master.scala 154:24]
  wire  _GEN_17529 = _T_136 ? _GEN_17521 : _GEN_17257; // @[sequencer-master.scala 154:24]
  wire  _GEN_17530 = _GEN_32729 | _GEN_17274; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17531 = _GEN_32730 | _GEN_17275; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17532 = _GEN_32731 | _GEN_17276; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17533 = _GEN_32732 | _GEN_17277; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17534 = _GEN_32733 | _GEN_17278; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17535 = _GEN_32734 | _GEN_17279; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17536 = _GEN_32735 | _GEN_17280; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17537 = _GEN_32736 | _GEN_17281; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17538 = _T_158 ? _GEN_17530 : _GEN_17274; // @[sequencer-master.scala 154:24]
  wire  _GEN_17539 = _T_158 ? _GEN_17531 : _GEN_17275; // @[sequencer-master.scala 154:24]
  wire  _GEN_17540 = _T_158 ? _GEN_17532 : _GEN_17276; // @[sequencer-master.scala 154:24]
  wire  _GEN_17541 = _T_158 ? _GEN_17533 : _GEN_17277; // @[sequencer-master.scala 154:24]
  wire  _GEN_17542 = _T_158 ? _GEN_17534 : _GEN_17278; // @[sequencer-master.scala 154:24]
  wire  _GEN_17543 = _T_158 ? _GEN_17535 : _GEN_17279; // @[sequencer-master.scala 154:24]
  wire  _GEN_17544 = _T_158 ? _GEN_17536 : _GEN_17280; // @[sequencer-master.scala 154:24]
  wire  _GEN_17545 = _T_158 ? _GEN_17537 : _GEN_17281; // @[sequencer-master.scala 154:24]
  wire  _GEN_17546 = _GEN_32729 | _GEN_17298; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17547 = _GEN_32730 | _GEN_17299; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17548 = _GEN_32731 | _GEN_17300; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17549 = _GEN_32732 | _GEN_17301; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17550 = _GEN_32733 | _GEN_17302; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17551 = _GEN_32734 | _GEN_17303; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17552 = _GEN_32735 | _GEN_17304; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17553 = _GEN_32736 | _GEN_17305; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17554 = _T_180 ? _GEN_17546 : _GEN_17298; // @[sequencer-master.scala 154:24]
  wire  _GEN_17555 = _T_180 ? _GEN_17547 : _GEN_17299; // @[sequencer-master.scala 154:24]
  wire  _GEN_17556 = _T_180 ? _GEN_17548 : _GEN_17300; // @[sequencer-master.scala 154:24]
  wire  _GEN_17557 = _T_180 ? _GEN_17549 : _GEN_17301; // @[sequencer-master.scala 154:24]
  wire  _GEN_17558 = _T_180 ? _GEN_17550 : _GEN_17302; // @[sequencer-master.scala 154:24]
  wire  _GEN_17559 = _T_180 ? _GEN_17551 : _GEN_17303; // @[sequencer-master.scala 154:24]
  wire  _GEN_17560 = _T_180 ? _GEN_17552 : _GEN_17304; // @[sequencer-master.scala 154:24]
  wire  _GEN_17561 = _T_180 ? _GEN_17553 : _GEN_17305; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_17562 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_16086; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17563 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_16087; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17564 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_16088; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17565 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_16089; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17566 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_16090; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17567 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_16091; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17568 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_16092; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17569 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_16093; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17570 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_17090; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17571 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_17091; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17572 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_17092; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17573 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_17093; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17574 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_17094; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17575 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_17095; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17576 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_17096; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17577 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_17097; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17578 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_16094; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17579 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_16095; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17580 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_16096; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17581 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_16097; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17582 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_16098; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17583 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_16099; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17584 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_16100; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17585 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_16101; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17586 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_16102; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17587 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_16103; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17588 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_16104; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17589 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_16105; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17590 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_16106; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17591 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_16107; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17592 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_16108; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_17593 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_16109; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17594 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_16110; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17595 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_16111; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17596 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_16112; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17597 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_16113; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17598 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_16114; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17599 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_16115; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17600 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_16116; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_17601 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_16117; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_17602 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_16118; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17603 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_16119; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17604 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_16120; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17605 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_16121; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17606 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_16122; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17607 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_16123; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17608 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_16124; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_17609 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_16125; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_17610 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_16126; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17611 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_16127; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17612 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_16128; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17613 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_16129; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17614 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_16130; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17615 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_16131; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17616 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_16132; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17617 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_16133; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_17618 = _T_189 ? _GEN_17610 : _GEN_16126; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17619 = _T_189 ? _GEN_17611 : _GEN_16127; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17620 = _T_189 ? _GEN_17612 : _GEN_16128; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17621 = _T_189 ? _GEN_17613 : _GEN_16129; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17622 = _T_189 ? _GEN_17614 : _GEN_16130; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17623 = _T_189 ? _GEN_17615 : _GEN_16131; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17624 = _T_189 ? _GEN_17616 : _GEN_16132; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_17625 = _T_189 ? _GEN_17617 : _GEN_16133; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_17626 = io_op_bits_base_vs1_valid ? _GEN_17562 : _GEN_16086; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17627 = io_op_bits_base_vs1_valid ? _GEN_17563 : _GEN_16087; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17628 = io_op_bits_base_vs1_valid ? _GEN_17564 : _GEN_16088; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17629 = io_op_bits_base_vs1_valid ? _GEN_17565 : _GEN_16089; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17630 = io_op_bits_base_vs1_valid ? _GEN_17566 : _GEN_16090; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17631 = io_op_bits_base_vs1_valid ? _GEN_17567 : _GEN_16091; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17632 = io_op_bits_base_vs1_valid ? _GEN_17568 : _GEN_16092; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17633 = io_op_bits_base_vs1_valid ? _GEN_17569 : _GEN_16093; // @[sequencer-master.scala 328:47]
  wire  _GEN_17634 = io_op_bits_base_vs1_valid ? _GEN_17570 : _GEN_17090; // @[sequencer-master.scala 328:47]
  wire  _GEN_17635 = io_op_bits_base_vs1_valid ? _GEN_17571 : _GEN_17091; // @[sequencer-master.scala 328:47]
  wire  _GEN_17636 = io_op_bits_base_vs1_valid ? _GEN_17572 : _GEN_17092; // @[sequencer-master.scala 328:47]
  wire  _GEN_17637 = io_op_bits_base_vs1_valid ? _GEN_17573 : _GEN_17093; // @[sequencer-master.scala 328:47]
  wire  _GEN_17638 = io_op_bits_base_vs1_valid ? _GEN_17574 : _GEN_17094; // @[sequencer-master.scala 328:47]
  wire  _GEN_17639 = io_op_bits_base_vs1_valid ? _GEN_17575 : _GEN_17095; // @[sequencer-master.scala 328:47]
  wire  _GEN_17640 = io_op_bits_base_vs1_valid ? _GEN_17576 : _GEN_17096; // @[sequencer-master.scala 328:47]
  wire  _GEN_17641 = io_op_bits_base_vs1_valid ? _GEN_17577 : _GEN_17097; // @[sequencer-master.scala 328:47]
  wire  _GEN_17642 = io_op_bits_base_vs1_valid ? _GEN_17578 : _GEN_16094; // @[sequencer-master.scala 328:47]
  wire  _GEN_17643 = io_op_bits_base_vs1_valid ? _GEN_17579 : _GEN_16095; // @[sequencer-master.scala 328:47]
  wire  _GEN_17644 = io_op_bits_base_vs1_valid ? _GEN_17580 : _GEN_16096; // @[sequencer-master.scala 328:47]
  wire  _GEN_17645 = io_op_bits_base_vs1_valid ? _GEN_17581 : _GEN_16097; // @[sequencer-master.scala 328:47]
  wire  _GEN_17646 = io_op_bits_base_vs1_valid ? _GEN_17582 : _GEN_16098; // @[sequencer-master.scala 328:47]
  wire  _GEN_17647 = io_op_bits_base_vs1_valid ? _GEN_17583 : _GEN_16099; // @[sequencer-master.scala 328:47]
  wire  _GEN_17648 = io_op_bits_base_vs1_valid ? _GEN_17584 : _GEN_16100; // @[sequencer-master.scala 328:47]
  wire  _GEN_17649 = io_op_bits_base_vs1_valid ? _GEN_17585 : _GEN_16101; // @[sequencer-master.scala 328:47]
  wire  _GEN_17650 = io_op_bits_base_vs1_valid ? _GEN_17586 : _GEN_16102; // @[sequencer-master.scala 328:47]
  wire  _GEN_17651 = io_op_bits_base_vs1_valid ? _GEN_17587 : _GEN_16103; // @[sequencer-master.scala 328:47]
  wire  _GEN_17652 = io_op_bits_base_vs1_valid ? _GEN_17588 : _GEN_16104; // @[sequencer-master.scala 328:47]
  wire  _GEN_17653 = io_op_bits_base_vs1_valid ? _GEN_17589 : _GEN_16105; // @[sequencer-master.scala 328:47]
  wire  _GEN_17654 = io_op_bits_base_vs1_valid ? _GEN_17590 : _GEN_16106; // @[sequencer-master.scala 328:47]
  wire  _GEN_17655 = io_op_bits_base_vs1_valid ? _GEN_17591 : _GEN_16107; // @[sequencer-master.scala 328:47]
  wire  _GEN_17656 = io_op_bits_base_vs1_valid ? _GEN_17592 : _GEN_16108; // @[sequencer-master.scala 328:47]
  wire  _GEN_17657 = io_op_bits_base_vs1_valid ? _GEN_17593 : _GEN_16109; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17658 = io_op_bits_base_vs1_valid ? _GEN_17594 : _GEN_16110; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17659 = io_op_bits_base_vs1_valid ? _GEN_17595 : _GEN_16111; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17660 = io_op_bits_base_vs1_valid ? _GEN_17596 : _GEN_16112; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17661 = io_op_bits_base_vs1_valid ? _GEN_17597 : _GEN_16113; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17662 = io_op_bits_base_vs1_valid ? _GEN_17598 : _GEN_16114; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17663 = io_op_bits_base_vs1_valid ? _GEN_17599 : _GEN_16115; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17664 = io_op_bits_base_vs1_valid ? _GEN_17600 : _GEN_16116; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_17665 = io_op_bits_base_vs1_valid ? _GEN_17601 : _GEN_16117; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17666 = io_op_bits_base_vs1_valid ? _GEN_17602 : _GEN_16118; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17667 = io_op_bits_base_vs1_valid ? _GEN_17603 : _GEN_16119; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17668 = io_op_bits_base_vs1_valid ? _GEN_17604 : _GEN_16120; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17669 = io_op_bits_base_vs1_valid ? _GEN_17605 : _GEN_16121; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17670 = io_op_bits_base_vs1_valid ? _GEN_17606 : _GEN_16122; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17671 = io_op_bits_base_vs1_valid ? _GEN_17607 : _GEN_16123; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17672 = io_op_bits_base_vs1_valid ? _GEN_17608 : _GEN_16124; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_17673 = io_op_bits_base_vs1_valid ? _GEN_17609 : _GEN_16125; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17674 = io_op_bits_base_vs1_valid ? _GEN_17618 : _GEN_16126; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17675 = io_op_bits_base_vs1_valid ? _GEN_17619 : _GEN_16127; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17676 = io_op_bits_base_vs1_valid ? _GEN_17620 : _GEN_16128; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17677 = io_op_bits_base_vs1_valid ? _GEN_17621 : _GEN_16129; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17678 = io_op_bits_base_vs1_valid ? _GEN_17622 : _GEN_16130; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17679 = io_op_bits_base_vs1_valid ? _GEN_17623 : _GEN_16131; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17680 = io_op_bits_base_vs1_valid ? _GEN_17624 : _GEN_16132; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_17681 = io_op_bits_base_vs1_valid ? _GEN_17625 : _GEN_16133; // @[sequencer-master.scala 328:47]
  wire  _GEN_17682 = _GEN_32729 | _GEN_17442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17683 = _GEN_32730 | _GEN_17443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17684 = _GEN_32731 | _GEN_17444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17685 = _GEN_32732 | _GEN_17445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17686 = _GEN_32733 | _GEN_17446; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17687 = _GEN_32734 | _GEN_17447; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17688 = _GEN_32735 | _GEN_17448; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17689 = _GEN_32736 | _GEN_17449; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17690 = _T_203 ? _GEN_17682 : _GEN_17442; // @[sequencer-master.scala 154:24]
  wire  _GEN_17691 = _T_203 ? _GEN_17683 : _GEN_17443; // @[sequencer-master.scala 154:24]
  wire  _GEN_17692 = _T_203 ? _GEN_17684 : _GEN_17444; // @[sequencer-master.scala 154:24]
  wire  _GEN_17693 = _T_203 ? _GEN_17685 : _GEN_17445; // @[sequencer-master.scala 154:24]
  wire  _GEN_17694 = _T_203 ? _GEN_17686 : _GEN_17446; // @[sequencer-master.scala 154:24]
  wire  _GEN_17695 = _T_203 ? _GEN_17687 : _GEN_17447; // @[sequencer-master.scala 154:24]
  wire  _GEN_17696 = _T_203 ? _GEN_17688 : _GEN_17448; // @[sequencer-master.scala 154:24]
  wire  _GEN_17697 = _T_203 ? _GEN_17689 : _GEN_17449; // @[sequencer-master.scala 154:24]
  wire  _GEN_17698 = _GEN_32729 | _GEN_17458; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17699 = _GEN_32730 | _GEN_17459; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17700 = _GEN_32731 | _GEN_17460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17701 = _GEN_32732 | _GEN_17461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17702 = _GEN_32733 | _GEN_17462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17703 = _GEN_32734 | _GEN_17463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17704 = _GEN_32735 | _GEN_17464; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17705 = _GEN_32736 | _GEN_17465; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17706 = _T_225 ? _GEN_17698 : _GEN_17458; // @[sequencer-master.scala 154:24]
  wire  _GEN_17707 = _T_225 ? _GEN_17699 : _GEN_17459; // @[sequencer-master.scala 154:24]
  wire  _GEN_17708 = _T_225 ? _GEN_17700 : _GEN_17460; // @[sequencer-master.scala 154:24]
  wire  _GEN_17709 = _T_225 ? _GEN_17701 : _GEN_17461; // @[sequencer-master.scala 154:24]
  wire  _GEN_17710 = _T_225 ? _GEN_17702 : _GEN_17462; // @[sequencer-master.scala 154:24]
  wire  _GEN_17711 = _T_225 ? _GEN_17703 : _GEN_17463; // @[sequencer-master.scala 154:24]
  wire  _GEN_17712 = _T_225 ? _GEN_17704 : _GEN_17464; // @[sequencer-master.scala 154:24]
  wire  _GEN_17713 = _T_225 ? _GEN_17705 : _GEN_17465; // @[sequencer-master.scala 154:24]
  wire  _GEN_17714 = _GEN_32729 | _GEN_17474; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17715 = _GEN_32730 | _GEN_17475; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17716 = _GEN_32731 | _GEN_17476; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17717 = _GEN_32732 | _GEN_17477; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17718 = _GEN_32733 | _GEN_17478; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17719 = _GEN_32734 | _GEN_17479; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17720 = _GEN_32735 | _GEN_17480; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17721 = _GEN_32736 | _GEN_17481; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17722 = _T_247 ? _GEN_17714 : _GEN_17474; // @[sequencer-master.scala 154:24]
  wire  _GEN_17723 = _T_247 ? _GEN_17715 : _GEN_17475; // @[sequencer-master.scala 154:24]
  wire  _GEN_17724 = _T_247 ? _GEN_17716 : _GEN_17476; // @[sequencer-master.scala 154:24]
  wire  _GEN_17725 = _T_247 ? _GEN_17717 : _GEN_17477; // @[sequencer-master.scala 154:24]
  wire  _GEN_17726 = _T_247 ? _GEN_17718 : _GEN_17478; // @[sequencer-master.scala 154:24]
  wire  _GEN_17727 = _T_247 ? _GEN_17719 : _GEN_17479; // @[sequencer-master.scala 154:24]
  wire  _GEN_17728 = _T_247 ? _GEN_17720 : _GEN_17480; // @[sequencer-master.scala 154:24]
  wire  _GEN_17729 = _T_247 ? _GEN_17721 : _GEN_17481; // @[sequencer-master.scala 154:24]
  wire  _GEN_17730 = _GEN_32729 | _GEN_17490; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17731 = _GEN_32730 | _GEN_17491; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17732 = _GEN_32731 | _GEN_17492; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17733 = _GEN_32732 | _GEN_17493; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17734 = _GEN_32733 | _GEN_17494; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17735 = _GEN_32734 | _GEN_17495; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17736 = _GEN_32735 | _GEN_17496; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17737 = _GEN_32736 | _GEN_17497; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17738 = _T_269 ? _GEN_17730 : _GEN_17490; // @[sequencer-master.scala 154:24]
  wire  _GEN_17739 = _T_269 ? _GEN_17731 : _GEN_17491; // @[sequencer-master.scala 154:24]
  wire  _GEN_17740 = _T_269 ? _GEN_17732 : _GEN_17492; // @[sequencer-master.scala 154:24]
  wire  _GEN_17741 = _T_269 ? _GEN_17733 : _GEN_17493; // @[sequencer-master.scala 154:24]
  wire  _GEN_17742 = _T_269 ? _GEN_17734 : _GEN_17494; // @[sequencer-master.scala 154:24]
  wire  _GEN_17743 = _T_269 ? _GEN_17735 : _GEN_17495; // @[sequencer-master.scala 154:24]
  wire  _GEN_17744 = _T_269 ? _GEN_17736 : _GEN_17496; // @[sequencer-master.scala 154:24]
  wire  _GEN_17745 = _T_269 ? _GEN_17737 : _GEN_17497; // @[sequencer-master.scala 154:24]
  wire  _GEN_17746 = _GEN_32729 | _GEN_17506; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17747 = _GEN_32730 | _GEN_17507; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17748 = _GEN_32731 | _GEN_17508; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17749 = _GEN_32732 | _GEN_17509; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17750 = _GEN_32733 | _GEN_17510; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17751 = _GEN_32734 | _GEN_17511; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17752 = _GEN_32735 | _GEN_17512; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17753 = _GEN_32736 | _GEN_17513; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17754 = _T_291 ? _GEN_17746 : _GEN_17506; // @[sequencer-master.scala 154:24]
  wire  _GEN_17755 = _T_291 ? _GEN_17747 : _GEN_17507; // @[sequencer-master.scala 154:24]
  wire  _GEN_17756 = _T_291 ? _GEN_17748 : _GEN_17508; // @[sequencer-master.scala 154:24]
  wire  _GEN_17757 = _T_291 ? _GEN_17749 : _GEN_17509; // @[sequencer-master.scala 154:24]
  wire  _GEN_17758 = _T_291 ? _GEN_17750 : _GEN_17510; // @[sequencer-master.scala 154:24]
  wire  _GEN_17759 = _T_291 ? _GEN_17751 : _GEN_17511; // @[sequencer-master.scala 154:24]
  wire  _GEN_17760 = _T_291 ? _GEN_17752 : _GEN_17512; // @[sequencer-master.scala 154:24]
  wire  _GEN_17761 = _T_291 ? _GEN_17753 : _GEN_17513; // @[sequencer-master.scala 154:24]
  wire  _GEN_17762 = _GEN_32729 | _GEN_17522; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17763 = _GEN_32730 | _GEN_17523; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17764 = _GEN_32731 | _GEN_17524; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17765 = _GEN_32732 | _GEN_17525; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17766 = _GEN_32733 | _GEN_17526; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17767 = _GEN_32734 | _GEN_17527; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17768 = _GEN_32735 | _GEN_17528; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17769 = _GEN_32736 | _GEN_17529; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17770 = _T_313 ? _GEN_17762 : _GEN_17522; // @[sequencer-master.scala 154:24]
  wire  _GEN_17771 = _T_313 ? _GEN_17763 : _GEN_17523; // @[sequencer-master.scala 154:24]
  wire  _GEN_17772 = _T_313 ? _GEN_17764 : _GEN_17524; // @[sequencer-master.scala 154:24]
  wire  _GEN_17773 = _T_313 ? _GEN_17765 : _GEN_17525; // @[sequencer-master.scala 154:24]
  wire  _GEN_17774 = _T_313 ? _GEN_17766 : _GEN_17526; // @[sequencer-master.scala 154:24]
  wire  _GEN_17775 = _T_313 ? _GEN_17767 : _GEN_17527; // @[sequencer-master.scala 154:24]
  wire  _GEN_17776 = _T_313 ? _GEN_17768 : _GEN_17528; // @[sequencer-master.scala 154:24]
  wire  _GEN_17777 = _T_313 ? _GEN_17769 : _GEN_17529; // @[sequencer-master.scala 154:24]
  wire  _GEN_17778 = _GEN_32729 | _GEN_17538; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17779 = _GEN_32730 | _GEN_17539; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17780 = _GEN_32731 | _GEN_17540; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17781 = _GEN_32732 | _GEN_17541; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17782 = _GEN_32733 | _GEN_17542; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17783 = _GEN_32734 | _GEN_17543; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17784 = _GEN_32735 | _GEN_17544; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17785 = _GEN_32736 | _GEN_17545; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17786 = _T_335 ? _GEN_17778 : _GEN_17538; // @[sequencer-master.scala 154:24]
  wire  _GEN_17787 = _T_335 ? _GEN_17779 : _GEN_17539; // @[sequencer-master.scala 154:24]
  wire  _GEN_17788 = _T_335 ? _GEN_17780 : _GEN_17540; // @[sequencer-master.scala 154:24]
  wire  _GEN_17789 = _T_335 ? _GEN_17781 : _GEN_17541; // @[sequencer-master.scala 154:24]
  wire  _GEN_17790 = _T_335 ? _GEN_17782 : _GEN_17542; // @[sequencer-master.scala 154:24]
  wire  _GEN_17791 = _T_335 ? _GEN_17783 : _GEN_17543; // @[sequencer-master.scala 154:24]
  wire  _GEN_17792 = _T_335 ? _GEN_17784 : _GEN_17544; // @[sequencer-master.scala 154:24]
  wire  _GEN_17793 = _T_335 ? _GEN_17785 : _GEN_17545; // @[sequencer-master.scala 154:24]
  wire  _GEN_17794 = _GEN_32729 | _GEN_17554; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17795 = _GEN_32730 | _GEN_17555; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17796 = _GEN_32731 | _GEN_17556; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17797 = _GEN_32732 | _GEN_17557; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17798 = _GEN_32733 | _GEN_17558; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17799 = _GEN_32734 | _GEN_17559; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17800 = _GEN_32735 | _GEN_17560; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17801 = _GEN_32736 | _GEN_17561; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_17802 = _T_357 ? _GEN_17794 : _GEN_17554; // @[sequencer-master.scala 154:24]
  wire  _GEN_17803 = _T_357 ? _GEN_17795 : _GEN_17555; // @[sequencer-master.scala 154:24]
  wire  _GEN_17804 = _T_357 ? _GEN_17796 : _GEN_17556; // @[sequencer-master.scala 154:24]
  wire  _GEN_17805 = _T_357 ? _GEN_17797 : _GEN_17557; // @[sequencer-master.scala 154:24]
  wire  _GEN_17806 = _T_357 ? _GEN_17798 : _GEN_17558; // @[sequencer-master.scala 154:24]
  wire  _GEN_17807 = _T_357 ? _GEN_17799 : _GEN_17559; // @[sequencer-master.scala 154:24]
  wire  _GEN_17808 = _T_357 ? _GEN_17800 : _GEN_17560; // @[sequencer-master.scala 154:24]
  wire  _GEN_17809 = _T_357 ? _GEN_17801 : _GEN_17561; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_17810 = 3'h0 == tail ? _T_1615[1:0] : _GEN_17040; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17811 = 3'h1 == tail ? _T_1615[1:0] : _GEN_17041; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17812 = 3'h2 == tail ? _T_1615[1:0] : _GEN_17042; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17813 = 3'h3 == tail ? _T_1615[1:0] : _GEN_17043; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17814 = 3'h4 == tail ? _T_1615[1:0] : _GEN_17044; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17815 = 3'h5 == tail ? _T_1615[1:0] : _GEN_17045; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17816 = 3'h6 == tail ? _T_1615[1:0] : _GEN_17046; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_17817 = 3'h7 == tail ? _T_1615[1:0] : _GEN_17047; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_17818 = 3'h0 == tail ? 4'h0 : _GEN_17048; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17819 = 3'h1 == tail ? 4'h0 : _GEN_17049; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17820 = 3'h2 == tail ? 4'h0 : _GEN_17050; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17821 = 3'h3 == tail ? 4'h0 : _GEN_17051; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17822 = 3'h4 == tail ? 4'h0 : _GEN_17052; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17823 = 3'h5 == tail ? 4'h0 : _GEN_17053; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17824 = 3'h6 == tail ? 4'h0 : _GEN_17054; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_17825 = 3'h7 == tail ? 4'h0 : _GEN_17055; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_17826 = 3'h0 == tail ? 3'h0 : _GEN_17056; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17827 = 3'h1 == tail ? 3'h0 : _GEN_17057; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17828 = 3'h2 == tail ? 3'h0 : _GEN_17058; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17829 = 3'h3 == tail ? 3'h0 : _GEN_17059; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17830 = 3'h4 == tail ? 3'h0 : _GEN_17060; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17831 = 3'h5 == tail ? 3'h0 : _GEN_17061; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17832 = 3'h6 == tail ? 3'h0 : _GEN_17062; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_17833 = 3'h7 == tail ? 3'h0 : _GEN_17063; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_17834 = io_op_bits_active_vrfirst ? _GEN_17066 : _GEN_16720; // @[sequencer-master.scala 649:42]
  wire  _GEN_17835 = io_op_bits_active_vrfirst ? _GEN_17067 : _GEN_16721; // @[sequencer-master.scala 649:42]
  wire  _GEN_17836 = io_op_bits_active_vrfirst ? _GEN_17068 : _GEN_16722; // @[sequencer-master.scala 649:42]
  wire  _GEN_17837 = io_op_bits_active_vrfirst ? _GEN_17069 : _GEN_16723; // @[sequencer-master.scala 649:42]
  wire  _GEN_17838 = io_op_bits_active_vrfirst ? _GEN_17070 : _GEN_16724; // @[sequencer-master.scala 649:42]
  wire  _GEN_17839 = io_op_bits_active_vrfirst ? _GEN_17071 : _GEN_16725; // @[sequencer-master.scala 649:42]
  wire  _GEN_17840 = io_op_bits_active_vrfirst ? _GEN_17072 : _GEN_16726; // @[sequencer-master.scala 649:42]
  wire  _GEN_17841 = io_op_bits_active_vrfirst ? _GEN_17073 : _GEN_16727; // @[sequencer-master.scala 649:42]
  wire  _GEN_17850 = io_op_bits_active_vrfirst ? _GEN_17402 : _GEN_16736; // @[sequencer-master.scala 649:42]
  wire  _GEN_17851 = io_op_bits_active_vrfirst ? _GEN_17403 : _GEN_16737; // @[sequencer-master.scala 649:42]
  wire  _GEN_17852 = io_op_bits_active_vrfirst ? _GEN_17404 : _GEN_16738; // @[sequencer-master.scala 649:42]
  wire  _GEN_17853 = io_op_bits_active_vrfirst ? _GEN_17405 : _GEN_16739; // @[sequencer-master.scala 649:42]
  wire  _GEN_17854 = io_op_bits_active_vrfirst ? _GEN_17406 : _GEN_16740; // @[sequencer-master.scala 649:42]
  wire  _GEN_17855 = io_op_bits_active_vrfirst ? _GEN_17407 : _GEN_16741; // @[sequencer-master.scala 649:42]
  wire  _GEN_17856 = io_op_bits_active_vrfirst ? _GEN_17408 : _GEN_16742; // @[sequencer-master.scala 649:42]
  wire  _GEN_17857 = io_op_bits_active_vrfirst ? _GEN_17409 : _GEN_16743; // @[sequencer-master.scala 649:42]
  wire  _GEN_17858 = io_op_bits_active_vrfirst ? _GEN_17634 : _GEN_16744; // @[sequencer-master.scala 649:42]
  wire  _GEN_17859 = io_op_bits_active_vrfirst ? _GEN_17635 : _GEN_16745; // @[sequencer-master.scala 649:42]
  wire  _GEN_17860 = io_op_bits_active_vrfirst ? _GEN_17636 : _GEN_16746; // @[sequencer-master.scala 649:42]
  wire  _GEN_17861 = io_op_bits_active_vrfirst ? _GEN_17637 : _GEN_16747; // @[sequencer-master.scala 649:42]
  wire  _GEN_17862 = io_op_bits_active_vrfirst ? _GEN_17638 : _GEN_16748; // @[sequencer-master.scala 649:42]
  wire  _GEN_17863 = io_op_bits_active_vrfirst ? _GEN_17639 : _GEN_16749; // @[sequencer-master.scala 649:42]
  wire  _GEN_17864 = io_op_bits_active_vrfirst ? _GEN_17640 : _GEN_16750; // @[sequencer-master.scala 649:42]
  wire  _GEN_17865 = io_op_bits_active_vrfirst ? _GEN_17641 : _GEN_16751; // @[sequencer-master.scala 649:42]
  wire  _GEN_17866 = io_op_bits_active_vrfirst ? _GEN_17098 : _GEN_16752; // @[sequencer-master.scala 649:42]
  wire  _GEN_17867 = io_op_bits_active_vrfirst ? _GEN_17099 : _GEN_16753; // @[sequencer-master.scala 649:42]
  wire  _GEN_17868 = io_op_bits_active_vrfirst ? _GEN_17100 : _GEN_16754; // @[sequencer-master.scala 649:42]
  wire  _GEN_17869 = io_op_bits_active_vrfirst ? _GEN_17101 : _GEN_16755; // @[sequencer-master.scala 649:42]
  wire  _GEN_17870 = io_op_bits_active_vrfirst ? _GEN_17102 : _GEN_16756; // @[sequencer-master.scala 649:42]
  wire  _GEN_17871 = io_op_bits_active_vrfirst ? _GEN_17103 : _GEN_16757; // @[sequencer-master.scala 649:42]
  wire  _GEN_17872 = io_op_bits_active_vrfirst ? _GEN_17104 : _GEN_16758; // @[sequencer-master.scala 649:42]
  wire  _GEN_17873 = io_op_bits_active_vrfirst ? _GEN_17105 : _GEN_16759; // @[sequencer-master.scala 649:42]
  wire  _GEN_17874 = io_op_bits_active_vrfirst ? _GEN_17106 : _GEN_16760; // @[sequencer-master.scala 649:42]
  wire  _GEN_17875 = io_op_bits_active_vrfirst ? _GEN_17107 : _GEN_16761; // @[sequencer-master.scala 649:42]
  wire  _GEN_17876 = io_op_bits_active_vrfirst ? _GEN_17108 : _GEN_16762; // @[sequencer-master.scala 649:42]
  wire  _GEN_17877 = io_op_bits_active_vrfirst ? _GEN_17109 : _GEN_16763; // @[sequencer-master.scala 649:42]
  wire  _GEN_17878 = io_op_bits_active_vrfirst ? _GEN_17110 : _GEN_16764; // @[sequencer-master.scala 649:42]
  wire  _GEN_17879 = io_op_bits_active_vrfirst ? _GEN_17111 : _GEN_16765; // @[sequencer-master.scala 649:42]
  wire  _GEN_17880 = io_op_bits_active_vrfirst ? _GEN_17112 : _GEN_16766; // @[sequencer-master.scala 649:42]
  wire  _GEN_17881 = io_op_bits_active_vrfirst ? _GEN_17113 : _GEN_16767; // @[sequencer-master.scala 649:42]
  wire  _GEN_17882 = io_op_bits_active_vrfirst ? _GEN_17114 : _GEN_16768; // @[sequencer-master.scala 649:42]
  wire  _GEN_17883 = io_op_bits_active_vrfirst ? _GEN_17115 : _GEN_16769; // @[sequencer-master.scala 649:42]
  wire  _GEN_17884 = io_op_bits_active_vrfirst ? _GEN_17116 : _GEN_16770; // @[sequencer-master.scala 649:42]
  wire  _GEN_17885 = io_op_bits_active_vrfirst ? _GEN_17117 : _GEN_16771; // @[sequencer-master.scala 649:42]
  wire  _GEN_17886 = io_op_bits_active_vrfirst ? _GEN_17118 : _GEN_16772; // @[sequencer-master.scala 649:42]
  wire  _GEN_17887 = io_op_bits_active_vrfirst ? _GEN_17119 : _GEN_16773; // @[sequencer-master.scala 649:42]
  wire  _GEN_17888 = io_op_bits_active_vrfirst ? _GEN_17120 : _GEN_16774; // @[sequencer-master.scala 649:42]
  wire  _GEN_17889 = io_op_bits_active_vrfirst ? _GEN_17121 : _GEN_16775; // @[sequencer-master.scala 649:42]
  wire  _GEN_17890 = io_op_bits_active_vrfirst ? _GEN_17122 : _GEN_16776; // @[sequencer-master.scala 649:42]
  wire  _GEN_17891 = io_op_bits_active_vrfirst ? _GEN_17123 : _GEN_16777; // @[sequencer-master.scala 649:42]
  wire  _GEN_17892 = io_op_bits_active_vrfirst ? _GEN_17124 : _GEN_16778; // @[sequencer-master.scala 649:42]
  wire  _GEN_17893 = io_op_bits_active_vrfirst ? _GEN_17125 : _GEN_16779; // @[sequencer-master.scala 649:42]
  wire  _GEN_17894 = io_op_bits_active_vrfirst ? _GEN_17126 : _GEN_16780; // @[sequencer-master.scala 649:42]
  wire  _GEN_17895 = io_op_bits_active_vrfirst ? _GEN_17127 : _GEN_16781; // @[sequencer-master.scala 649:42]
  wire  _GEN_17896 = io_op_bits_active_vrfirst ? _GEN_17128 : _GEN_16782; // @[sequencer-master.scala 649:42]
  wire  _GEN_17897 = io_op_bits_active_vrfirst ? _GEN_17129 : _GEN_16783; // @[sequencer-master.scala 649:42]
  wire  _GEN_17898 = io_op_bits_active_vrfirst ? _GEN_17690 : _GEN_16784; // @[sequencer-master.scala 649:42]
  wire  _GEN_17899 = io_op_bits_active_vrfirst ? _GEN_17691 : _GEN_16785; // @[sequencer-master.scala 649:42]
  wire  _GEN_17900 = io_op_bits_active_vrfirst ? _GEN_17692 : _GEN_16786; // @[sequencer-master.scala 649:42]
  wire  _GEN_17901 = io_op_bits_active_vrfirst ? _GEN_17693 : _GEN_16787; // @[sequencer-master.scala 649:42]
  wire  _GEN_17902 = io_op_bits_active_vrfirst ? _GEN_17694 : _GEN_16788; // @[sequencer-master.scala 649:42]
  wire  _GEN_17903 = io_op_bits_active_vrfirst ? _GEN_17695 : _GEN_16789; // @[sequencer-master.scala 649:42]
  wire  _GEN_17904 = io_op_bits_active_vrfirst ? _GEN_17696 : _GEN_16790; // @[sequencer-master.scala 649:42]
  wire  _GEN_17905 = io_op_bits_active_vrfirst ? _GEN_17697 : _GEN_16791; // @[sequencer-master.scala 649:42]
  wire  _GEN_17906 = io_op_bits_active_vrfirst ? _GEN_17138 : _GEN_16792; // @[sequencer-master.scala 649:42]
  wire  _GEN_17907 = io_op_bits_active_vrfirst ? _GEN_17139 : _GEN_16793; // @[sequencer-master.scala 649:42]
  wire  _GEN_17908 = io_op_bits_active_vrfirst ? _GEN_17140 : _GEN_16794; // @[sequencer-master.scala 649:42]
  wire  _GEN_17909 = io_op_bits_active_vrfirst ? _GEN_17141 : _GEN_16795; // @[sequencer-master.scala 649:42]
  wire  _GEN_17910 = io_op_bits_active_vrfirst ? _GEN_17142 : _GEN_16796; // @[sequencer-master.scala 649:42]
  wire  _GEN_17911 = io_op_bits_active_vrfirst ? _GEN_17143 : _GEN_16797; // @[sequencer-master.scala 649:42]
  wire  _GEN_17912 = io_op_bits_active_vrfirst ? _GEN_17144 : _GEN_16798; // @[sequencer-master.scala 649:42]
  wire  _GEN_17913 = io_op_bits_active_vrfirst ? _GEN_17145 : _GEN_16799; // @[sequencer-master.scala 649:42]
  wire  _GEN_17914 = io_op_bits_active_vrfirst ? _GEN_17146 : _GEN_16800; // @[sequencer-master.scala 649:42]
  wire  _GEN_17915 = io_op_bits_active_vrfirst ? _GEN_17147 : _GEN_16801; // @[sequencer-master.scala 649:42]
  wire  _GEN_17916 = io_op_bits_active_vrfirst ? _GEN_17148 : _GEN_16802; // @[sequencer-master.scala 649:42]
  wire  _GEN_17917 = io_op_bits_active_vrfirst ? _GEN_17149 : _GEN_16803; // @[sequencer-master.scala 649:42]
  wire  _GEN_17918 = io_op_bits_active_vrfirst ? _GEN_17150 : _GEN_16804; // @[sequencer-master.scala 649:42]
  wire  _GEN_17919 = io_op_bits_active_vrfirst ? _GEN_17151 : _GEN_16805; // @[sequencer-master.scala 649:42]
  wire  _GEN_17920 = io_op_bits_active_vrfirst ? _GEN_17152 : _GEN_16806; // @[sequencer-master.scala 649:42]
  wire  _GEN_17921 = io_op_bits_active_vrfirst ? _GEN_17153 : _GEN_16807; // @[sequencer-master.scala 649:42]
  wire  _GEN_17922 = io_op_bits_active_vrfirst ? _GEN_17706 : _GEN_16808; // @[sequencer-master.scala 649:42]
  wire  _GEN_17923 = io_op_bits_active_vrfirst ? _GEN_17707 : _GEN_16809; // @[sequencer-master.scala 649:42]
  wire  _GEN_17924 = io_op_bits_active_vrfirst ? _GEN_17708 : _GEN_16810; // @[sequencer-master.scala 649:42]
  wire  _GEN_17925 = io_op_bits_active_vrfirst ? _GEN_17709 : _GEN_16811; // @[sequencer-master.scala 649:42]
  wire  _GEN_17926 = io_op_bits_active_vrfirst ? _GEN_17710 : _GEN_16812; // @[sequencer-master.scala 649:42]
  wire  _GEN_17927 = io_op_bits_active_vrfirst ? _GEN_17711 : _GEN_16813; // @[sequencer-master.scala 649:42]
  wire  _GEN_17928 = io_op_bits_active_vrfirst ? _GEN_17712 : _GEN_16814; // @[sequencer-master.scala 649:42]
  wire  _GEN_17929 = io_op_bits_active_vrfirst ? _GEN_17713 : _GEN_16815; // @[sequencer-master.scala 649:42]
  wire  _GEN_17930 = io_op_bits_active_vrfirst ? _GEN_17162 : _GEN_16816; // @[sequencer-master.scala 649:42]
  wire  _GEN_17931 = io_op_bits_active_vrfirst ? _GEN_17163 : _GEN_16817; // @[sequencer-master.scala 649:42]
  wire  _GEN_17932 = io_op_bits_active_vrfirst ? _GEN_17164 : _GEN_16818; // @[sequencer-master.scala 649:42]
  wire  _GEN_17933 = io_op_bits_active_vrfirst ? _GEN_17165 : _GEN_16819; // @[sequencer-master.scala 649:42]
  wire  _GEN_17934 = io_op_bits_active_vrfirst ? _GEN_17166 : _GEN_16820; // @[sequencer-master.scala 649:42]
  wire  _GEN_17935 = io_op_bits_active_vrfirst ? _GEN_17167 : _GEN_16821; // @[sequencer-master.scala 649:42]
  wire  _GEN_17936 = io_op_bits_active_vrfirst ? _GEN_17168 : _GEN_16822; // @[sequencer-master.scala 649:42]
  wire  _GEN_17937 = io_op_bits_active_vrfirst ? _GEN_17169 : _GEN_16823; // @[sequencer-master.scala 649:42]
  wire  _GEN_17938 = io_op_bits_active_vrfirst ? _GEN_17170 : _GEN_16824; // @[sequencer-master.scala 649:42]
  wire  _GEN_17939 = io_op_bits_active_vrfirst ? _GEN_17171 : _GEN_16825; // @[sequencer-master.scala 649:42]
  wire  _GEN_17940 = io_op_bits_active_vrfirst ? _GEN_17172 : _GEN_16826; // @[sequencer-master.scala 649:42]
  wire  _GEN_17941 = io_op_bits_active_vrfirst ? _GEN_17173 : _GEN_16827; // @[sequencer-master.scala 649:42]
  wire  _GEN_17942 = io_op_bits_active_vrfirst ? _GEN_17174 : _GEN_16828; // @[sequencer-master.scala 649:42]
  wire  _GEN_17943 = io_op_bits_active_vrfirst ? _GEN_17175 : _GEN_16829; // @[sequencer-master.scala 649:42]
  wire  _GEN_17944 = io_op_bits_active_vrfirst ? _GEN_17176 : _GEN_16830; // @[sequencer-master.scala 649:42]
  wire  _GEN_17945 = io_op_bits_active_vrfirst ? _GEN_17177 : _GEN_16831; // @[sequencer-master.scala 649:42]
  wire  _GEN_17946 = io_op_bits_active_vrfirst ? _GEN_17722 : _GEN_16832; // @[sequencer-master.scala 649:42]
  wire  _GEN_17947 = io_op_bits_active_vrfirst ? _GEN_17723 : _GEN_16833; // @[sequencer-master.scala 649:42]
  wire  _GEN_17948 = io_op_bits_active_vrfirst ? _GEN_17724 : _GEN_16834; // @[sequencer-master.scala 649:42]
  wire  _GEN_17949 = io_op_bits_active_vrfirst ? _GEN_17725 : _GEN_16835; // @[sequencer-master.scala 649:42]
  wire  _GEN_17950 = io_op_bits_active_vrfirst ? _GEN_17726 : _GEN_16836; // @[sequencer-master.scala 649:42]
  wire  _GEN_17951 = io_op_bits_active_vrfirst ? _GEN_17727 : _GEN_16837; // @[sequencer-master.scala 649:42]
  wire  _GEN_17952 = io_op_bits_active_vrfirst ? _GEN_17728 : _GEN_16838; // @[sequencer-master.scala 649:42]
  wire  _GEN_17953 = io_op_bits_active_vrfirst ? _GEN_17729 : _GEN_16839; // @[sequencer-master.scala 649:42]
  wire  _GEN_17954 = io_op_bits_active_vrfirst ? _GEN_17186 : _GEN_16840; // @[sequencer-master.scala 649:42]
  wire  _GEN_17955 = io_op_bits_active_vrfirst ? _GEN_17187 : _GEN_16841; // @[sequencer-master.scala 649:42]
  wire  _GEN_17956 = io_op_bits_active_vrfirst ? _GEN_17188 : _GEN_16842; // @[sequencer-master.scala 649:42]
  wire  _GEN_17957 = io_op_bits_active_vrfirst ? _GEN_17189 : _GEN_16843; // @[sequencer-master.scala 649:42]
  wire  _GEN_17958 = io_op_bits_active_vrfirst ? _GEN_17190 : _GEN_16844; // @[sequencer-master.scala 649:42]
  wire  _GEN_17959 = io_op_bits_active_vrfirst ? _GEN_17191 : _GEN_16845; // @[sequencer-master.scala 649:42]
  wire  _GEN_17960 = io_op_bits_active_vrfirst ? _GEN_17192 : _GEN_16846; // @[sequencer-master.scala 649:42]
  wire  _GEN_17961 = io_op_bits_active_vrfirst ? _GEN_17193 : _GEN_16847; // @[sequencer-master.scala 649:42]
  wire  _GEN_17962 = io_op_bits_active_vrfirst ? _GEN_17194 : _GEN_16848; // @[sequencer-master.scala 649:42]
  wire  _GEN_17963 = io_op_bits_active_vrfirst ? _GEN_17195 : _GEN_16849; // @[sequencer-master.scala 649:42]
  wire  _GEN_17964 = io_op_bits_active_vrfirst ? _GEN_17196 : _GEN_16850; // @[sequencer-master.scala 649:42]
  wire  _GEN_17965 = io_op_bits_active_vrfirst ? _GEN_17197 : _GEN_16851; // @[sequencer-master.scala 649:42]
  wire  _GEN_17966 = io_op_bits_active_vrfirst ? _GEN_17198 : _GEN_16852; // @[sequencer-master.scala 649:42]
  wire  _GEN_17967 = io_op_bits_active_vrfirst ? _GEN_17199 : _GEN_16853; // @[sequencer-master.scala 649:42]
  wire  _GEN_17968 = io_op_bits_active_vrfirst ? _GEN_17200 : _GEN_16854; // @[sequencer-master.scala 649:42]
  wire  _GEN_17969 = io_op_bits_active_vrfirst ? _GEN_17201 : _GEN_16855; // @[sequencer-master.scala 649:42]
  wire  _GEN_17970 = io_op_bits_active_vrfirst ? _GEN_17738 : _GEN_16856; // @[sequencer-master.scala 649:42]
  wire  _GEN_17971 = io_op_bits_active_vrfirst ? _GEN_17739 : _GEN_16857; // @[sequencer-master.scala 649:42]
  wire  _GEN_17972 = io_op_bits_active_vrfirst ? _GEN_17740 : _GEN_16858; // @[sequencer-master.scala 649:42]
  wire  _GEN_17973 = io_op_bits_active_vrfirst ? _GEN_17741 : _GEN_16859; // @[sequencer-master.scala 649:42]
  wire  _GEN_17974 = io_op_bits_active_vrfirst ? _GEN_17742 : _GEN_16860; // @[sequencer-master.scala 649:42]
  wire  _GEN_17975 = io_op_bits_active_vrfirst ? _GEN_17743 : _GEN_16861; // @[sequencer-master.scala 649:42]
  wire  _GEN_17976 = io_op_bits_active_vrfirst ? _GEN_17744 : _GEN_16862; // @[sequencer-master.scala 649:42]
  wire  _GEN_17977 = io_op_bits_active_vrfirst ? _GEN_17745 : _GEN_16863; // @[sequencer-master.scala 649:42]
  wire  _GEN_17978 = io_op_bits_active_vrfirst ? _GEN_17210 : _GEN_16864; // @[sequencer-master.scala 649:42]
  wire  _GEN_17979 = io_op_bits_active_vrfirst ? _GEN_17211 : _GEN_16865; // @[sequencer-master.scala 649:42]
  wire  _GEN_17980 = io_op_bits_active_vrfirst ? _GEN_17212 : _GEN_16866; // @[sequencer-master.scala 649:42]
  wire  _GEN_17981 = io_op_bits_active_vrfirst ? _GEN_17213 : _GEN_16867; // @[sequencer-master.scala 649:42]
  wire  _GEN_17982 = io_op_bits_active_vrfirst ? _GEN_17214 : _GEN_16868; // @[sequencer-master.scala 649:42]
  wire  _GEN_17983 = io_op_bits_active_vrfirst ? _GEN_17215 : _GEN_16869; // @[sequencer-master.scala 649:42]
  wire  _GEN_17984 = io_op_bits_active_vrfirst ? _GEN_17216 : _GEN_16870; // @[sequencer-master.scala 649:42]
  wire  _GEN_17985 = io_op_bits_active_vrfirst ? _GEN_17217 : _GEN_16871; // @[sequencer-master.scala 649:42]
  wire  _GEN_17986 = io_op_bits_active_vrfirst ? _GEN_17218 : _GEN_16872; // @[sequencer-master.scala 649:42]
  wire  _GEN_17987 = io_op_bits_active_vrfirst ? _GEN_17219 : _GEN_16873; // @[sequencer-master.scala 649:42]
  wire  _GEN_17988 = io_op_bits_active_vrfirst ? _GEN_17220 : _GEN_16874; // @[sequencer-master.scala 649:42]
  wire  _GEN_17989 = io_op_bits_active_vrfirst ? _GEN_17221 : _GEN_16875; // @[sequencer-master.scala 649:42]
  wire  _GEN_17990 = io_op_bits_active_vrfirst ? _GEN_17222 : _GEN_16876; // @[sequencer-master.scala 649:42]
  wire  _GEN_17991 = io_op_bits_active_vrfirst ? _GEN_17223 : _GEN_16877; // @[sequencer-master.scala 649:42]
  wire  _GEN_17992 = io_op_bits_active_vrfirst ? _GEN_17224 : _GEN_16878; // @[sequencer-master.scala 649:42]
  wire  _GEN_17993 = io_op_bits_active_vrfirst ? _GEN_17225 : _GEN_16879; // @[sequencer-master.scala 649:42]
  wire  _GEN_17994 = io_op_bits_active_vrfirst ? _GEN_17754 : _GEN_16880; // @[sequencer-master.scala 649:42]
  wire  _GEN_17995 = io_op_bits_active_vrfirst ? _GEN_17755 : _GEN_16881; // @[sequencer-master.scala 649:42]
  wire  _GEN_17996 = io_op_bits_active_vrfirst ? _GEN_17756 : _GEN_16882; // @[sequencer-master.scala 649:42]
  wire  _GEN_17997 = io_op_bits_active_vrfirst ? _GEN_17757 : _GEN_16883; // @[sequencer-master.scala 649:42]
  wire  _GEN_17998 = io_op_bits_active_vrfirst ? _GEN_17758 : _GEN_16884; // @[sequencer-master.scala 649:42]
  wire  _GEN_17999 = io_op_bits_active_vrfirst ? _GEN_17759 : _GEN_16885; // @[sequencer-master.scala 649:42]
  wire  _GEN_18000 = io_op_bits_active_vrfirst ? _GEN_17760 : _GEN_16886; // @[sequencer-master.scala 649:42]
  wire  _GEN_18001 = io_op_bits_active_vrfirst ? _GEN_17761 : _GEN_16887; // @[sequencer-master.scala 649:42]
  wire  _GEN_18002 = io_op_bits_active_vrfirst ? _GEN_17234 : _GEN_16888; // @[sequencer-master.scala 649:42]
  wire  _GEN_18003 = io_op_bits_active_vrfirst ? _GEN_17235 : _GEN_16889; // @[sequencer-master.scala 649:42]
  wire  _GEN_18004 = io_op_bits_active_vrfirst ? _GEN_17236 : _GEN_16890; // @[sequencer-master.scala 649:42]
  wire  _GEN_18005 = io_op_bits_active_vrfirst ? _GEN_17237 : _GEN_16891; // @[sequencer-master.scala 649:42]
  wire  _GEN_18006 = io_op_bits_active_vrfirst ? _GEN_17238 : _GEN_16892; // @[sequencer-master.scala 649:42]
  wire  _GEN_18007 = io_op_bits_active_vrfirst ? _GEN_17239 : _GEN_16893; // @[sequencer-master.scala 649:42]
  wire  _GEN_18008 = io_op_bits_active_vrfirst ? _GEN_17240 : _GEN_16894; // @[sequencer-master.scala 649:42]
  wire  _GEN_18009 = io_op_bits_active_vrfirst ? _GEN_17241 : _GEN_16895; // @[sequencer-master.scala 649:42]
  wire  _GEN_18010 = io_op_bits_active_vrfirst ? _GEN_17242 : _GEN_16896; // @[sequencer-master.scala 649:42]
  wire  _GEN_18011 = io_op_bits_active_vrfirst ? _GEN_17243 : _GEN_16897; // @[sequencer-master.scala 649:42]
  wire  _GEN_18012 = io_op_bits_active_vrfirst ? _GEN_17244 : _GEN_16898; // @[sequencer-master.scala 649:42]
  wire  _GEN_18013 = io_op_bits_active_vrfirst ? _GEN_17245 : _GEN_16899; // @[sequencer-master.scala 649:42]
  wire  _GEN_18014 = io_op_bits_active_vrfirst ? _GEN_17246 : _GEN_16900; // @[sequencer-master.scala 649:42]
  wire  _GEN_18015 = io_op_bits_active_vrfirst ? _GEN_17247 : _GEN_16901; // @[sequencer-master.scala 649:42]
  wire  _GEN_18016 = io_op_bits_active_vrfirst ? _GEN_17248 : _GEN_16902; // @[sequencer-master.scala 649:42]
  wire  _GEN_18017 = io_op_bits_active_vrfirst ? _GEN_17249 : _GEN_16903; // @[sequencer-master.scala 649:42]
  wire  _GEN_18018 = io_op_bits_active_vrfirst ? _GEN_17770 : _GEN_16904; // @[sequencer-master.scala 649:42]
  wire  _GEN_18019 = io_op_bits_active_vrfirst ? _GEN_17771 : _GEN_16905; // @[sequencer-master.scala 649:42]
  wire  _GEN_18020 = io_op_bits_active_vrfirst ? _GEN_17772 : _GEN_16906; // @[sequencer-master.scala 649:42]
  wire  _GEN_18021 = io_op_bits_active_vrfirst ? _GEN_17773 : _GEN_16907; // @[sequencer-master.scala 649:42]
  wire  _GEN_18022 = io_op_bits_active_vrfirst ? _GEN_17774 : _GEN_16908; // @[sequencer-master.scala 649:42]
  wire  _GEN_18023 = io_op_bits_active_vrfirst ? _GEN_17775 : _GEN_16909; // @[sequencer-master.scala 649:42]
  wire  _GEN_18024 = io_op_bits_active_vrfirst ? _GEN_17776 : _GEN_16910; // @[sequencer-master.scala 649:42]
  wire  _GEN_18025 = io_op_bits_active_vrfirst ? _GEN_17777 : _GEN_16911; // @[sequencer-master.scala 649:42]
  wire  _GEN_18026 = io_op_bits_active_vrfirst ? _GEN_17258 : _GEN_16912; // @[sequencer-master.scala 649:42]
  wire  _GEN_18027 = io_op_bits_active_vrfirst ? _GEN_17259 : _GEN_16913; // @[sequencer-master.scala 649:42]
  wire  _GEN_18028 = io_op_bits_active_vrfirst ? _GEN_17260 : _GEN_16914; // @[sequencer-master.scala 649:42]
  wire  _GEN_18029 = io_op_bits_active_vrfirst ? _GEN_17261 : _GEN_16915; // @[sequencer-master.scala 649:42]
  wire  _GEN_18030 = io_op_bits_active_vrfirst ? _GEN_17262 : _GEN_16916; // @[sequencer-master.scala 649:42]
  wire  _GEN_18031 = io_op_bits_active_vrfirst ? _GEN_17263 : _GEN_16917; // @[sequencer-master.scala 649:42]
  wire  _GEN_18032 = io_op_bits_active_vrfirst ? _GEN_17264 : _GEN_16918; // @[sequencer-master.scala 649:42]
  wire  _GEN_18033 = io_op_bits_active_vrfirst ? _GEN_17265 : _GEN_16919; // @[sequencer-master.scala 649:42]
  wire  _GEN_18034 = io_op_bits_active_vrfirst ? _GEN_17266 : _GEN_16920; // @[sequencer-master.scala 649:42]
  wire  _GEN_18035 = io_op_bits_active_vrfirst ? _GEN_17267 : _GEN_16921; // @[sequencer-master.scala 649:42]
  wire  _GEN_18036 = io_op_bits_active_vrfirst ? _GEN_17268 : _GEN_16922; // @[sequencer-master.scala 649:42]
  wire  _GEN_18037 = io_op_bits_active_vrfirst ? _GEN_17269 : _GEN_16923; // @[sequencer-master.scala 649:42]
  wire  _GEN_18038 = io_op_bits_active_vrfirst ? _GEN_17270 : _GEN_16924; // @[sequencer-master.scala 649:42]
  wire  _GEN_18039 = io_op_bits_active_vrfirst ? _GEN_17271 : _GEN_16925; // @[sequencer-master.scala 649:42]
  wire  _GEN_18040 = io_op_bits_active_vrfirst ? _GEN_17272 : _GEN_16926; // @[sequencer-master.scala 649:42]
  wire  _GEN_18041 = io_op_bits_active_vrfirst ? _GEN_17273 : _GEN_16927; // @[sequencer-master.scala 649:42]
  wire  _GEN_18042 = io_op_bits_active_vrfirst ? _GEN_17786 : _GEN_16928; // @[sequencer-master.scala 649:42]
  wire  _GEN_18043 = io_op_bits_active_vrfirst ? _GEN_17787 : _GEN_16929; // @[sequencer-master.scala 649:42]
  wire  _GEN_18044 = io_op_bits_active_vrfirst ? _GEN_17788 : _GEN_16930; // @[sequencer-master.scala 649:42]
  wire  _GEN_18045 = io_op_bits_active_vrfirst ? _GEN_17789 : _GEN_16931; // @[sequencer-master.scala 649:42]
  wire  _GEN_18046 = io_op_bits_active_vrfirst ? _GEN_17790 : _GEN_16932; // @[sequencer-master.scala 649:42]
  wire  _GEN_18047 = io_op_bits_active_vrfirst ? _GEN_17791 : _GEN_16933; // @[sequencer-master.scala 649:42]
  wire  _GEN_18048 = io_op_bits_active_vrfirst ? _GEN_17792 : _GEN_16934; // @[sequencer-master.scala 649:42]
  wire  _GEN_18049 = io_op_bits_active_vrfirst ? _GEN_17793 : _GEN_16935; // @[sequencer-master.scala 649:42]
  wire  _GEN_18050 = io_op_bits_active_vrfirst ? _GEN_17282 : _GEN_16936; // @[sequencer-master.scala 649:42]
  wire  _GEN_18051 = io_op_bits_active_vrfirst ? _GEN_17283 : _GEN_16937; // @[sequencer-master.scala 649:42]
  wire  _GEN_18052 = io_op_bits_active_vrfirst ? _GEN_17284 : _GEN_16938; // @[sequencer-master.scala 649:42]
  wire  _GEN_18053 = io_op_bits_active_vrfirst ? _GEN_17285 : _GEN_16939; // @[sequencer-master.scala 649:42]
  wire  _GEN_18054 = io_op_bits_active_vrfirst ? _GEN_17286 : _GEN_16940; // @[sequencer-master.scala 649:42]
  wire  _GEN_18055 = io_op_bits_active_vrfirst ? _GEN_17287 : _GEN_16941; // @[sequencer-master.scala 649:42]
  wire  _GEN_18056 = io_op_bits_active_vrfirst ? _GEN_17288 : _GEN_16942; // @[sequencer-master.scala 649:42]
  wire  _GEN_18057 = io_op_bits_active_vrfirst ? _GEN_17289 : _GEN_16943; // @[sequencer-master.scala 649:42]
  wire  _GEN_18058 = io_op_bits_active_vrfirst ? _GEN_17290 : _GEN_16944; // @[sequencer-master.scala 649:42]
  wire  _GEN_18059 = io_op_bits_active_vrfirst ? _GEN_17291 : _GEN_16945; // @[sequencer-master.scala 649:42]
  wire  _GEN_18060 = io_op_bits_active_vrfirst ? _GEN_17292 : _GEN_16946; // @[sequencer-master.scala 649:42]
  wire  _GEN_18061 = io_op_bits_active_vrfirst ? _GEN_17293 : _GEN_16947; // @[sequencer-master.scala 649:42]
  wire  _GEN_18062 = io_op_bits_active_vrfirst ? _GEN_17294 : _GEN_16948; // @[sequencer-master.scala 649:42]
  wire  _GEN_18063 = io_op_bits_active_vrfirst ? _GEN_17295 : _GEN_16949; // @[sequencer-master.scala 649:42]
  wire  _GEN_18064 = io_op_bits_active_vrfirst ? _GEN_17296 : _GEN_16950; // @[sequencer-master.scala 649:42]
  wire  _GEN_18065 = io_op_bits_active_vrfirst ? _GEN_17297 : _GEN_16951; // @[sequencer-master.scala 649:42]
  wire  _GEN_18066 = io_op_bits_active_vrfirst ? _GEN_17802 : _GEN_16952; // @[sequencer-master.scala 649:42]
  wire  _GEN_18067 = io_op_bits_active_vrfirst ? _GEN_17803 : _GEN_16953; // @[sequencer-master.scala 649:42]
  wire  _GEN_18068 = io_op_bits_active_vrfirst ? _GEN_17804 : _GEN_16954; // @[sequencer-master.scala 649:42]
  wire  _GEN_18069 = io_op_bits_active_vrfirst ? _GEN_17805 : _GEN_16955; // @[sequencer-master.scala 649:42]
  wire  _GEN_18070 = io_op_bits_active_vrfirst ? _GEN_17806 : _GEN_16956; // @[sequencer-master.scala 649:42]
  wire  _GEN_18071 = io_op_bits_active_vrfirst ? _GEN_17807 : _GEN_16957; // @[sequencer-master.scala 649:42]
  wire  _GEN_18072 = io_op_bits_active_vrfirst ? _GEN_17808 : _GEN_16958; // @[sequencer-master.scala 649:42]
  wire  _GEN_18073 = io_op_bits_active_vrfirst ? _GEN_17809 : _GEN_16959; // @[sequencer-master.scala 649:42]
  wire  _GEN_18074 = io_op_bits_active_vrfirst ? _GEN_17306 : _GEN_16960; // @[sequencer-master.scala 649:42]
  wire  _GEN_18075 = io_op_bits_active_vrfirst ? _GEN_17307 : _GEN_16961; // @[sequencer-master.scala 649:42]
  wire  _GEN_18076 = io_op_bits_active_vrfirst ? _GEN_17308 : _GEN_16962; // @[sequencer-master.scala 649:42]
  wire  _GEN_18077 = io_op_bits_active_vrfirst ? _GEN_17309 : _GEN_16963; // @[sequencer-master.scala 649:42]
  wire  _GEN_18078 = io_op_bits_active_vrfirst ? _GEN_17310 : _GEN_16964; // @[sequencer-master.scala 649:42]
  wire  _GEN_18079 = io_op_bits_active_vrfirst ? _GEN_17311 : _GEN_16965; // @[sequencer-master.scala 649:42]
  wire  _GEN_18080 = io_op_bits_active_vrfirst ? _GEN_17312 : _GEN_16966; // @[sequencer-master.scala 649:42]
  wire  _GEN_18081 = io_op_bits_active_vrfirst ? _GEN_17313 : _GEN_16967; // @[sequencer-master.scala 649:42]
  wire  _GEN_18082 = io_op_bits_active_vrfirst ? _GEN_17314 : _GEN_16968; // @[sequencer-master.scala 649:42]
  wire  _GEN_18083 = io_op_bits_active_vrfirst ? _GEN_17315 : _GEN_16969; // @[sequencer-master.scala 649:42]
  wire  _GEN_18084 = io_op_bits_active_vrfirst ? _GEN_17316 : _GEN_16970; // @[sequencer-master.scala 649:42]
  wire  _GEN_18085 = io_op_bits_active_vrfirst ? _GEN_17317 : _GEN_16971; // @[sequencer-master.scala 649:42]
  wire  _GEN_18086 = io_op_bits_active_vrfirst ? _GEN_17318 : _GEN_16972; // @[sequencer-master.scala 649:42]
  wire  _GEN_18087 = io_op_bits_active_vrfirst ? _GEN_17319 : _GEN_16973; // @[sequencer-master.scala 649:42]
  wire  _GEN_18088 = io_op_bits_active_vrfirst ? _GEN_17320 : _GEN_16974; // @[sequencer-master.scala 649:42]
  wire  _GEN_18089 = io_op_bits_active_vrfirst ? _GEN_17321 : _GEN_16975; // @[sequencer-master.scala 649:42]
  wire  _GEN_18090 = io_op_bits_active_vrfirst ? _GEN_17322 : _GEN_16976; // @[sequencer-master.scala 649:42]
  wire  _GEN_18091 = io_op_bits_active_vrfirst ? _GEN_17323 : _GEN_16977; // @[sequencer-master.scala 649:42]
  wire  _GEN_18092 = io_op_bits_active_vrfirst ? _GEN_17324 : _GEN_16978; // @[sequencer-master.scala 649:42]
  wire  _GEN_18093 = io_op_bits_active_vrfirst ? _GEN_17325 : _GEN_16979; // @[sequencer-master.scala 649:42]
  wire  _GEN_18094 = io_op_bits_active_vrfirst ? _GEN_17326 : _GEN_16980; // @[sequencer-master.scala 649:42]
  wire  _GEN_18095 = io_op_bits_active_vrfirst ? _GEN_17327 : _GEN_16981; // @[sequencer-master.scala 649:42]
  wire  _GEN_18096 = io_op_bits_active_vrfirst ? _GEN_17328 : _GEN_16982; // @[sequencer-master.scala 649:42]
  wire  _GEN_18097 = io_op_bits_active_vrfirst ? _GEN_17329 : _GEN_16983; // @[sequencer-master.scala 649:42]
  wire  _GEN_18106 = io_op_bits_active_vrfirst ? _GEN_17338 : _GEN_16992; // @[sequencer-master.scala 649:42]
  wire  _GEN_18107 = io_op_bits_active_vrfirst ? _GEN_17339 : _GEN_16993; // @[sequencer-master.scala 649:42]
  wire  _GEN_18108 = io_op_bits_active_vrfirst ? _GEN_17340 : _GEN_16994; // @[sequencer-master.scala 649:42]
  wire  _GEN_18109 = io_op_bits_active_vrfirst ? _GEN_17341 : _GEN_16995; // @[sequencer-master.scala 649:42]
  wire  _GEN_18110 = io_op_bits_active_vrfirst ? _GEN_17342 : _GEN_16996; // @[sequencer-master.scala 649:42]
  wire  _GEN_18111 = io_op_bits_active_vrfirst ? _GEN_17343 : _GEN_16997; // @[sequencer-master.scala 649:42]
  wire  _GEN_18112 = io_op_bits_active_vrfirst ? _GEN_17344 : _GEN_16998; // @[sequencer-master.scala 649:42]
  wire  _GEN_18113 = io_op_bits_active_vrfirst ? _GEN_17345 : _GEN_16999; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18114 = io_op_bits_active_vrfirst ? _GEN_17346 : _GEN_17000; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18115 = io_op_bits_active_vrfirst ? _GEN_17347 : _GEN_17001; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18116 = io_op_bits_active_vrfirst ? _GEN_17348 : _GEN_17002; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18117 = io_op_bits_active_vrfirst ? _GEN_17349 : _GEN_17003; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18118 = io_op_bits_active_vrfirst ? _GEN_17350 : _GEN_17004; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18119 = io_op_bits_active_vrfirst ? _GEN_17351 : _GEN_17005; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18120 = io_op_bits_active_vrfirst ? _GEN_17352 : _GEN_17006; // @[sequencer-master.scala 649:42]
  wire [9:0] _GEN_18121 = io_op_bits_active_vrfirst ? _GEN_17353 : _GEN_17007; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18122 = io_op_bits_active_vrfirst ? _GEN_17394 : _GEN_17008; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18123 = io_op_bits_active_vrfirst ? _GEN_17395 : _GEN_17009; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18124 = io_op_bits_active_vrfirst ? _GEN_17396 : _GEN_17010; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18125 = io_op_bits_active_vrfirst ? _GEN_17397 : _GEN_17011; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18126 = io_op_bits_active_vrfirst ? _GEN_17398 : _GEN_17012; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18127 = io_op_bits_active_vrfirst ? _GEN_17399 : _GEN_17013; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18128 = io_op_bits_active_vrfirst ? _GEN_17400 : _GEN_17014; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18129 = io_op_bits_active_vrfirst ? _GEN_17401 : _GEN_17015; // @[sequencer-master.scala 649:42]
  wire  _GEN_18130 = io_op_bits_active_vrfirst ? _GEN_17410 : _GEN_17016; // @[sequencer-master.scala 649:42]
  wire  _GEN_18131 = io_op_bits_active_vrfirst ? _GEN_17411 : _GEN_17017; // @[sequencer-master.scala 649:42]
  wire  _GEN_18132 = io_op_bits_active_vrfirst ? _GEN_17412 : _GEN_17018; // @[sequencer-master.scala 649:42]
  wire  _GEN_18133 = io_op_bits_active_vrfirst ? _GEN_17413 : _GEN_17019; // @[sequencer-master.scala 649:42]
  wire  _GEN_18134 = io_op_bits_active_vrfirst ? _GEN_17414 : _GEN_17020; // @[sequencer-master.scala 649:42]
  wire  _GEN_18135 = io_op_bits_active_vrfirst ? _GEN_17415 : _GEN_17021; // @[sequencer-master.scala 649:42]
  wire  _GEN_18136 = io_op_bits_active_vrfirst ? _GEN_17416 : _GEN_17022; // @[sequencer-master.scala 649:42]
  wire  _GEN_18137 = io_op_bits_active_vrfirst ? _GEN_17417 : _GEN_17023; // @[sequencer-master.scala 649:42]
  wire  _GEN_18138 = io_op_bits_active_vrfirst ? _GEN_17418 : _GEN_17024; // @[sequencer-master.scala 649:42]
  wire  _GEN_18139 = io_op_bits_active_vrfirst ? _GEN_17419 : _GEN_17025; // @[sequencer-master.scala 649:42]
  wire  _GEN_18140 = io_op_bits_active_vrfirst ? _GEN_17420 : _GEN_17026; // @[sequencer-master.scala 649:42]
  wire  _GEN_18141 = io_op_bits_active_vrfirst ? _GEN_17421 : _GEN_17027; // @[sequencer-master.scala 649:42]
  wire  _GEN_18142 = io_op_bits_active_vrfirst ? _GEN_17422 : _GEN_17028; // @[sequencer-master.scala 649:42]
  wire  _GEN_18143 = io_op_bits_active_vrfirst ? _GEN_17423 : _GEN_17029; // @[sequencer-master.scala 649:42]
  wire  _GEN_18144 = io_op_bits_active_vrfirst ? _GEN_17424 : _GEN_17030; // @[sequencer-master.scala 649:42]
  wire  _GEN_18145 = io_op_bits_active_vrfirst ? _GEN_17425 : _GEN_17031; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18146 = io_op_bits_active_vrfirst ? _GEN_17426 : _GEN_17032; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18147 = io_op_bits_active_vrfirst ? _GEN_17427 : _GEN_17033; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18148 = io_op_bits_active_vrfirst ? _GEN_17428 : _GEN_17034; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18149 = io_op_bits_active_vrfirst ? _GEN_17429 : _GEN_17035; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18150 = io_op_bits_active_vrfirst ? _GEN_17430 : _GEN_17036; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18151 = io_op_bits_active_vrfirst ? _GEN_17431 : _GEN_17037; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18152 = io_op_bits_active_vrfirst ? _GEN_17432 : _GEN_17038; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18153 = io_op_bits_active_vrfirst ? _GEN_17433 : _GEN_17039; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18154 = io_op_bits_active_vrfirst ? _GEN_17626 : _GEN_16086; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18155 = io_op_bits_active_vrfirst ? _GEN_17627 : _GEN_16087; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18156 = io_op_bits_active_vrfirst ? _GEN_17628 : _GEN_16088; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18157 = io_op_bits_active_vrfirst ? _GEN_17629 : _GEN_16089; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18158 = io_op_bits_active_vrfirst ? _GEN_17630 : _GEN_16090; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18159 = io_op_bits_active_vrfirst ? _GEN_17631 : _GEN_16091; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18160 = io_op_bits_active_vrfirst ? _GEN_17632 : _GEN_16092; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18161 = io_op_bits_active_vrfirst ? _GEN_17633 : _GEN_16093; // @[sequencer-master.scala 649:42]
  wire  _GEN_18162 = io_op_bits_active_vrfirst ? _GEN_17642 : _GEN_16094; // @[sequencer-master.scala 649:42]
  wire  _GEN_18163 = io_op_bits_active_vrfirst ? _GEN_17643 : _GEN_16095; // @[sequencer-master.scala 649:42]
  wire  _GEN_18164 = io_op_bits_active_vrfirst ? _GEN_17644 : _GEN_16096; // @[sequencer-master.scala 649:42]
  wire  _GEN_18165 = io_op_bits_active_vrfirst ? _GEN_17645 : _GEN_16097; // @[sequencer-master.scala 649:42]
  wire  _GEN_18166 = io_op_bits_active_vrfirst ? _GEN_17646 : _GEN_16098; // @[sequencer-master.scala 649:42]
  wire  _GEN_18167 = io_op_bits_active_vrfirst ? _GEN_17647 : _GEN_16099; // @[sequencer-master.scala 649:42]
  wire  _GEN_18168 = io_op_bits_active_vrfirst ? _GEN_17648 : _GEN_16100; // @[sequencer-master.scala 649:42]
  wire  _GEN_18169 = io_op_bits_active_vrfirst ? _GEN_17649 : _GEN_16101; // @[sequencer-master.scala 649:42]
  wire  _GEN_18170 = io_op_bits_active_vrfirst ? _GEN_17650 : _GEN_16102; // @[sequencer-master.scala 649:42]
  wire  _GEN_18171 = io_op_bits_active_vrfirst ? _GEN_17651 : _GEN_16103; // @[sequencer-master.scala 649:42]
  wire  _GEN_18172 = io_op_bits_active_vrfirst ? _GEN_17652 : _GEN_16104; // @[sequencer-master.scala 649:42]
  wire  _GEN_18173 = io_op_bits_active_vrfirst ? _GEN_17653 : _GEN_16105; // @[sequencer-master.scala 649:42]
  wire  _GEN_18174 = io_op_bits_active_vrfirst ? _GEN_17654 : _GEN_16106; // @[sequencer-master.scala 649:42]
  wire  _GEN_18175 = io_op_bits_active_vrfirst ? _GEN_17655 : _GEN_16107; // @[sequencer-master.scala 649:42]
  wire  _GEN_18176 = io_op_bits_active_vrfirst ? _GEN_17656 : _GEN_16108; // @[sequencer-master.scala 649:42]
  wire  _GEN_18177 = io_op_bits_active_vrfirst ? _GEN_17657 : _GEN_16109; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18178 = io_op_bits_active_vrfirst ? _GEN_17658 : _GEN_16110; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18179 = io_op_bits_active_vrfirst ? _GEN_17659 : _GEN_16111; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18180 = io_op_bits_active_vrfirst ? _GEN_17660 : _GEN_16112; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18181 = io_op_bits_active_vrfirst ? _GEN_17661 : _GEN_16113; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18182 = io_op_bits_active_vrfirst ? _GEN_17662 : _GEN_16114; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18183 = io_op_bits_active_vrfirst ? _GEN_17663 : _GEN_16115; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18184 = io_op_bits_active_vrfirst ? _GEN_17664 : _GEN_16116; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18185 = io_op_bits_active_vrfirst ? _GEN_17665 : _GEN_16117; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18186 = io_op_bits_active_vrfirst ? _GEN_17666 : _GEN_16118; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18187 = io_op_bits_active_vrfirst ? _GEN_17667 : _GEN_16119; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18188 = io_op_bits_active_vrfirst ? _GEN_17668 : _GEN_16120; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18189 = io_op_bits_active_vrfirst ? _GEN_17669 : _GEN_16121; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18190 = io_op_bits_active_vrfirst ? _GEN_17670 : _GEN_16122; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18191 = io_op_bits_active_vrfirst ? _GEN_17671 : _GEN_16123; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18192 = io_op_bits_active_vrfirst ? _GEN_17672 : _GEN_16124; // @[sequencer-master.scala 649:42]
  wire [7:0] _GEN_18193 = io_op_bits_active_vrfirst ? _GEN_17673 : _GEN_16125; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18194 = io_op_bits_active_vrfirst ? _GEN_17674 : _GEN_16126; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18195 = io_op_bits_active_vrfirst ? _GEN_17675 : _GEN_16127; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18196 = io_op_bits_active_vrfirst ? _GEN_17676 : _GEN_16128; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18197 = io_op_bits_active_vrfirst ? _GEN_17677 : _GEN_16129; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18198 = io_op_bits_active_vrfirst ? _GEN_17678 : _GEN_16130; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18199 = io_op_bits_active_vrfirst ? _GEN_17679 : _GEN_16131; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18200 = io_op_bits_active_vrfirst ? _GEN_17680 : _GEN_16132; // @[sequencer-master.scala 649:42]
  wire [63:0] _GEN_18201 = io_op_bits_active_vrfirst ? _GEN_17681 : _GEN_16133; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18202 = io_op_bits_active_vrfirst ? _GEN_17810 : _GEN_17040; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18203 = io_op_bits_active_vrfirst ? _GEN_17811 : _GEN_17041; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18204 = io_op_bits_active_vrfirst ? _GEN_17812 : _GEN_17042; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18205 = io_op_bits_active_vrfirst ? _GEN_17813 : _GEN_17043; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18206 = io_op_bits_active_vrfirst ? _GEN_17814 : _GEN_17044; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18207 = io_op_bits_active_vrfirst ? _GEN_17815 : _GEN_17045; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18208 = io_op_bits_active_vrfirst ? _GEN_17816 : _GEN_17046; // @[sequencer-master.scala 649:42]
  wire [1:0] _GEN_18209 = io_op_bits_active_vrfirst ? _GEN_17817 : _GEN_17047; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18210 = io_op_bits_active_vrfirst ? _GEN_17818 : _GEN_17048; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18211 = io_op_bits_active_vrfirst ? _GEN_17819 : _GEN_17049; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18212 = io_op_bits_active_vrfirst ? _GEN_17820 : _GEN_17050; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18213 = io_op_bits_active_vrfirst ? _GEN_17821 : _GEN_17051; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18214 = io_op_bits_active_vrfirst ? _GEN_17822 : _GEN_17052; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18215 = io_op_bits_active_vrfirst ? _GEN_17823 : _GEN_17053; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18216 = io_op_bits_active_vrfirst ? _GEN_17824 : _GEN_17054; // @[sequencer-master.scala 649:42]
  wire [3:0] _GEN_18217 = io_op_bits_active_vrfirst ? _GEN_17825 : _GEN_17055; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18218 = io_op_bits_active_vrfirst ? _GEN_17826 : _GEN_17056; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18219 = io_op_bits_active_vrfirst ? _GEN_17827 : _GEN_17057; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18220 = io_op_bits_active_vrfirst ? _GEN_17828 : _GEN_17058; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18221 = io_op_bits_active_vrfirst ? _GEN_17829 : _GEN_17059; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18222 = io_op_bits_active_vrfirst ? _GEN_17830 : _GEN_17060; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18223 = io_op_bits_active_vrfirst ? _GEN_17831 : _GEN_17061; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18224 = io_op_bits_active_vrfirst ? _GEN_17832 : _GEN_17062; // @[sequencer-master.scala 649:42]
  wire [2:0] _GEN_18225 = io_op_bits_active_vrfirst ? _GEN_17833 : _GEN_17063; // @[sequencer-master.scala 649:42]
  wire  _GEN_18226 = io_op_bits_active_vrfirst | _GEN_17064; // @[sequencer-master.scala 649:42 sequencer-master.scala 265:41]
  wire [2:0] _GEN_18227 = io_op_bits_active_vrfirst ? _T_1645 : _GEN_17065; // @[sequencer-master.scala 649:42 sequencer-master.scala 265:66]
  wire  _GEN_18244 = 3'h0 == tail ? 1'h0 : _GEN_17850; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18245 = 3'h1 == tail ? 1'h0 : _GEN_17851; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18246 = 3'h2 == tail ? 1'h0 : _GEN_17852; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18247 = 3'h3 == tail ? 1'h0 : _GEN_17853; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18248 = 3'h4 == tail ? 1'h0 : _GEN_17854; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18249 = 3'h5 == tail ? 1'h0 : _GEN_17855; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18250 = 3'h6 == tail ? 1'h0 : _GEN_17856; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18251 = 3'h7 == tail ? 1'h0 : _GEN_17857; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_18252 = 3'h0 == tail ? 1'h0 : _GEN_17858; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18253 = 3'h1 == tail ? 1'h0 : _GEN_17859; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18254 = 3'h2 == tail ? 1'h0 : _GEN_17860; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18255 = 3'h3 == tail ? 1'h0 : _GEN_17861; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18256 = 3'h4 == tail ? 1'h0 : _GEN_17862; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18257 = 3'h5 == tail ? 1'h0 : _GEN_17863; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18258 = 3'h6 == tail ? 1'h0 : _GEN_17864; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18259 = 3'h7 == tail ? 1'h0 : _GEN_17865; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_18260 = 3'h0 == tail ? 1'h0 : _GEN_17866; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18261 = 3'h1 == tail ? 1'h0 : _GEN_17867; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18262 = 3'h2 == tail ? 1'h0 : _GEN_17868; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18263 = 3'h3 == tail ? 1'h0 : _GEN_17869; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18264 = 3'h4 == tail ? 1'h0 : _GEN_17870; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18265 = 3'h5 == tail ? 1'h0 : _GEN_17871; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18266 = 3'h6 == tail ? 1'h0 : _GEN_17872; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18267 = 3'h7 == tail ? 1'h0 : _GEN_17873; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_18268 = 3'h0 == tail ? 1'h0 : _GEN_17874; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18269 = 3'h1 == tail ? 1'h0 : _GEN_17875; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18270 = 3'h2 == tail ? 1'h0 : _GEN_17876; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18271 = 3'h3 == tail ? 1'h0 : _GEN_17877; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18272 = 3'h4 == tail ? 1'h0 : _GEN_17878; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18273 = 3'h5 == tail ? 1'h0 : _GEN_17879; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18274 = 3'h6 == tail ? 1'h0 : _GEN_17880; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18275 = 3'h7 == tail ? 1'h0 : _GEN_17881; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_18276 = 3'h0 == tail ? 1'h0 : _GEN_17882; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18277 = 3'h1 == tail ? 1'h0 : _GEN_17883; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18278 = 3'h2 == tail ? 1'h0 : _GEN_17884; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18279 = 3'h3 == tail ? 1'h0 : _GEN_17885; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18280 = 3'h4 == tail ? 1'h0 : _GEN_17886; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18281 = 3'h5 == tail ? 1'h0 : _GEN_17887; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18282 = 3'h6 == tail ? 1'h0 : _GEN_17888; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18283 = 3'h7 == tail ? 1'h0 : _GEN_17889; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_18292 = 3'h0 == tail ? 1'h0 : _GEN_17898; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18293 = 3'h1 == tail ? 1'h0 : _GEN_17899; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18294 = 3'h2 == tail ? 1'h0 : _GEN_17900; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18295 = 3'h3 == tail ? 1'h0 : _GEN_17901; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18296 = 3'h4 == tail ? 1'h0 : _GEN_17902; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18297 = 3'h5 == tail ? 1'h0 : _GEN_17903; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18298 = 3'h6 == tail ? 1'h0 : _GEN_17904; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18299 = 3'h7 == tail ? 1'h0 : _GEN_17905; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18300 = 3'h0 == tail ? 1'h0 : _GEN_17906; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18301 = 3'h1 == tail ? 1'h0 : _GEN_17907; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18302 = 3'h2 == tail ? 1'h0 : _GEN_17908; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18303 = 3'h3 == tail ? 1'h0 : _GEN_17909; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18304 = 3'h4 == tail ? 1'h0 : _GEN_17910; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18305 = 3'h5 == tail ? 1'h0 : _GEN_17911; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18306 = 3'h6 == tail ? 1'h0 : _GEN_17912; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18307 = 3'h7 == tail ? 1'h0 : _GEN_17913; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18308 = 3'h0 == tail ? 1'h0 : _GEN_17914; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18309 = 3'h1 == tail ? 1'h0 : _GEN_17915; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18310 = 3'h2 == tail ? 1'h0 : _GEN_17916; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18311 = 3'h3 == tail ? 1'h0 : _GEN_17917; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18312 = 3'h4 == tail ? 1'h0 : _GEN_17918; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18313 = 3'h5 == tail ? 1'h0 : _GEN_17919; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18314 = 3'h6 == tail ? 1'h0 : _GEN_17920; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18315 = 3'h7 == tail ? 1'h0 : _GEN_17921; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18316 = 3'h0 == tail ? 1'h0 : _GEN_17922; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18317 = 3'h1 == tail ? 1'h0 : _GEN_17923; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18318 = 3'h2 == tail ? 1'h0 : _GEN_17924; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18319 = 3'h3 == tail ? 1'h0 : _GEN_17925; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18320 = 3'h4 == tail ? 1'h0 : _GEN_17926; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18321 = 3'h5 == tail ? 1'h0 : _GEN_17927; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18322 = 3'h6 == tail ? 1'h0 : _GEN_17928; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18323 = 3'h7 == tail ? 1'h0 : _GEN_17929; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18324 = 3'h0 == tail ? 1'h0 : _GEN_17930; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18325 = 3'h1 == tail ? 1'h0 : _GEN_17931; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18326 = 3'h2 == tail ? 1'h0 : _GEN_17932; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18327 = 3'h3 == tail ? 1'h0 : _GEN_17933; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18328 = 3'h4 == tail ? 1'h0 : _GEN_17934; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18329 = 3'h5 == tail ? 1'h0 : _GEN_17935; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18330 = 3'h6 == tail ? 1'h0 : _GEN_17936; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18331 = 3'h7 == tail ? 1'h0 : _GEN_17937; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18332 = 3'h0 == tail ? 1'h0 : _GEN_17938; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18333 = 3'h1 == tail ? 1'h0 : _GEN_17939; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18334 = 3'h2 == tail ? 1'h0 : _GEN_17940; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18335 = 3'h3 == tail ? 1'h0 : _GEN_17941; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18336 = 3'h4 == tail ? 1'h0 : _GEN_17942; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18337 = 3'h5 == tail ? 1'h0 : _GEN_17943; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18338 = 3'h6 == tail ? 1'h0 : _GEN_17944; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18339 = 3'h7 == tail ? 1'h0 : _GEN_17945; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18340 = 3'h0 == tail ? 1'h0 : _GEN_17946; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18341 = 3'h1 == tail ? 1'h0 : _GEN_17947; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18342 = 3'h2 == tail ? 1'h0 : _GEN_17948; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18343 = 3'h3 == tail ? 1'h0 : _GEN_17949; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18344 = 3'h4 == tail ? 1'h0 : _GEN_17950; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18345 = 3'h5 == tail ? 1'h0 : _GEN_17951; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18346 = 3'h6 == tail ? 1'h0 : _GEN_17952; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18347 = 3'h7 == tail ? 1'h0 : _GEN_17953; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18348 = 3'h0 == tail ? 1'h0 : _GEN_17954; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18349 = 3'h1 == tail ? 1'h0 : _GEN_17955; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18350 = 3'h2 == tail ? 1'h0 : _GEN_17956; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18351 = 3'h3 == tail ? 1'h0 : _GEN_17957; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18352 = 3'h4 == tail ? 1'h0 : _GEN_17958; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18353 = 3'h5 == tail ? 1'h0 : _GEN_17959; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18354 = 3'h6 == tail ? 1'h0 : _GEN_17960; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18355 = 3'h7 == tail ? 1'h0 : _GEN_17961; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18356 = 3'h0 == tail ? 1'h0 : _GEN_17962; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18357 = 3'h1 == tail ? 1'h0 : _GEN_17963; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18358 = 3'h2 == tail ? 1'h0 : _GEN_17964; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18359 = 3'h3 == tail ? 1'h0 : _GEN_17965; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18360 = 3'h4 == tail ? 1'h0 : _GEN_17966; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18361 = 3'h5 == tail ? 1'h0 : _GEN_17967; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18362 = 3'h6 == tail ? 1'h0 : _GEN_17968; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18363 = 3'h7 == tail ? 1'h0 : _GEN_17969; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18364 = 3'h0 == tail ? 1'h0 : _GEN_17970; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18365 = 3'h1 == tail ? 1'h0 : _GEN_17971; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18366 = 3'h2 == tail ? 1'h0 : _GEN_17972; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18367 = 3'h3 == tail ? 1'h0 : _GEN_17973; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18368 = 3'h4 == tail ? 1'h0 : _GEN_17974; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18369 = 3'h5 == tail ? 1'h0 : _GEN_17975; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18370 = 3'h6 == tail ? 1'h0 : _GEN_17976; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18371 = 3'h7 == tail ? 1'h0 : _GEN_17977; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18372 = 3'h0 == tail ? 1'h0 : _GEN_17978; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18373 = 3'h1 == tail ? 1'h0 : _GEN_17979; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18374 = 3'h2 == tail ? 1'h0 : _GEN_17980; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18375 = 3'h3 == tail ? 1'h0 : _GEN_17981; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18376 = 3'h4 == tail ? 1'h0 : _GEN_17982; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18377 = 3'h5 == tail ? 1'h0 : _GEN_17983; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18378 = 3'h6 == tail ? 1'h0 : _GEN_17984; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18379 = 3'h7 == tail ? 1'h0 : _GEN_17985; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18380 = 3'h0 == tail ? 1'h0 : _GEN_17986; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18381 = 3'h1 == tail ? 1'h0 : _GEN_17987; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18382 = 3'h2 == tail ? 1'h0 : _GEN_17988; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18383 = 3'h3 == tail ? 1'h0 : _GEN_17989; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18384 = 3'h4 == tail ? 1'h0 : _GEN_17990; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18385 = 3'h5 == tail ? 1'h0 : _GEN_17991; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18386 = 3'h6 == tail ? 1'h0 : _GEN_17992; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18387 = 3'h7 == tail ? 1'h0 : _GEN_17993; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18388 = 3'h0 == tail ? 1'h0 : _GEN_17994; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18389 = 3'h1 == tail ? 1'h0 : _GEN_17995; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18390 = 3'h2 == tail ? 1'h0 : _GEN_17996; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18391 = 3'h3 == tail ? 1'h0 : _GEN_17997; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18392 = 3'h4 == tail ? 1'h0 : _GEN_17998; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18393 = 3'h5 == tail ? 1'h0 : _GEN_17999; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18394 = 3'h6 == tail ? 1'h0 : _GEN_18000; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18395 = 3'h7 == tail ? 1'h0 : _GEN_18001; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18396 = 3'h0 == tail ? 1'h0 : _GEN_18002; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18397 = 3'h1 == tail ? 1'h0 : _GEN_18003; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18398 = 3'h2 == tail ? 1'h0 : _GEN_18004; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18399 = 3'h3 == tail ? 1'h0 : _GEN_18005; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18400 = 3'h4 == tail ? 1'h0 : _GEN_18006; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18401 = 3'h5 == tail ? 1'h0 : _GEN_18007; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18402 = 3'h6 == tail ? 1'h0 : _GEN_18008; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18403 = 3'h7 == tail ? 1'h0 : _GEN_18009; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18404 = 3'h0 == tail ? 1'h0 : _GEN_18010; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18405 = 3'h1 == tail ? 1'h0 : _GEN_18011; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18406 = 3'h2 == tail ? 1'h0 : _GEN_18012; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18407 = 3'h3 == tail ? 1'h0 : _GEN_18013; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18408 = 3'h4 == tail ? 1'h0 : _GEN_18014; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18409 = 3'h5 == tail ? 1'h0 : _GEN_18015; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18410 = 3'h6 == tail ? 1'h0 : _GEN_18016; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18411 = 3'h7 == tail ? 1'h0 : _GEN_18017; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18412 = 3'h0 == tail ? 1'h0 : _GEN_18018; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18413 = 3'h1 == tail ? 1'h0 : _GEN_18019; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18414 = 3'h2 == tail ? 1'h0 : _GEN_18020; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18415 = 3'h3 == tail ? 1'h0 : _GEN_18021; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18416 = 3'h4 == tail ? 1'h0 : _GEN_18022; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18417 = 3'h5 == tail ? 1'h0 : _GEN_18023; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18418 = 3'h6 == tail ? 1'h0 : _GEN_18024; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18419 = 3'h7 == tail ? 1'h0 : _GEN_18025; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18420 = 3'h0 == tail ? 1'h0 : _GEN_18026; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18421 = 3'h1 == tail ? 1'h0 : _GEN_18027; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18422 = 3'h2 == tail ? 1'h0 : _GEN_18028; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18423 = 3'h3 == tail ? 1'h0 : _GEN_18029; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18424 = 3'h4 == tail ? 1'h0 : _GEN_18030; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18425 = 3'h5 == tail ? 1'h0 : _GEN_18031; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18426 = 3'h6 == tail ? 1'h0 : _GEN_18032; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18427 = 3'h7 == tail ? 1'h0 : _GEN_18033; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18428 = 3'h0 == tail ? 1'h0 : _GEN_18034; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18429 = 3'h1 == tail ? 1'h0 : _GEN_18035; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18430 = 3'h2 == tail ? 1'h0 : _GEN_18036; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18431 = 3'h3 == tail ? 1'h0 : _GEN_18037; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18432 = 3'h4 == tail ? 1'h0 : _GEN_18038; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18433 = 3'h5 == tail ? 1'h0 : _GEN_18039; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18434 = 3'h6 == tail ? 1'h0 : _GEN_18040; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18435 = 3'h7 == tail ? 1'h0 : _GEN_18041; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18436 = 3'h0 == tail ? 1'h0 : _GEN_18042; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18437 = 3'h1 == tail ? 1'h0 : _GEN_18043; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18438 = 3'h2 == tail ? 1'h0 : _GEN_18044; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18439 = 3'h3 == tail ? 1'h0 : _GEN_18045; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18440 = 3'h4 == tail ? 1'h0 : _GEN_18046; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18441 = 3'h5 == tail ? 1'h0 : _GEN_18047; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18442 = 3'h6 == tail ? 1'h0 : _GEN_18048; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18443 = 3'h7 == tail ? 1'h0 : _GEN_18049; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18444 = 3'h0 == tail ? 1'h0 : _GEN_18050; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18445 = 3'h1 == tail ? 1'h0 : _GEN_18051; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18446 = 3'h2 == tail ? 1'h0 : _GEN_18052; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18447 = 3'h3 == tail ? 1'h0 : _GEN_18053; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18448 = 3'h4 == tail ? 1'h0 : _GEN_18054; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18449 = 3'h5 == tail ? 1'h0 : _GEN_18055; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18450 = 3'h6 == tail ? 1'h0 : _GEN_18056; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18451 = 3'h7 == tail ? 1'h0 : _GEN_18057; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18452 = 3'h0 == tail ? 1'h0 : _GEN_18058; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18453 = 3'h1 == tail ? 1'h0 : _GEN_18059; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18454 = 3'h2 == tail ? 1'h0 : _GEN_18060; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18455 = 3'h3 == tail ? 1'h0 : _GEN_18061; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18456 = 3'h4 == tail ? 1'h0 : _GEN_18062; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18457 = 3'h5 == tail ? 1'h0 : _GEN_18063; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18458 = 3'h6 == tail ? 1'h0 : _GEN_18064; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18459 = 3'h7 == tail ? 1'h0 : _GEN_18065; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18460 = 3'h0 == tail ? 1'h0 : _GEN_18066; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18461 = 3'h1 == tail ? 1'h0 : _GEN_18067; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18462 = 3'h2 == tail ? 1'h0 : _GEN_18068; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18463 = 3'h3 == tail ? 1'h0 : _GEN_18069; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18464 = 3'h4 == tail ? 1'h0 : _GEN_18070; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18465 = 3'h5 == tail ? 1'h0 : _GEN_18071; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18466 = 3'h6 == tail ? 1'h0 : _GEN_18072; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18467 = 3'h7 == tail ? 1'h0 : _GEN_18073; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_18468 = 3'h0 == tail ? 1'h0 : _GEN_18074; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18469 = 3'h1 == tail ? 1'h0 : _GEN_18075; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18470 = 3'h2 == tail ? 1'h0 : _GEN_18076; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18471 = 3'h3 == tail ? 1'h0 : _GEN_18077; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18472 = 3'h4 == tail ? 1'h0 : _GEN_18078; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18473 = 3'h5 == tail ? 1'h0 : _GEN_18079; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18474 = 3'h6 == tail ? 1'h0 : _GEN_18080; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18475 = 3'h7 == tail ? 1'h0 : _GEN_18081; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_18476 = 3'h0 == tail ? 1'h0 : _GEN_18082; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18477 = 3'h1 == tail ? 1'h0 : _GEN_18083; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18478 = 3'h2 == tail ? 1'h0 : _GEN_18084; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18479 = 3'h3 == tail ? 1'h0 : _GEN_18085; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18480 = 3'h4 == tail ? 1'h0 : _GEN_18086; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18481 = 3'h5 == tail ? 1'h0 : _GEN_18087; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18482 = 3'h6 == tail ? 1'h0 : _GEN_18088; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18483 = 3'h7 == tail ? 1'h0 : _GEN_18089; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_18484 = 3'h0 == tail ? 1'h0 : _GEN_18090; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18485 = 3'h1 == tail ? 1'h0 : _GEN_18091; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18486 = 3'h2 == tail ? 1'h0 : _GEN_18092; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18487 = 3'h3 == tail ? 1'h0 : _GEN_18093; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18488 = 3'h4 == tail ? 1'h0 : _GEN_18094; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18489 = 3'h5 == tail ? 1'h0 : _GEN_18095; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18490 = 3'h6 == tail ? 1'h0 : _GEN_18096; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18491 = 3'h7 == tail ? 1'h0 : _GEN_18097; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_18500 = _GEN_32729 | e_0_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18501 = _GEN_32730 | e_1_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18502 = _GEN_32731 | e_2_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18503 = _GEN_32732 | e_3_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18504 = _GEN_32733 | e_4_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18505 = _GEN_32734 | e_5_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18506 = _GEN_32735 | e_6_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_18507 = _GEN_32736 | e_7_active_vgu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_18508 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_18114; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18509 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_18115; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18510 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_18116; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18511 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_18117; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18512 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_18118; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18513 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_18119; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18514 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_18120; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_18515 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_18121; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_18516 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_18122; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18517 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_18123; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18518 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_18124; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18519 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_18125; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18520 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_18126; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18521 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_18127; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18522 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_18128; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_18523 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_18129; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18524 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_18244; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18525 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_18245; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18526 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_18246; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18527 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_18247; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18528 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_18248; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18529 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_18249; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18530 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_18250; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18531 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_18251; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18532 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_18130; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18533 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_18131; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18534 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_18132; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18535 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_18133; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18536 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_18134; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18537 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_18135; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18538 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_18136; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18539 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_18137; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18540 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_18138; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18541 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_18139; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18542 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_18140; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18543 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_18141; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18544 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_18142; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18545 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_18143; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18546 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_18144; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_18547 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_18145; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_18548 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_18146; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18549 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_18147; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18550 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_18148; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18551 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_18149; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18552 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_18150; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18553 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_18151; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18554 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_18152; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_18555 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_18153; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_18556 = io_op_bits_base_vp_valid ? _GEN_18516 : _GEN_18122; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18557 = io_op_bits_base_vp_valid ? _GEN_18517 : _GEN_18123; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18558 = io_op_bits_base_vp_valid ? _GEN_18518 : _GEN_18124; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18559 = io_op_bits_base_vp_valid ? _GEN_18519 : _GEN_18125; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18560 = io_op_bits_base_vp_valid ? _GEN_18520 : _GEN_18126; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18561 = io_op_bits_base_vp_valid ? _GEN_18521 : _GEN_18127; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18562 = io_op_bits_base_vp_valid ? _GEN_18522 : _GEN_18128; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_18563 = io_op_bits_base_vp_valid ? _GEN_18523 : _GEN_18129; // @[sequencer-master.scala 320:41]
  wire  _GEN_18564 = io_op_bits_base_vp_valid ? _GEN_18524 : _GEN_18244; // @[sequencer-master.scala 320:41]
  wire  _GEN_18565 = io_op_bits_base_vp_valid ? _GEN_18525 : _GEN_18245; // @[sequencer-master.scala 320:41]
  wire  _GEN_18566 = io_op_bits_base_vp_valid ? _GEN_18526 : _GEN_18246; // @[sequencer-master.scala 320:41]
  wire  _GEN_18567 = io_op_bits_base_vp_valid ? _GEN_18527 : _GEN_18247; // @[sequencer-master.scala 320:41]
  wire  _GEN_18568 = io_op_bits_base_vp_valid ? _GEN_18528 : _GEN_18248; // @[sequencer-master.scala 320:41]
  wire  _GEN_18569 = io_op_bits_base_vp_valid ? _GEN_18529 : _GEN_18249; // @[sequencer-master.scala 320:41]
  wire  _GEN_18570 = io_op_bits_base_vp_valid ? _GEN_18530 : _GEN_18250; // @[sequencer-master.scala 320:41]
  wire  _GEN_18571 = io_op_bits_base_vp_valid ? _GEN_18531 : _GEN_18251; // @[sequencer-master.scala 320:41]
  wire  _GEN_18572 = io_op_bits_base_vp_valid ? _GEN_18532 : _GEN_18130; // @[sequencer-master.scala 320:41]
  wire  _GEN_18573 = io_op_bits_base_vp_valid ? _GEN_18533 : _GEN_18131; // @[sequencer-master.scala 320:41]
  wire  _GEN_18574 = io_op_bits_base_vp_valid ? _GEN_18534 : _GEN_18132; // @[sequencer-master.scala 320:41]
  wire  _GEN_18575 = io_op_bits_base_vp_valid ? _GEN_18535 : _GEN_18133; // @[sequencer-master.scala 320:41]
  wire  _GEN_18576 = io_op_bits_base_vp_valid ? _GEN_18536 : _GEN_18134; // @[sequencer-master.scala 320:41]
  wire  _GEN_18577 = io_op_bits_base_vp_valid ? _GEN_18537 : _GEN_18135; // @[sequencer-master.scala 320:41]
  wire  _GEN_18578 = io_op_bits_base_vp_valid ? _GEN_18538 : _GEN_18136; // @[sequencer-master.scala 320:41]
  wire  _GEN_18579 = io_op_bits_base_vp_valid ? _GEN_18539 : _GEN_18137; // @[sequencer-master.scala 320:41]
  wire  _GEN_18580 = io_op_bits_base_vp_valid ? _GEN_18540 : _GEN_18138; // @[sequencer-master.scala 320:41]
  wire  _GEN_18581 = io_op_bits_base_vp_valid ? _GEN_18541 : _GEN_18139; // @[sequencer-master.scala 320:41]
  wire  _GEN_18582 = io_op_bits_base_vp_valid ? _GEN_18542 : _GEN_18140; // @[sequencer-master.scala 320:41]
  wire  _GEN_18583 = io_op_bits_base_vp_valid ? _GEN_18543 : _GEN_18141; // @[sequencer-master.scala 320:41]
  wire  _GEN_18584 = io_op_bits_base_vp_valid ? _GEN_18544 : _GEN_18142; // @[sequencer-master.scala 320:41]
  wire  _GEN_18585 = io_op_bits_base_vp_valid ? _GEN_18545 : _GEN_18143; // @[sequencer-master.scala 320:41]
  wire  _GEN_18586 = io_op_bits_base_vp_valid ? _GEN_18546 : _GEN_18144; // @[sequencer-master.scala 320:41]
  wire  _GEN_18587 = io_op_bits_base_vp_valid ? _GEN_18547 : _GEN_18145; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18588 = io_op_bits_base_vp_valid ? _GEN_18548 : _GEN_18146; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18589 = io_op_bits_base_vp_valid ? _GEN_18549 : _GEN_18147; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18590 = io_op_bits_base_vp_valid ? _GEN_18550 : _GEN_18148; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18591 = io_op_bits_base_vp_valid ? _GEN_18551 : _GEN_18149; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18592 = io_op_bits_base_vp_valid ? _GEN_18552 : _GEN_18150; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18593 = io_op_bits_base_vp_valid ? _GEN_18553 : _GEN_18151; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18594 = io_op_bits_base_vp_valid ? _GEN_18554 : _GEN_18152; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_18595 = io_op_bits_base_vp_valid ? _GEN_18555 : _GEN_18153; // @[sequencer-master.scala 320:41]
  wire  _GEN_18596 = _GEN_32729 | _GEN_18292; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18597 = _GEN_32730 | _GEN_18293; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18598 = _GEN_32731 | _GEN_18294; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18599 = _GEN_32732 | _GEN_18295; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18600 = _GEN_32733 | _GEN_18296; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18601 = _GEN_32734 | _GEN_18297; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18602 = _GEN_32735 | _GEN_18298; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18603 = _GEN_32736 | _GEN_18299; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18604 = _T_26 ? _GEN_18596 : _GEN_18292; // @[sequencer-master.scala 154:24]
  wire  _GEN_18605 = _T_26 ? _GEN_18597 : _GEN_18293; // @[sequencer-master.scala 154:24]
  wire  _GEN_18606 = _T_26 ? _GEN_18598 : _GEN_18294; // @[sequencer-master.scala 154:24]
  wire  _GEN_18607 = _T_26 ? _GEN_18599 : _GEN_18295; // @[sequencer-master.scala 154:24]
  wire  _GEN_18608 = _T_26 ? _GEN_18600 : _GEN_18296; // @[sequencer-master.scala 154:24]
  wire  _GEN_18609 = _T_26 ? _GEN_18601 : _GEN_18297; // @[sequencer-master.scala 154:24]
  wire  _GEN_18610 = _T_26 ? _GEN_18602 : _GEN_18298; // @[sequencer-master.scala 154:24]
  wire  _GEN_18611 = _T_26 ? _GEN_18603 : _GEN_18299; // @[sequencer-master.scala 154:24]
  wire  _GEN_18612 = _GEN_32729 | _GEN_18316; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18613 = _GEN_32730 | _GEN_18317; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18614 = _GEN_32731 | _GEN_18318; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18615 = _GEN_32732 | _GEN_18319; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18616 = _GEN_32733 | _GEN_18320; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18617 = _GEN_32734 | _GEN_18321; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18618 = _GEN_32735 | _GEN_18322; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18619 = _GEN_32736 | _GEN_18323; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18620 = _T_48 ? _GEN_18612 : _GEN_18316; // @[sequencer-master.scala 154:24]
  wire  _GEN_18621 = _T_48 ? _GEN_18613 : _GEN_18317; // @[sequencer-master.scala 154:24]
  wire  _GEN_18622 = _T_48 ? _GEN_18614 : _GEN_18318; // @[sequencer-master.scala 154:24]
  wire  _GEN_18623 = _T_48 ? _GEN_18615 : _GEN_18319; // @[sequencer-master.scala 154:24]
  wire  _GEN_18624 = _T_48 ? _GEN_18616 : _GEN_18320; // @[sequencer-master.scala 154:24]
  wire  _GEN_18625 = _T_48 ? _GEN_18617 : _GEN_18321; // @[sequencer-master.scala 154:24]
  wire  _GEN_18626 = _T_48 ? _GEN_18618 : _GEN_18322; // @[sequencer-master.scala 154:24]
  wire  _GEN_18627 = _T_48 ? _GEN_18619 : _GEN_18323; // @[sequencer-master.scala 154:24]
  wire  _GEN_18628 = _GEN_32729 | _GEN_18340; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18629 = _GEN_32730 | _GEN_18341; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18630 = _GEN_32731 | _GEN_18342; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18631 = _GEN_32732 | _GEN_18343; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18632 = _GEN_32733 | _GEN_18344; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18633 = _GEN_32734 | _GEN_18345; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18634 = _GEN_32735 | _GEN_18346; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18635 = _GEN_32736 | _GEN_18347; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18636 = _T_70 ? _GEN_18628 : _GEN_18340; // @[sequencer-master.scala 154:24]
  wire  _GEN_18637 = _T_70 ? _GEN_18629 : _GEN_18341; // @[sequencer-master.scala 154:24]
  wire  _GEN_18638 = _T_70 ? _GEN_18630 : _GEN_18342; // @[sequencer-master.scala 154:24]
  wire  _GEN_18639 = _T_70 ? _GEN_18631 : _GEN_18343; // @[sequencer-master.scala 154:24]
  wire  _GEN_18640 = _T_70 ? _GEN_18632 : _GEN_18344; // @[sequencer-master.scala 154:24]
  wire  _GEN_18641 = _T_70 ? _GEN_18633 : _GEN_18345; // @[sequencer-master.scala 154:24]
  wire  _GEN_18642 = _T_70 ? _GEN_18634 : _GEN_18346; // @[sequencer-master.scala 154:24]
  wire  _GEN_18643 = _T_70 ? _GEN_18635 : _GEN_18347; // @[sequencer-master.scala 154:24]
  wire  _GEN_18644 = _GEN_32729 | _GEN_18364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18645 = _GEN_32730 | _GEN_18365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18646 = _GEN_32731 | _GEN_18366; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18647 = _GEN_32732 | _GEN_18367; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18648 = _GEN_32733 | _GEN_18368; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18649 = _GEN_32734 | _GEN_18369; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18650 = _GEN_32735 | _GEN_18370; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18651 = _GEN_32736 | _GEN_18371; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18652 = _T_92 ? _GEN_18644 : _GEN_18364; // @[sequencer-master.scala 154:24]
  wire  _GEN_18653 = _T_92 ? _GEN_18645 : _GEN_18365; // @[sequencer-master.scala 154:24]
  wire  _GEN_18654 = _T_92 ? _GEN_18646 : _GEN_18366; // @[sequencer-master.scala 154:24]
  wire  _GEN_18655 = _T_92 ? _GEN_18647 : _GEN_18367; // @[sequencer-master.scala 154:24]
  wire  _GEN_18656 = _T_92 ? _GEN_18648 : _GEN_18368; // @[sequencer-master.scala 154:24]
  wire  _GEN_18657 = _T_92 ? _GEN_18649 : _GEN_18369; // @[sequencer-master.scala 154:24]
  wire  _GEN_18658 = _T_92 ? _GEN_18650 : _GEN_18370; // @[sequencer-master.scala 154:24]
  wire  _GEN_18659 = _T_92 ? _GEN_18651 : _GEN_18371; // @[sequencer-master.scala 154:24]
  wire  _GEN_18660 = _GEN_32729 | _GEN_18388; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18661 = _GEN_32730 | _GEN_18389; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18662 = _GEN_32731 | _GEN_18390; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18663 = _GEN_32732 | _GEN_18391; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18664 = _GEN_32733 | _GEN_18392; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18665 = _GEN_32734 | _GEN_18393; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18666 = _GEN_32735 | _GEN_18394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18667 = _GEN_32736 | _GEN_18395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18668 = _T_114 ? _GEN_18660 : _GEN_18388; // @[sequencer-master.scala 154:24]
  wire  _GEN_18669 = _T_114 ? _GEN_18661 : _GEN_18389; // @[sequencer-master.scala 154:24]
  wire  _GEN_18670 = _T_114 ? _GEN_18662 : _GEN_18390; // @[sequencer-master.scala 154:24]
  wire  _GEN_18671 = _T_114 ? _GEN_18663 : _GEN_18391; // @[sequencer-master.scala 154:24]
  wire  _GEN_18672 = _T_114 ? _GEN_18664 : _GEN_18392; // @[sequencer-master.scala 154:24]
  wire  _GEN_18673 = _T_114 ? _GEN_18665 : _GEN_18393; // @[sequencer-master.scala 154:24]
  wire  _GEN_18674 = _T_114 ? _GEN_18666 : _GEN_18394; // @[sequencer-master.scala 154:24]
  wire  _GEN_18675 = _T_114 ? _GEN_18667 : _GEN_18395; // @[sequencer-master.scala 154:24]
  wire  _GEN_18676 = _GEN_32729 | _GEN_18412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18677 = _GEN_32730 | _GEN_18413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18678 = _GEN_32731 | _GEN_18414; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18679 = _GEN_32732 | _GEN_18415; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18680 = _GEN_32733 | _GEN_18416; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18681 = _GEN_32734 | _GEN_18417; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18682 = _GEN_32735 | _GEN_18418; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18683 = _GEN_32736 | _GEN_18419; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18684 = _T_136 ? _GEN_18676 : _GEN_18412; // @[sequencer-master.scala 154:24]
  wire  _GEN_18685 = _T_136 ? _GEN_18677 : _GEN_18413; // @[sequencer-master.scala 154:24]
  wire  _GEN_18686 = _T_136 ? _GEN_18678 : _GEN_18414; // @[sequencer-master.scala 154:24]
  wire  _GEN_18687 = _T_136 ? _GEN_18679 : _GEN_18415; // @[sequencer-master.scala 154:24]
  wire  _GEN_18688 = _T_136 ? _GEN_18680 : _GEN_18416; // @[sequencer-master.scala 154:24]
  wire  _GEN_18689 = _T_136 ? _GEN_18681 : _GEN_18417; // @[sequencer-master.scala 154:24]
  wire  _GEN_18690 = _T_136 ? _GEN_18682 : _GEN_18418; // @[sequencer-master.scala 154:24]
  wire  _GEN_18691 = _T_136 ? _GEN_18683 : _GEN_18419; // @[sequencer-master.scala 154:24]
  wire  _GEN_18692 = _GEN_32729 | _GEN_18436; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18693 = _GEN_32730 | _GEN_18437; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18694 = _GEN_32731 | _GEN_18438; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18695 = _GEN_32732 | _GEN_18439; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18696 = _GEN_32733 | _GEN_18440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18697 = _GEN_32734 | _GEN_18441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18698 = _GEN_32735 | _GEN_18442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18699 = _GEN_32736 | _GEN_18443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18700 = _T_158 ? _GEN_18692 : _GEN_18436; // @[sequencer-master.scala 154:24]
  wire  _GEN_18701 = _T_158 ? _GEN_18693 : _GEN_18437; // @[sequencer-master.scala 154:24]
  wire  _GEN_18702 = _T_158 ? _GEN_18694 : _GEN_18438; // @[sequencer-master.scala 154:24]
  wire  _GEN_18703 = _T_158 ? _GEN_18695 : _GEN_18439; // @[sequencer-master.scala 154:24]
  wire  _GEN_18704 = _T_158 ? _GEN_18696 : _GEN_18440; // @[sequencer-master.scala 154:24]
  wire  _GEN_18705 = _T_158 ? _GEN_18697 : _GEN_18441; // @[sequencer-master.scala 154:24]
  wire  _GEN_18706 = _T_158 ? _GEN_18698 : _GEN_18442; // @[sequencer-master.scala 154:24]
  wire  _GEN_18707 = _T_158 ? _GEN_18699 : _GEN_18443; // @[sequencer-master.scala 154:24]
  wire  _GEN_18708 = _GEN_32729 | _GEN_18460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18709 = _GEN_32730 | _GEN_18461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18710 = _GEN_32731 | _GEN_18462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18711 = _GEN_32732 | _GEN_18463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18712 = _GEN_32733 | _GEN_18464; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18713 = _GEN_32734 | _GEN_18465; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18714 = _GEN_32735 | _GEN_18466; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18715 = _GEN_32736 | _GEN_18467; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18716 = _T_180 ? _GEN_18708 : _GEN_18460; // @[sequencer-master.scala 154:24]
  wire  _GEN_18717 = _T_180 ? _GEN_18709 : _GEN_18461; // @[sequencer-master.scala 154:24]
  wire  _GEN_18718 = _T_180 ? _GEN_18710 : _GEN_18462; // @[sequencer-master.scala 154:24]
  wire  _GEN_18719 = _T_180 ? _GEN_18711 : _GEN_18463; // @[sequencer-master.scala 154:24]
  wire  _GEN_18720 = _T_180 ? _GEN_18712 : _GEN_18464; // @[sequencer-master.scala 154:24]
  wire  _GEN_18721 = _T_180 ? _GEN_18713 : _GEN_18465; // @[sequencer-master.scala 154:24]
  wire  _GEN_18722 = _T_180 ? _GEN_18714 : _GEN_18466; // @[sequencer-master.scala 154:24]
  wire  _GEN_18723 = _T_180 ? _GEN_18715 : _GEN_18467; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_18724 = 3'h0 == tail ? io_op_bits_base_vs1_id : _GEN_18154; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18725 = 3'h1 == tail ? io_op_bits_base_vs1_id : _GEN_18155; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18726 = 3'h2 == tail ? io_op_bits_base_vs1_id : _GEN_18156; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18727 = 3'h3 == tail ? io_op_bits_base_vs1_id : _GEN_18157; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18728 = 3'h4 == tail ? io_op_bits_base_vs1_id : _GEN_18158; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18729 = 3'h5 == tail ? io_op_bits_base_vs1_id : _GEN_18159; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18730 = 3'h6 == tail ? io_op_bits_base_vs1_id : _GEN_18160; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18731 = 3'h7 == tail ? io_op_bits_base_vs1_id : _GEN_18161; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18732 = 3'h0 == tail ? io_op_bits_base_vs1_valid : _GEN_18252; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18733 = 3'h1 == tail ? io_op_bits_base_vs1_valid : _GEN_18253; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18734 = 3'h2 == tail ? io_op_bits_base_vs1_valid : _GEN_18254; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18735 = 3'h3 == tail ? io_op_bits_base_vs1_valid : _GEN_18255; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18736 = 3'h4 == tail ? io_op_bits_base_vs1_valid : _GEN_18256; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18737 = 3'h5 == tail ? io_op_bits_base_vs1_valid : _GEN_18257; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18738 = 3'h6 == tail ? io_op_bits_base_vs1_valid : _GEN_18258; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18739 = 3'h7 == tail ? io_op_bits_base_vs1_valid : _GEN_18259; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18740 = 3'h0 == tail ? io_op_bits_base_vs1_scalar : _GEN_18162; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18741 = 3'h1 == tail ? io_op_bits_base_vs1_scalar : _GEN_18163; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18742 = 3'h2 == tail ? io_op_bits_base_vs1_scalar : _GEN_18164; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18743 = 3'h3 == tail ? io_op_bits_base_vs1_scalar : _GEN_18165; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18744 = 3'h4 == tail ? io_op_bits_base_vs1_scalar : _GEN_18166; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18745 = 3'h5 == tail ? io_op_bits_base_vs1_scalar : _GEN_18167; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18746 = 3'h6 == tail ? io_op_bits_base_vs1_scalar : _GEN_18168; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18747 = 3'h7 == tail ? io_op_bits_base_vs1_scalar : _GEN_18169; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18748 = 3'h0 == tail ? io_op_bits_base_vs1_pred : _GEN_18170; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18749 = 3'h1 == tail ? io_op_bits_base_vs1_pred : _GEN_18171; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18750 = 3'h2 == tail ? io_op_bits_base_vs1_pred : _GEN_18172; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18751 = 3'h3 == tail ? io_op_bits_base_vs1_pred : _GEN_18173; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18752 = 3'h4 == tail ? io_op_bits_base_vs1_pred : _GEN_18174; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18753 = 3'h5 == tail ? io_op_bits_base_vs1_pred : _GEN_18175; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18754 = 3'h6 == tail ? io_op_bits_base_vs1_pred : _GEN_18176; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_18755 = 3'h7 == tail ? io_op_bits_base_vs1_pred : _GEN_18177; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18756 = 3'h0 == tail ? io_op_bits_base_vs1_prec : _GEN_18178; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18757 = 3'h1 == tail ? io_op_bits_base_vs1_prec : _GEN_18179; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18758 = 3'h2 == tail ? io_op_bits_base_vs1_prec : _GEN_18180; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18759 = 3'h3 == tail ? io_op_bits_base_vs1_prec : _GEN_18181; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18760 = 3'h4 == tail ? io_op_bits_base_vs1_prec : _GEN_18182; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18761 = 3'h5 == tail ? io_op_bits_base_vs1_prec : _GEN_18183; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18762 = 3'h6 == tail ? io_op_bits_base_vs1_prec : _GEN_18184; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_18763 = 3'h7 == tail ? io_op_bits_base_vs1_prec : _GEN_18185; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_18764 = 3'h0 == tail ? io_op_bits_reg_vs1_id : _GEN_18186; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18765 = 3'h1 == tail ? io_op_bits_reg_vs1_id : _GEN_18187; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18766 = 3'h2 == tail ? io_op_bits_reg_vs1_id : _GEN_18188; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18767 = 3'h3 == tail ? io_op_bits_reg_vs1_id : _GEN_18189; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18768 = 3'h4 == tail ? io_op_bits_reg_vs1_id : _GEN_18190; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18769 = 3'h5 == tail ? io_op_bits_reg_vs1_id : _GEN_18191; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18770 = 3'h6 == tail ? io_op_bits_reg_vs1_id : _GEN_18192; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_18771 = 3'h7 == tail ? io_op_bits_reg_vs1_id : _GEN_18193; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_18772 = 3'h0 == tail ? io_op_bits_sreg_ss1 : _GEN_18194; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18773 = 3'h1 == tail ? io_op_bits_sreg_ss1 : _GEN_18195; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18774 = 3'h2 == tail ? io_op_bits_sreg_ss1 : _GEN_18196; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18775 = 3'h3 == tail ? io_op_bits_sreg_ss1 : _GEN_18197; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18776 = 3'h4 == tail ? io_op_bits_sreg_ss1 : _GEN_18198; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18777 = 3'h5 == tail ? io_op_bits_sreg_ss1 : _GEN_18199; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18778 = 3'h6 == tail ? io_op_bits_sreg_ss1 : _GEN_18200; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18779 = 3'h7 == tail ? io_op_bits_sreg_ss1 : _GEN_18201; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_18780 = _T_189 ? _GEN_18772 : _GEN_18194; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18781 = _T_189 ? _GEN_18773 : _GEN_18195; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18782 = _T_189 ? _GEN_18774 : _GEN_18196; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18783 = _T_189 ? _GEN_18775 : _GEN_18197; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18784 = _T_189 ? _GEN_18776 : _GEN_18198; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18785 = _T_189 ? _GEN_18777 : _GEN_18199; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18786 = _T_189 ? _GEN_18778 : _GEN_18200; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_18787 = _T_189 ? _GEN_18779 : _GEN_18201; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_18788 = io_op_bits_base_vs1_valid ? _GEN_18724 : _GEN_18154; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18789 = io_op_bits_base_vs1_valid ? _GEN_18725 : _GEN_18155; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18790 = io_op_bits_base_vs1_valid ? _GEN_18726 : _GEN_18156; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18791 = io_op_bits_base_vs1_valid ? _GEN_18727 : _GEN_18157; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18792 = io_op_bits_base_vs1_valid ? _GEN_18728 : _GEN_18158; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18793 = io_op_bits_base_vs1_valid ? _GEN_18729 : _GEN_18159; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18794 = io_op_bits_base_vs1_valid ? _GEN_18730 : _GEN_18160; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18795 = io_op_bits_base_vs1_valid ? _GEN_18731 : _GEN_18161; // @[sequencer-master.scala 328:47]
  wire  _GEN_18796 = io_op_bits_base_vs1_valid ? _GEN_18732 : _GEN_18252; // @[sequencer-master.scala 328:47]
  wire  _GEN_18797 = io_op_bits_base_vs1_valid ? _GEN_18733 : _GEN_18253; // @[sequencer-master.scala 328:47]
  wire  _GEN_18798 = io_op_bits_base_vs1_valid ? _GEN_18734 : _GEN_18254; // @[sequencer-master.scala 328:47]
  wire  _GEN_18799 = io_op_bits_base_vs1_valid ? _GEN_18735 : _GEN_18255; // @[sequencer-master.scala 328:47]
  wire  _GEN_18800 = io_op_bits_base_vs1_valid ? _GEN_18736 : _GEN_18256; // @[sequencer-master.scala 328:47]
  wire  _GEN_18801 = io_op_bits_base_vs1_valid ? _GEN_18737 : _GEN_18257; // @[sequencer-master.scala 328:47]
  wire  _GEN_18802 = io_op_bits_base_vs1_valid ? _GEN_18738 : _GEN_18258; // @[sequencer-master.scala 328:47]
  wire  _GEN_18803 = io_op_bits_base_vs1_valid ? _GEN_18739 : _GEN_18259; // @[sequencer-master.scala 328:47]
  wire  _GEN_18804 = io_op_bits_base_vs1_valid ? _GEN_18740 : _GEN_18162; // @[sequencer-master.scala 328:47]
  wire  _GEN_18805 = io_op_bits_base_vs1_valid ? _GEN_18741 : _GEN_18163; // @[sequencer-master.scala 328:47]
  wire  _GEN_18806 = io_op_bits_base_vs1_valid ? _GEN_18742 : _GEN_18164; // @[sequencer-master.scala 328:47]
  wire  _GEN_18807 = io_op_bits_base_vs1_valid ? _GEN_18743 : _GEN_18165; // @[sequencer-master.scala 328:47]
  wire  _GEN_18808 = io_op_bits_base_vs1_valid ? _GEN_18744 : _GEN_18166; // @[sequencer-master.scala 328:47]
  wire  _GEN_18809 = io_op_bits_base_vs1_valid ? _GEN_18745 : _GEN_18167; // @[sequencer-master.scala 328:47]
  wire  _GEN_18810 = io_op_bits_base_vs1_valid ? _GEN_18746 : _GEN_18168; // @[sequencer-master.scala 328:47]
  wire  _GEN_18811 = io_op_bits_base_vs1_valid ? _GEN_18747 : _GEN_18169; // @[sequencer-master.scala 328:47]
  wire  _GEN_18812 = io_op_bits_base_vs1_valid ? _GEN_18748 : _GEN_18170; // @[sequencer-master.scala 328:47]
  wire  _GEN_18813 = io_op_bits_base_vs1_valid ? _GEN_18749 : _GEN_18171; // @[sequencer-master.scala 328:47]
  wire  _GEN_18814 = io_op_bits_base_vs1_valid ? _GEN_18750 : _GEN_18172; // @[sequencer-master.scala 328:47]
  wire  _GEN_18815 = io_op_bits_base_vs1_valid ? _GEN_18751 : _GEN_18173; // @[sequencer-master.scala 328:47]
  wire  _GEN_18816 = io_op_bits_base_vs1_valid ? _GEN_18752 : _GEN_18174; // @[sequencer-master.scala 328:47]
  wire  _GEN_18817 = io_op_bits_base_vs1_valid ? _GEN_18753 : _GEN_18175; // @[sequencer-master.scala 328:47]
  wire  _GEN_18818 = io_op_bits_base_vs1_valid ? _GEN_18754 : _GEN_18176; // @[sequencer-master.scala 328:47]
  wire  _GEN_18819 = io_op_bits_base_vs1_valid ? _GEN_18755 : _GEN_18177; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18820 = io_op_bits_base_vs1_valid ? _GEN_18756 : _GEN_18178; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18821 = io_op_bits_base_vs1_valid ? _GEN_18757 : _GEN_18179; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18822 = io_op_bits_base_vs1_valid ? _GEN_18758 : _GEN_18180; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18823 = io_op_bits_base_vs1_valid ? _GEN_18759 : _GEN_18181; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18824 = io_op_bits_base_vs1_valid ? _GEN_18760 : _GEN_18182; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18825 = io_op_bits_base_vs1_valid ? _GEN_18761 : _GEN_18183; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18826 = io_op_bits_base_vs1_valid ? _GEN_18762 : _GEN_18184; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_18827 = io_op_bits_base_vs1_valid ? _GEN_18763 : _GEN_18185; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18828 = io_op_bits_base_vs1_valid ? _GEN_18764 : _GEN_18186; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18829 = io_op_bits_base_vs1_valid ? _GEN_18765 : _GEN_18187; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18830 = io_op_bits_base_vs1_valid ? _GEN_18766 : _GEN_18188; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18831 = io_op_bits_base_vs1_valid ? _GEN_18767 : _GEN_18189; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18832 = io_op_bits_base_vs1_valid ? _GEN_18768 : _GEN_18190; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18833 = io_op_bits_base_vs1_valid ? _GEN_18769 : _GEN_18191; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18834 = io_op_bits_base_vs1_valid ? _GEN_18770 : _GEN_18192; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_18835 = io_op_bits_base_vs1_valid ? _GEN_18771 : _GEN_18193; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18836 = io_op_bits_base_vs1_valid ? _GEN_18780 : _GEN_18194; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18837 = io_op_bits_base_vs1_valid ? _GEN_18781 : _GEN_18195; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18838 = io_op_bits_base_vs1_valid ? _GEN_18782 : _GEN_18196; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18839 = io_op_bits_base_vs1_valid ? _GEN_18783 : _GEN_18197; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18840 = io_op_bits_base_vs1_valid ? _GEN_18784 : _GEN_18198; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18841 = io_op_bits_base_vs1_valid ? _GEN_18785 : _GEN_18199; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18842 = io_op_bits_base_vs1_valid ? _GEN_18786 : _GEN_18200; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_18843 = io_op_bits_base_vs1_valid ? _GEN_18787 : _GEN_18201; // @[sequencer-master.scala 328:47]
  wire  _GEN_18844 = _GEN_32729 | _GEN_18604; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18845 = _GEN_32730 | _GEN_18605; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18846 = _GEN_32731 | _GEN_18606; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18847 = _GEN_32732 | _GEN_18607; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18848 = _GEN_32733 | _GEN_18608; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18849 = _GEN_32734 | _GEN_18609; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18850 = _GEN_32735 | _GEN_18610; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18851 = _GEN_32736 | _GEN_18611; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18852 = _T_203 ? _GEN_18844 : _GEN_18604; // @[sequencer-master.scala 154:24]
  wire  _GEN_18853 = _T_203 ? _GEN_18845 : _GEN_18605; // @[sequencer-master.scala 154:24]
  wire  _GEN_18854 = _T_203 ? _GEN_18846 : _GEN_18606; // @[sequencer-master.scala 154:24]
  wire  _GEN_18855 = _T_203 ? _GEN_18847 : _GEN_18607; // @[sequencer-master.scala 154:24]
  wire  _GEN_18856 = _T_203 ? _GEN_18848 : _GEN_18608; // @[sequencer-master.scala 154:24]
  wire  _GEN_18857 = _T_203 ? _GEN_18849 : _GEN_18609; // @[sequencer-master.scala 154:24]
  wire  _GEN_18858 = _T_203 ? _GEN_18850 : _GEN_18610; // @[sequencer-master.scala 154:24]
  wire  _GEN_18859 = _T_203 ? _GEN_18851 : _GEN_18611; // @[sequencer-master.scala 154:24]
  wire  _GEN_18860 = _GEN_32729 | _GEN_18620; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18861 = _GEN_32730 | _GEN_18621; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18862 = _GEN_32731 | _GEN_18622; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18863 = _GEN_32732 | _GEN_18623; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18864 = _GEN_32733 | _GEN_18624; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18865 = _GEN_32734 | _GEN_18625; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18866 = _GEN_32735 | _GEN_18626; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18867 = _GEN_32736 | _GEN_18627; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18868 = _T_225 ? _GEN_18860 : _GEN_18620; // @[sequencer-master.scala 154:24]
  wire  _GEN_18869 = _T_225 ? _GEN_18861 : _GEN_18621; // @[sequencer-master.scala 154:24]
  wire  _GEN_18870 = _T_225 ? _GEN_18862 : _GEN_18622; // @[sequencer-master.scala 154:24]
  wire  _GEN_18871 = _T_225 ? _GEN_18863 : _GEN_18623; // @[sequencer-master.scala 154:24]
  wire  _GEN_18872 = _T_225 ? _GEN_18864 : _GEN_18624; // @[sequencer-master.scala 154:24]
  wire  _GEN_18873 = _T_225 ? _GEN_18865 : _GEN_18625; // @[sequencer-master.scala 154:24]
  wire  _GEN_18874 = _T_225 ? _GEN_18866 : _GEN_18626; // @[sequencer-master.scala 154:24]
  wire  _GEN_18875 = _T_225 ? _GEN_18867 : _GEN_18627; // @[sequencer-master.scala 154:24]
  wire  _GEN_18876 = _GEN_32729 | _GEN_18636; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18877 = _GEN_32730 | _GEN_18637; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18878 = _GEN_32731 | _GEN_18638; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18879 = _GEN_32732 | _GEN_18639; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18880 = _GEN_32733 | _GEN_18640; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18881 = _GEN_32734 | _GEN_18641; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18882 = _GEN_32735 | _GEN_18642; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18883 = _GEN_32736 | _GEN_18643; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18884 = _T_247 ? _GEN_18876 : _GEN_18636; // @[sequencer-master.scala 154:24]
  wire  _GEN_18885 = _T_247 ? _GEN_18877 : _GEN_18637; // @[sequencer-master.scala 154:24]
  wire  _GEN_18886 = _T_247 ? _GEN_18878 : _GEN_18638; // @[sequencer-master.scala 154:24]
  wire  _GEN_18887 = _T_247 ? _GEN_18879 : _GEN_18639; // @[sequencer-master.scala 154:24]
  wire  _GEN_18888 = _T_247 ? _GEN_18880 : _GEN_18640; // @[sequencer-master.scala 154:24]
  wire  _GEN_18889 = _T_247 ? _GEN_18881 : _GEN_18641; // @[sequencer-master.scala 154:24]
  wire  _GEN_18890 = _T_247 ? _GEN_18882 : _GEN_18642; // @[sequencer-master.scala 154:24]
  wire  _GEN_18891 = _T_247 ? _GEN_18883 : _GEN_18643; // @[sequencer-master.scala 154:24]
  wire  _GEN_18892 = _GEN_32729 | _GEN_18652; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18893 = _GEN_32730 | _GEN_18653; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18894 = _GEN_32731 | _GEN_18654; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18895 = _GEN_32732 | _GEN_18655; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18896 = _GEN_32733 | _GEN_18656; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18897 = _GEN_32734 | _GEN_18657; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18898 = _GEN_32735 | _GEN_18658; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18899 = _GEN_32736 | _GEN_18659; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18900 = _T_269 ? _GEN_18892 : _GEN_18652; // @[sequencer-master.scala 154:24]
  wire  _GEN_18901 = _T_269 ? _GEN_18893 : _GEN_18653; // @[sequencer-master.scala 154:24]
  wire  _GEN_18902 = _T_269 ? _GEN_18894 : _GEN_18654; // @[sequencer-master.scala 154:24]
  wire  _GEN_18903 = _T_269 ? _GEN_18895 : _GEN_18655; // @[sequencer-master.scala 154:24]
  wire  _GEN_18904 = _T_269 ? _GEN_18896 : _GEN_18656; // @[sequencer-master.scala 154:24]
  wire  _GEN_18905 = _T_269 ? _GEN_18897 : _GEN_18657; // @[sequencer-master.scala 154:24]
  wire  _GEN_18906 = _T_269 ? _GEN_18898 : _GEN_18658; // @[sequencer-master.scala 154:24]
  wire  _GEN_18907 = _T_269 ? _GEN_18899 : _GEN_18659; // @[sequencer-master.scala 154:24]
  wire  _GEN_18908 = _GEN_32729 | _GEN_18668; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18909 = _GEN_32730 | _GEN_18669; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18910 = _GEN_32731 | _GEN_18670; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18911 = _GEN_32732 | _GEN_18671; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18912 = _GEN_32733 | _GEN_18672; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18913 = _GEN_32734 | _GEN_18673; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18914 = _GEN_32735 | _GEN_18674; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18915 = _GEN_32736 | _GEN_18675; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18916 = _T_291 ? _GEN_18908 : _GEN_18668; // @[sequencer-master.scala 154:24]
  wire  _GEN_18917 = _T_291 ? _GEN_18909 : _GEN_18669; // @[sequencer-master.scala 154:24]
  wire  _GEN_18918 = _T_291 ? _GEN_18910 : _GEN_18670; // @[sequencer-master.scala 154:24]
  wire  _GEN_18919 = _T_291 ? _GEN_18911 : _GEN_18671; // @[sequencer-master.scala 154:24]
  wire  _GEN_18920 = _T_291 ? _GEN_18912 : _GEN_18672; // @[sequencer-master.scala 154:24]
  wire  _GEN_18921 = _T_291 ? _GEN_18913 : _GEN_18673; // @[sequencer-master.scala 154:24]
  wire  _GEN_18922 = _T_291 ? _GEN_18914 : _GEN_18674; // @[sequencer-master.scala 154:24]
  wire  _GEN_18923 = _T_291 ? _GEN_18915 : _GEN_18675; // @[sequencer-master.scala 154:24]
  wire  _GEN_18924 = _GEN_32729 | _GEN_18684; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18925 = _GEN_32730 | _GEN_18685; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18926 = _GEN_32731 | _GEN_18686; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18927 = _GEN_32732 | _GEN_18687; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18928 = _GEN_32733 | _GEN_18688; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18929 = _GEN_32734 | _GEN_18689; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18930 = _GEN_32735 | _GEN_18690; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18931 = _GEN_32736 | _GEN_18691; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18932 = _T_313 ? _GEN_18924 : _GEN_18684; // @[sequencer-master.scala 154:24]
  wire  _GEN_18933 = _T_313 ? _GEN_18925 : _GEN_18685; // @[sequencer-master.scala 154:24]
  wire  _GEN_18934 = _T_313 ? _GEN_18926 : _GEN_18686; // @[sequencer-master.scala 154:24]
  wire  _GEN_18935 = _T_313 ? _GEN_18927 : _GEN_18687; // @[sequencer-master.scala 154:24]
  wire  _GEN_18936 = _T_313 ? _GEN_18928 : _GEN_18688; // @[sequencer-master.scala 154:24]
  wire  _GEN_18937 = _T_313 ? _GEN_18929 : _GEN_18689; // @[sequencer-master.scala 154:24]
  wire  _GEN_18938 = _T_313 ? _GEN_18930 : _GEN_18690; // @[sequencer-master.scala 154:24]
  wire  _GEN_18939 = _T_313 ? _GEN_18931 : _GEN_18691; // @[sequencer-master.scala 154:24]
  wire  _GEN_18940 = _GEN_32729 | _GEN_18700; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18941 = _GEN_32730 | _GEN_18701; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18942 = _GEN_32731 | _GEN_18702; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18943 = _GEN_32732 | _GEN_18703; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18944 = _GEN_32733 | _GEN_18704; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18945 = _GEN_32734 | _GEN_18705; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18946 = _GEN_32735 | _GEN_18706; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18947 = _GEN_32736 | _GEN_18707; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18948 = _T_335 ? _GEN_18940 : _GEN_18700; // @[sequencer-master.scala 154:24]
  wire  _GEN_18949 = _T_335 ? _GEN_18941 : _GEN_18701; // @[sequencer-master.scala 154:24]
  wire  _GEN_18950 = _T_335 ? _GEN_18942 : _GEN_18702; // @[sequencer-master.scala 154:24]
  wire  _GEN_18951 = _T_335 ? _GEN_18943 : _GEN_18703; // @[sequencer-master.scala 154:24]
  wire  _GEN_18952 = _T_335 ? _GEN_18944 : _GEN_18704; // @[sequencer-master.scala 154:24]
  wire  _GEN_18953 = _T_335 ? _GEN_18945 : _GEN_18705; // @[sequencer-master.scala 154:24]
  wire  _GEN_18954 = _T_335 ? _GEN_18946 : _GEN_18706; // @[sequencer-master.scala 154:24]
  wire  _GEN_18955 = _T_335 ? _GEN_18947 : _GEN_18707; // @[sequencer-master.scala 154:24]
  wire  _GEN_18956 = _GEN_32729 | _GEN_18716; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18957 = _GEN_32730 | _GEN_18717; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18958 = _GEN_32731 | _GEN_18718; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18959 = _GEN_32732 | _GEN_18719; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18960 = _GEN_32733 | _GEN_18720; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18961 = _GEN_32734 | _GEN_18721; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18962 = _GEN_32735 | _GEN_18722; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18963 = _GEN_32736 | _GEN_18723; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_18964 = _T_357 ? _GEN_18956 : _GEN_18716; // @[sequencer-master.scala 154:24]
  wire  _GEN_18965 = _T_357 ? _GEN_18957 : _GEN_18717; // @[sequencer-master.scala 154:24]
  wire  _GEN_18966 = _T_357 ? _GEN_18958 : _GEN_18718; // @[sequencer-master.scala 154:24]
  wire  _GEN_18967 = _T_357 ? _GEN_18959 : _GEN_18719; // @[sequencer-master.scala 154:24]
  wire  _GEN_18968 = _T_357 ? _GEN_18960 : _GEN_18720; // @[sequencer-master.scala 154:24]
  wire  _GEN_18969 = _T_357 ? _GEN_18961 : _GEN_18721; // @[sequencer-master.scala 154:24]
  wire  _GEN_18970 = _T_357 ? _GEN_18962 : _GEN_18722; // @[sequencer-master.scala 154:24]
  wire  _GEN_18971 = _T_357 ? _GEN_18963 : _GEN_18723; // @[sequencer-master.scala 154:24]
  wire [1:0] _e_tail_rports_9 = {{1'd0}, _T_1623}; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18972 = 3'h0 == tail ? _e_tail_rports_9 : _GEN_18202; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18973 = 3'h1 == tail ? _e_tail_rports_9 : _GEN_18203; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18974 = 3'h2 == tail ? _e_tail_rports_9 : _GEN_18204; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18975 = 3'h3 == tail ? _e_tail_rports_9 : _GEN_18205; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18976 = 3'h4 == tail ? _e_tail_rports_9 : _GEN_18206; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18977 = 3'h5 == tail ? _e_tail_rports_9 : _GEN_18207; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18978 = 3'h6 == tail ? _e_tail_rports_9 : _GEN_18208; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_18979 = 3'h7 == tail ? _e_tail_rports_9 : _GEN_18209; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_18980 = 3'h0 == tail ? 4'h0 : _GEN_18210; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18981 = 3'h1 == tail ? 4'h0 : _GEN_18211; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18982 = 3'h2 == tail ? 4'h0 : _GEN_18212; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18983 = 3'h3 == tail ? 4'h0 : _GEN_18213; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18984 = 3'h4 == tail ? 4'h0 : _GEN_18214; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18985 = 3'h5 == tail ? 4'h0 : _GEN_18215; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18986 = 3'h6 == tail ? 4'h0 : _GEN_18216; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_18987 = 3'h7 == tail ? 4'h0 : _GEN_18217; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_18988 = 3'h0 == tail ? 3'h0 : _GEN_18218; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18989 = 3'h1 == tail ? 3'h0 : _GEN_18219; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18990 = 3'h2 == tail ? 3'h0 : _GEN_18220; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18991 = 3'h3 == tail ? 3'h0 : _GEN_18221; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18992 = 3'h4 == tail ? 3'h0 : _GEN_18222; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18993 = 3'h5 == tail ? 3'h0 : _GEN_18223; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18994 = 3'h6 == tail ? 3'h0 : _GEN_18224; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_18995 = 3'h7 == tail ? 3'h0 : _GEN_18225; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_19012 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18564; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19013 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18565; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19014 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18566; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19015 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18567; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19016 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18568; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19017 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18569; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19018 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18570; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19019 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18571; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19020 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18796; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19021 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18797; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19022 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18798; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19023 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18799; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19024 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18800; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19025 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18801; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19026 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18802; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19027 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18803; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19028 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18260; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19029 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18261; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19030 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18262; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19031 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18263; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19032 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18264; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19033 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18265; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19034 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18266; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19035 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18267; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19036 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18268; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19037 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18269; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19038 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18270; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19039 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18271; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19040 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18272; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19041 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18273; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19042 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18274; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19043 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18275; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19044 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18276; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19045 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18277; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19046 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18278; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19047 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18279; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19048 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18280; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19049 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18281; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19050 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18282; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19051 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18283; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19060 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18852; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19061 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18853; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19062 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18854; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19063 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18855; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19064 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18856; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19065 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18857; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19066 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18858; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19067 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18859; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19068 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18300; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19069 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18301; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19070 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18302; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19071 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18303; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19072 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18304; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19073 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18305; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19074 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18306; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19075 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18307; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19076 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18308; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19077 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18309; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19078 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18310; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19079 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18311; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19080 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18312; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19081 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18313; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19082 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18314; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19083 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18315; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19084 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18868; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19085 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18869; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19086 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18870; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19087 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18871; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19088 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18872; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19089 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18873; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19090 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18874; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19091 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18875; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19092 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18324; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19093 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18325; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19094 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18326; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19095 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18327; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19096 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18328; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19097 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18329; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19098 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18330; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19099 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18331; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19100 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18332; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19101 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18333; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19102 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18334; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19103 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18335; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19104 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18336; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19105 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18337; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19106 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18338; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19107 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18339; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19108 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18884; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19109 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18885; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19110 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18886; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19111 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18887; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19112 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18888; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19113 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18889; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19114 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18890; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19115 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18891; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19116 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18348; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19117 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18349; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19118 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18350; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19119 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18351; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19120 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18352; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19121 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18353; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19122 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18354; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19123 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18355; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19124 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18356; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19125 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18357; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19126 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18358; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19127 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18359; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19128 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18360; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19129 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18361; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19130 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18362; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19131 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18363; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19132 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18900; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19133 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18901; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19134 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18902; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19135 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18903; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19136 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18904; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19137 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18905; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19138 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18906; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19139 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18907; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19140 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18372; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19141 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18373; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19142 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18374; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19143 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18375; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19144 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18376; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19145 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18377; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19146 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18378; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19147 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18379; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19148 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18380; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19149 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18381; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19150 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18382; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19151 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18383; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19152 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18384; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19153 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18385; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19154 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18386; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19155 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18387; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19156 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18916; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19157 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18917; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19158 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18918; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19159 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18919; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19160 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18920; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19161 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18921; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19162 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18922; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19163 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18923; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19164 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18396; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19165 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18397; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19166 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18398; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19167 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18399; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19168 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18400; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19169 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18401; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19170 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18402; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19171 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18403; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19172 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18404; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19173 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18405; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19174 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18406; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19175 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18407; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19176 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18408; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19177 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18409; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19178 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18410; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19179 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18411; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19180 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18932; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19181 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18933; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19182 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18934; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19183 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18935; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19184 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18936; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19185 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18937; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19186 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18938; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19187 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18939; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19188 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18420; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19189 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18421; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19190 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18422; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19191 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18423; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19192 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18424; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19193 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18425; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19194 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18426; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19195 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18427; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19196 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18428; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19197 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18429; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19198 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18430; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19199 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18431; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19200 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18432; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19201 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18433; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19202 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18434; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19203 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18435; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19204 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18948; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19205 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18949; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19206 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18950; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19207 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18951; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19208 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18952; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19209 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18953; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19210 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18954; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19211 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18955; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19212 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18444; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19213 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18445; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19214 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18446; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19215 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18447; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19216 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18448; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19217 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18449; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19218 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18450; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19219 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18451; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19220 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18452; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19221 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18453; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19222 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18454; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19223 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18455; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19224 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18456; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19225 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18457; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19226 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18458; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19227 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18459; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19228 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18964; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19229 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18965; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19230 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18966; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19231 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18967; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19232 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18968; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19233 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18969; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19234 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18970; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19235 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18971; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19236 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18468; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19237 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18469; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19238 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18470; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19239 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18471; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19240 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18472; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19241 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18473; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19242 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18474; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19243 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18475; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19244 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18476; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19245 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18477; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19246 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18478; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19247 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18479; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19248 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18480; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19249 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18481; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19250 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18482; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19251 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18483; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19252 = 3'h0 == _T_1645 ? 1'h0 : _GEN_18484; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19253 = 3'h1 == _T_1645 ? 1'h0 : _GEN_18485; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19254 = 3'h2 == _T_1645 ? 1'h0 : _GEN_18486; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19255 = 3'h3 == _T_1645 ? 1'h0 : _GEN_18487; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19256 = 3'h4 == _T_1645 ? 1'h0 : _GEN_18488; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19257 = 3'h5 == _T_1645 ? 1'h0 : _GEN_18489; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19258 = 3'h6 == _T_1645 ? 1'h0 : _GEN_18490; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19259 = 3'h7 == _T_1645 ? 1'h0 : _GEN_18491; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19268 = _GEN_34121 | e_0_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19269 = _GEN_34122 | e_1_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19270 = _GEN_34123 | e_2_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19271 = _GEN_34124 | e_3_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19272 = _GEN_34125 | e_4_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19273 = _GEN_34126 | e_5_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19274 = _GEN_34127 | e_6_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19275 = _GEN_34128 | e_7_active_vcu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_19276 = 3'h0 == _T_1645 ? io_op_bits_fn_union : _GEN_18508; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19277 = 3'h1 == _T_1645 ? io_op_bits_fn_union : _GEN_18509; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19278 = 3'h2 == _T_1645 ? io_op_bits_fn_union : _GEN_18510; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19279 = 3'h3 == _T_1645 ? io_op_bits_fn_union : _GEN_18511; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19280 = 3'h4 == _T_1645 ? io_op_bits_fn_union : _GEN_18512; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19281 = 3'h5 == _T_1645 ? io_op_bits_fn_union : _GEN_18513; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19282 = 3'h6 == _T_1645 ? io_op_bits_fn_union : _GEN_18514; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19283 = 3'h7 == _T_1645 ? io_op_bits_fn_union : _GEN_18515; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [1:0] _GEN_19284 = 3'h0 == _T_1645 ? 2'h0 : _GEN_18972; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19285 = 3'h1 == _T_1645 ? 2'h0 : _GEN_18973; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19286 = 3'h2 == _T_1645 ? 2'h0 : _GEN_18974; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19287 = 3'h3 == _T_1645 ? 2'h0 : _GEN_18975; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19288 = 3'h4 == _T_1645 ? 2'h0 : _GEN_18976; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19289 = 3'h5 == _T_1645 ? 2'h0 : _GEN_18977; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19290 = 3'h6 == _T_1645 ? 2'h0 : _GEN_18978; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_19291 = 3'h7 == _T_1645 ? 2'h0 : _GEN_18979; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_19292 = 3'h0 == _T_1645 ? 4'h0 : _GEN_18980; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19293 = 3'h1 == _T_1645 ? 4'h0 : _GEN_18981; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19294 = 3'h2 == _T_1645 ? 4'h0 : _GEN_18982; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19295 = 3'h3 == _T_1645 ? 4'h0 : _GEN_18983; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19296 = 3'h4 == _T_1645 ? 4'h0 : _GEN_18984; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19297 = 3'h5 == _T_1645 ? 4'h0 : _GEN_18985; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19298 = 3'h6 == _T_1645 ? 4'h0 : _GEN_18986; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_19299 = 3'h7 == _T_1645 ? 4'h0 : _GEN_18987; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_19300 = 3'h0 == _T_1645 ? 3'h0 : _GEN_18988; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19301 = 3'h1 == _T_1645 ? 3'h0 : _GEN_18989; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19302 = 3'h2 == _T_1645 ? 3'h0 : _GEN_18990; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19303 = 3'h3 == _T_1645 ? 3'h0 : _GEN_18991; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19304 = 3'h4 == _T_1645 ? 3'h0 : _GEN_18992; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19305 = 3'h5 == _T_1645 ? 3'h0 : _GEN_18993; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19306 = 3'h6 == _T_1645 ? 3'h0 : _GEN_18994; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_19307 = 3'h7 == _T_1645 ? 3'h0 : _GEN_18995; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_19308 = _GEN_34121 | _GEN_19068; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19309 = _GEN_34122 | _GEN_19069; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19310 = _GEN_34123 | _GEN_19070; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19311 = _GEN_34124 | _GEN_19071; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19312 = _GEN_34125 | _GEN_19072; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19313 = _GEN_34126 | _GEN_19073; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19314 = _GEN_34127 | _GEN_19074; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19315 = _GEN_34128 | _GEN_19075; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19316 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19308 : _GEN_19068; // @[sequencer-master.scala 161:86]
  wire  _GEN_19317 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19309 : _GEN_19069; // @[sequencer-master.scala 161:86]
  wire  _GEN_19318 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19310 : _GEN_19070; // @[sequencer-master.scala 161:86]
  wire  _GEN_19319 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19311 : _GEN_19071; // @[sequencer-master.scala 161:86]
  wire  _GEN_19320 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19312 : _GEN_19072; // @[sequencer-master.scala 161:86]
  wire  _GEN_19321 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19313 : _GEN_19073; // @[sequencer-master.scala 161:86]
  wire  _GEN_19322 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19314 : _GEN_19074; // @[sequencer-master.scala 161:86]
  wire  _GEN_19323 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_19315 : _GEN_19075; // @[sequencer-master.scala 161:86]
  wire  _GEN_19324 = _GEN_34121 | _GEN_19092; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19325 = _GEN_34122 | _GEN_19093; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19326 = _GEN_34123 | _GEN_19094; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19327 = _GEN_34124 | _GEN_19095; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19328 = _GEN_34125 | _GEN_19096; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19329 = _GEN_34126 | _GEN_19097; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19330 = _GEN_34127 | _GEN_19098; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19331 = _GEN_34128 | _GEN_19099; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19332 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19324 : _GEN_19092; // @[sequencer-master.scala 161:86]
  wire  _GEN_19333 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19325 : _GEN_19093; // @[sequencer-master.scala 161:86]
  wire  _GEN_19334 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19326 : _GEN_19094; // @[sequencer-master.scala 161:86]
  wire  _GEN_19335 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19327 : _GEN_19095; // @[sequencer-master.scala 161:86]
  wire  _GEN_19336 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19328 : _GEN_19096; // @[sequencer-master.scala 161:86]
  wire  _GEN_19337 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19329 : _GEN_19097; // @[sequencer-master.scala 161:86]
  wire  _GEN_19338 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19330 : _GEN_19098; // @[sequencer-master.scala 161:86]
  wire  _GEN_19339 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_19331 : _GEN_19099; // @[sequencer-master.scala 161:86]
  wire  _GEN_19340 = _GEN_34121 | _GEN_19116; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19341 = _GEN_34122 | _GEN_19117; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19342 = _GEN_34123 | _GEN_19118; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19343 = _GEN_34124 | _GEN_19119; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19344 = _GEN_34125 | _GEN_19120; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19345 = _GEN_34126 | _GEN_19121; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19346 = _GEN_34127 | _GEN_19122; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19347 = _GEN_34128 | _GEN_19123; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19348 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19340 : _GEN_19116; // @[sequencer-master.scala 161:86]
  wire  _GEN_19349 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19341 : _GEN_19117; // @[sequencer-master.scala 161:86]
  wire  _GEN_19350 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19342 : _GEN_19118; // @[sequencer-master.scala 161:86]
  wire  _GEN_19351 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19343 : _GEN_19119; // @[sequencer-master.scala 161:86]
  wire  _GEN_19352 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19344 : _GEN_19120; // @[sequencer-master.scala 161:86]
  wire  _GEN_19353 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19345 : _GEN_19121; // @[sequencer-master.scala 161:86]
  wire  _GEN_19354 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19346 : _GEN_19122; // @[sequencer-master.scala 161:86]
  wire  _GEN_19355 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_19347 : _GEN_19123; // @[sequencer-master.scala 161:86]
  wire  _GEN_19356 = _GEN_34121 | _GEN_19140; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19357 = _GEN_34122 | _GEN_19141; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19358 = _GEN_34123 | _GEN_19142; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19359 = _GEN_34124 | _GEN_19143; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19360 = _GEN_34125 | _GEN_19144; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19361 = _GEN_34126 | _GEN_19145; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19362 = _GEN_34127 | _GEN_19146; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19363 = _GEN_34128 | _GEN_19147; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19364 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19356 : _GEN_19140; // @[sequencer-master.scala 161:86]
  wire  _GEN_19365 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19357 : _GEN_19141; // @[sequencer-master.scala 161:86]
  wire  _GEN_19366 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19358 : _GEN_19142; // @[sequencer-master.scala 161:86]
  wire  _GEN_19367 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19359 : _GEN_19143; // @[sequencer-master.scala 161:86]
  wire  _GEN_19368 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19360 : _GEN_19144; // @[sequencer-master.scala 161:86]
  wire  _GEN_19369 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19361 : _GEN_19145; // @[sequencer-master.scala 161:86]
  wire  _GEN_19370 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19362 : _GEN_19146; // @[sequencer-master.scala 161:86]
  wire  _GEN_19371 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_19363 : _GEN_19147; // @[sequencer-master.scala 161:86]
  wire  _GEN_19372 = _GEN_34121 | _GEN_19164; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19373 = _GEN_34122 | _GEN_19165; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19374 = _GEN_34123 | _GEN_19166; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19375 = _GEN_34124 | _GEN_19167; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19376 = _GEN_34125 | _GEN_19168; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19377 = _GEN_34126 | _GEN_19169; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19378 = _GEN_34127 | _GEN_19170; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19379 = _GEN_34128 | _GEN_19171; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19380 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19372 : _GEN_19164; // @[sequencer-master.scala 161:86]
  wire  _GEN_19381 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19373 : _GEN_19165; // @[sequencer-master.scala 161:86]
  wire  _GEN_19382 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19374 : _GEN_19166; // @[sequencer-master.scala 161:86]
  wire  _GEN_19383 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19375 : _GEN_19167; // @[sequencer-master.scala 161:86]
  wire  _GEN_19384 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19376 : _GEN_19168; // @[sequencer-master.scala 161:86]
  wire  _GEN_19385 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19377 : _GEN_19169; // @[sequencer-master.scala 161:86]
  wire  _GEN_19386 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19378 : _GEN_19170; // @[sequencer-master.scala 161:86]
  wire  _GEN_19387 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_19379 : _GEN_19171; // @[sequencer-master.scala 161:86]
  wire  _GEN_19388 = _GEN_34121 | _GEN_19188; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19389 = _GEN_34122 | _GEN_19189; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19390 = _GEN_34123 | _GEN_19190; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19391 = _GEN_34124 | _GEN_19191; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19392 = _GEN_34125 | _GEN_19192; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19393 = _GEN_34126 | _GEN_19193; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19394 = _GEN_34127 | _GEN_19194; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19395 = _GEN_34128 | _GEN_19195; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19396 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19388 : _GEN_19188; // @[sequencer-master.scala 161:86]
  wire  _GEN_19397 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19389 : _GEN_19189; // @[sequencer-master.scala 161:86]
  wire  _GEN_19398 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19390 : _GEN_19190; // @[sequencer-master.scala 161:86]
  wire  _GEN_19399 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19391 : _GEN_19191; // @[sequencer-master.scala 161:86]
  wire  _GEN_19400 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19392 : _GEN_19192; // @[sequencer-master.scala 161:86]
  wire  _GEN_19401 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19393 : _GEN_19193; // @[sequencer-master.scala 161:86]
  wire  _GEN_19402 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19394 : _GEN_19194; // @[sequencer-master.scala 161:86]
  wire  _GEN_19403 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_19395 : _GEN_19195; // @[sequencer-master.scala 161:86]
  wire  _GEN_19404 = _GEN_34121 | _GEN_19212; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19405 = _GEN_34122 | _GEN_19213; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19406 = _GEN_34123 | _GEN_19214; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19407 = _GEN_34124 | _GEN_19215; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19408 = _GEN_34125 | _GEN_19216; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19409 = _GEN_34126 | _GEN_19217; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19410 = _GEN_34127 | _GEN_19218; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19411 = _GEN_34128 | _GEN_19219; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19412 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19404 : _GEN_19212; // @[sequencer-master.scala 161:86]
  wire  _GEN_19413 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19405 : _GEN_19213; // @[sequencer-master.scala 161:86]
  wire  _GEN_19414 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19406 : _GEN_19214; // @[sequencer-master.scala 161:86]
  wire  _GEN_19415 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19407 : _GEN_19215; // @[sequencer-master.scala 161:86]
  wire  _GEN_19416 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19408 : _GEN_19216; // @[sequencer-master.scala 161:86]
  wire  _GEN_19417 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19409 : _GEN_19217; // @[sequencer-master.scala 161:86]
  wire  _GEN_19418 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19410 : _GEN_19218; // @[sequencer-master.scala 161:86]
  wire  _GEN_19419 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_19411 : _GEN_19219; // @[sequencer-master.scala 161:86]
  wire  _GEN_19420 = _GEN_34121 | _GEN_19236; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19421 = _GEN_34122 | _GEN_19237; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19422 = _GEN_34123 | _GEN_19238; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19423 = _GEN_34124 | _GEN_19239; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19424 = _GEN_34125 | _GEN_19240; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19425 = _GEN_34126 | _GEN_19241; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19426 = _GEN_34127 | _GEN_19242; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19427 = _GEN_34128 | _GEN_19243; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_19428 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19420 : _GEN_19236; // @[sequencer-master.scala 161:86]
  wire  _GEN_19429 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19421 : _GEN_19237; // @[sequencer-master.scala 161:86]
  wire  _GEN_19430 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19422 : _GEN_19238; // @[sequencer-master.scala 161:86]
  wire  _GEN_19431 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19423 : _GEN_19239; // @[sequencer-master.scala 161:86]
  wire  _GEN_19432 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19424 : _GEN_19240; // @[sequencer-master.scala 161:86]
  wire  _GEN_19433 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19425 : _GEN_19241; // @[sequencer-master.scala 161:86]
  wire  _GEN_19434 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19426 : _GEN_19242; // @[sequencer-master.scala 161:86]
  wire  _GEN_19435 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_19427 : _GEN_19243; // @[sequencer-master.scala 161:86]
  wire  _GEN_19436 = _GEN_34121 | _GEN_19076; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19437 = _GEN_34122 | _GEN_19077; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19438 = _GEN_34123 | _GEN_19078; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19439 = _GEN_34124 | _GEN_19079; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19440 = _GEN_34125 | _GEN_19080; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19441 = _GEN_34126 | _GEN_19081; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19442 = _GEN_34127 | _GEN_19082; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19443 = _GEN_34128 | _GEN_19083; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19444 = _T_1442 ? _GEN_19436 : _GEN_19076; // @[sequencer-master.scala 168:32]
  wire  _GEN_19445 = _T_1442 ? _GEN_19437 : _GEN_19077; // @[sequencer-master.scala 168:32]
  wire  _GEN_19446 = _T_1442 ? _GEN_19438 : _GEN_19078; // @[sequencer-master.scala 168:32]
  wire  _GEN_19447 = _T_1442 ? _GEN_19439 : _GEN_19079; // @[sequencer-master.scala 168:32]
  wire  _GEN_19448 = _T_1442 ? _GEN_19440 : _GEN_19080; // @[sequencer-master.scala 168:32]
  wire  _GEN_19449 = _T_1442 ? _GEN_19441 : _GEN_19081; // @[sequencer-master.scala 168:32]
  wire  _GEN_19450 = _T_1442 ? _GEN_19442 : _GEN_19082; // @[sequencer-master.scala 168:32]
  wire  _GEN_19451 = _T_1442 ? _GEN_19443 : _GEN_19083; // @[sequencer-master.scala 168:32]
  wire  _GEN_19452 = _GEN_34121 | _GEN_19100; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19453 = _GEN_34122 | _GEN_19101; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19454 = _GEN_34123 | _GEN_19102; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19455 = _GEN_34124 | _GEN_19103; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19456 = _GEN_34125 | _GEN_19104; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19457 = _GEN_34126 | _GEN_19105; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19458 = _GEN_34127 | _GEN_19106; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19459 = _GEN_34128 | _GEN_19107; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19460 = _T_1464 ? _GEN_19452 : _GEN_19100; // @[sequencer-master.scala 168:32]
  wire  _GEN_19461 = _T_1464 ? _GEN_19453 : _GEN_19101; // @[sequencer-master.scala 168:32]
  wire  _GEN_19462 = _T_1464 ? _GEN_19454 : _GEN_19102; // @[sequencer-master.scala 168:32]
  wire  _GEN_19463 = _T_1464 ? _GEN_19455 : _GEN_19103; // @[sequencer-master.scala 168:32]
  wire  _GEN_19464 = _T_1464 ? _GEN_19456 : _GEN_19104; // @[sequencer-master.scala 168:32]
  wire  _GEN_19465 = _T_1464 ? _GEN_19457 : _GEN_19105; // @[sequencer-master.scala 168:32]
  wire  _GEN_19466 = _T_1464 ? _GEN_19458 : _GEN_19106; // @[sequencer-master.scala 168:32]
  wire  _GEN_19467 = _T_1464 ? _GEN_19459 : _GEN_19107; // @[sequencer-master.scala 168:32]
  wire  _GEN_19468 = _GEN_34121 | _GEN_19124; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19469 = _GEN_34122 | _GEN_19125; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19470 = _GEN_34123 | _GEN_19126; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19471 = _GEN_34124 | _GEN_19127; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19472 = _GEN_34125 | _GEN_19128; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19473 = _GEN_34126 | _GEN_19129; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19474 = _GEN_34127 | _GEN_19130; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19475 = _GEN_34128 | _GEN_19131; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19476 = _T_1486 ? _GEN_19468 : _GEN_19124; // @[sequencer-master.scala 168:32]
  wire  _GEN_19477 = _T_1486 ? _GEN_19469 : _GEN_19125; // @[sequencer-master.scala 168:32]
  wire  _GEN_19478 = _T_1486 ? _GEN_19470 : _GEN_19126; // @[sequencer-master.scala 168:32]
  wire  _GEN_19479 = _T_1486 ? _GEN_19471 : _GEN_19127; // @[sequencer-master.scala 168:32]
  wire  _GEN_19480 = _T_1486 ? _GEN_19472 : _GEN_19128; // @[sequencer-master.scala 168:32]
  wire  _GEN_19481 = _T_1486 ? _GEN_19473 : _GEN_19129; // @[sequencer-master.scala 168:32]
  wire  _GEN_19482 = _T_1486 ? _GEN_19474 : _GEN_19130; // @[sequencer-master.scala 168:32]
  wire  _GEN_19483 = _T_1486 ? _GEN_19475 : _GEN_19131; // @[sequencer-master.scala 168:32]
  wire  _GEN_19484 = _GEN_34121 | _GEN_19148; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19485 = _GEN_34122 | _GEN_19149; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19486 = _GEN_34123 | _GEN_19150; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19487 = _GEN_34124 | _GEN_19151; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19488 = _GEN_34125 | _GEN_19152; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19489 = _GEN_34126 | _GEN_19153; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19490 = _GEN_34127 | _GEN_19154; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19491 = _GEN_34128 | _GEN_19155; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19492 = _T_1508 ? _GEN_19484 : _GEN_19148; // @[sequencer-master.scala 168:32]
  wire  _GEN_19493 = _T_1508 ? _GEN_19485 : _GEN_19149; // @[sequencer-master.scala 168:32]
  wire  _GEN_19494 = _T_1508 ? _GEN_19486 : _GEN_19150; // @[sequencer-master.scala 168:32]
  wire  _GEN_19495 = _T_1508 ? _GEN_19487 : _GEN_19151; // @[sequencer-master.scala 168:32]
  wire  _GEN_19496 = _T_1508 ? _GEN_19488 : _GEN_19152; // @[sequencer-master.scala 168:32]
  wire  _GEN_19497 = _T_1508 ? _GEN_19489 : _GEN_19153; // @[sequencer-master.scala 168:32]
  wire  _GEN_19498 = _T_1508 ? _GEN_19490 : _GEN_19154; // @[sequencer-master.scala 168:32]
  wire  _GEN_19499 = _T_1508 ? _GEN_19491 : _GEN_19155; // @[sequencer-master.scala 168:32]
  wire  _GEN_19500 = _GEN_34121 | _GEN_19172; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19501 = _GEN_34122 | _GEN_19173; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19502 = _GEN_34123 | _GEN_19174; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19503 = _GEN_34124 | _GEN_19175; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19504 = _GEN_34125 | _GEN_19176; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19505 = _GEN_34126 | _GEN_19177; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19506 = _GEN_34127 | _GEN_19178; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19507 = _GEN_34128 | _GEN_19179; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19508 = _T_1530 ? _GEN_19500 : _GEN_19172; // @[sequencer-master.scala 168:32]
  wire  _GEN_19509 = _T_1530 ? _GEN_19501 : _GEN_19173; // @[sequencer-master.scala 168:32]
  wire  _GEN_19510 = _T_1530 ? _GEN_19502 : _GEN_19174; // @[sequencer-master.scala 168:32]
  wire  _GEN_19511 = _T_1530 ? _GEN_19503 : _GEN_19175; // @[sequencer-master.scala 168:32]
  wire  _GEN_19512 = _T_1530 ? _GEN_19504 : _GEN_19176; // @[sequencer-master.scala 168:32]
  wire  _GEN_19513 = _T_1530 ? _GEN_19505 : _GEN_19177; // @[sequencer-master.scala 168:32]
  wire  _GEN_19514 = _T_1530 ? _GEN_19506 : _GEN_19178; // @[sequencer-master.scala 168:32]
  wire  _GEN_19515 = _T_1530 ? _GEN_19507 : _GEN_19179; // @[sequencer-master.scala 168:32]
  wire  _GEN_19516 = _GEN_34121 | _GEN_19196; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19517 = _GEN_34122 | _GEN_19197; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19518 = _GEN_34123 | _GEN_19198; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19519 = _GEN_34124 | _GEN_19199; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19520 = _GEN_34125 | _GEN_19200; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19521 = _GEN_34126 | _GEN_19201; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19522 = _GEN_34127 | _GEN_19202; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19523 = _GEN_34128 | _GEN_19203; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19524 = _T_1552 ? _GEN_19516 : _GEN_19196; // @[sequencer-master.scala 168:32]
  wire  _GEN_19525 = _T_1552 ? _GEN_19517 : _GEN_19197; // @[sequencer-master.scala 168:32]
  wire  _GEN_19526 = _T_1552 ? _GEN_19518 : _GEN_19198; // @[sequencer-master.scala 168:32]
  wire  _GEN_19527 = _T_1552 ? _GEN_19519 : _GEN_19199; // @[sequencer-master.scala 168:32]
  wire  _GEN_19528 = _T_1552 ? _GEN_19520 : _GEN_19200; // @[sequencer-master.scala 168:32]
  wire  _GEN_19529 = _T_1552 ? _GEN_19521 : _GEN_19201; // @[sequencer-master.scala 168:32]
  wire  _GEN_19530 = _T_1552 ? _GEN_19522 : _GEN_19202; // @[sequencer-master.scala 168:32]
  wire  _GEN_19531 = _T_1552 ? _GEN_19523 : _GEN_19203; // @[sequencer-master.scala 168:32]
  wire  _GEN_19532 = _GEN_34121 | _GEN_19220; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19533 = _GEN_34122 | _GEN_19221; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19534 = _GEN_34123 | _GEN_19222; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19535 = _GEN_34124 | _GEN_19223; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19536 = _GEN_34125 | _GEN_19224; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19537 = _GEN_34126 | _GEN_19225; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19538 = _GEN_34127 | _GEN_19226; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19539 = _GEN_34128 | _GEN_19227; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19540 = _T_1574 ? _GEN_19532 : _GEN_19220; // @[sequencer-master.scala 168:32]
  wire  _GEN_19541 = _T_1574 ? _GEN_19533 : _GEN_19221; // @[sequencer-master.scala 168:32]
  wire  _GEN_19542 = _T_1574 ? _GEN_19534 : _GEN_19222; // @[sequencer-master.scala 168:32]
  wire  _GEN_19543 = _T_1574 ? _GEN_19535 : _GEN_19223; // @[sequencer-master.scala 168:32]
  wire  _GEN_19544 = _T_1574 ? _GEN_19536 : _GEN_19224; // @[sequencer-master.scala 168:32]
  wire  _GEN_19545 = _T_1574 ? _GEN_19537 : _GEN_19225; // @[sequencer-master.scala 168:32]
  wire  _GEN_19546 = _T_1574 ? _GEN_19538 : _GEN_19226; // @[sequencer-master.scala 168:32]
  wire  _GEN_19547 = _T_1574 ? _GEN_19539 : _GEN_19227; // @[sequencer-master.scala 168:32]
  wire  _GEN_19548 = _GEN_34121 | _GEN_19244; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19549 = _GEN_34122 | _GEN_19245; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19550 = _GEN_34123 | _GEN_19246; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19551 = _GEN_34124 | _GEN_19247; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19552 = _GEN_34125 | _GEN_19248; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19553 = _GEN_34126 | _GEN_19249; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19554 = _GEN_34127 | _GEN_19250; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19555 = _GEN_34128 | _GEN_19251; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_19556 = _T_1596 ? _GEN_19548 : _GEN_19244; // @[sequencer-master.scala 168:32]
  wire  _GEN_19557 = _T_1596 ? _GEN_19549 : _GEN_19245; // @[sequencer-master.scala 168:32]
  wire  _GEN_19558 = _T_1596 ? _GEN_19550 : _GEN_19246; // @[sequencer-master.scala 168:32]
  wire  _GEN_19559 = _T_1596 ? _GEN_19551 : _GEN_19247; // @[sequencer-master.scala 168:32]
  wire  _GEN_19560 = _T_1596 ? _GEN_19552 : _GEN_19248; // @[sequencer-master.scala 168:32]
  wire  _GEN_19561 = _T_1596 ? _GEN_19553 : _GEN_19249; // @[sequencer-master.scala 168:32]
  wire  _GEN_19562 = _T_1596 ? _GEN_19554 : _GEN_19250; // @[sequencer-master.scala 168:32]
  wire  _GEN_19563 = _T_1596 ? _GEN_19555 : _GEN_19251; // @[sequencer-master.scala 168:32]
  wire  _GEN_36426 = 3'h0 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36427 = 3'h1 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36428 = 3'h2 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36429 = 3'h3 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36430 = 3'h4 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36431 = 3'h5 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36432 = 3'h6 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36433 = 3'h7 == _T_1647; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_19580 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19012; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19581 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19013; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19582 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19014; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19583 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19015; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19584 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19016; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19585 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19017; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19586 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19018; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19587 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19019; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_19588 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19020; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19589 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19021; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19590 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19022; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19591 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19023; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19592 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19024; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19593 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19025; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19594 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19026; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19595 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19027; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_19596 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19028; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19597 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19029; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19598 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19030; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19599 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19031; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19600 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19032; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19601 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19033; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19602 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19034; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19603 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19035; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_19604 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19036; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19605 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19037; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19606 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19038; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19607 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19039; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19608 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19040; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19609 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19041; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19610 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19042; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19611 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19043; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_19612 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19044; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19613 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19045; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19614 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19046; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19615 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19047; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19616 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19048; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19617 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19049; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19618 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19050; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19619 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19051; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_19628 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19060; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19629 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19061; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19630 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19062; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19631 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19063; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19632 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19064; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19633 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19065; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19634 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19066; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19635 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19067; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19636 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19316; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19637 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19317; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19638 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19318; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19639 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19319; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19640 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19320; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19641 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19321; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19642 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19322; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19643 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19323; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19644 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19444; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19645 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19445; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19646 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19446; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19647 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19447; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19648 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19448; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19649 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19449; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19650 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19450; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19651 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19451; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19652 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19084; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19653 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19085; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19654 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19086; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19655 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19087; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19656 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19088; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19657 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19089; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19658 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19090; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19659 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19091; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19660 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19332; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19661 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19333; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19662 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19334; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19663 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19335; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19664 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19336; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19665 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19337; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19666 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19338; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19667 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19339; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19668 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19460; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19669 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19461; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19670 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19462; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19671 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19463; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19672 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19464; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19673 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19465; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19674 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19466; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19675 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19467; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19676 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19108; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19677 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19109; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19678 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19110; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19679 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19111; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19680 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19112; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19681 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19113; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19682 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19114; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19683 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19115; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19684 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19348; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19685 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19349; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19686 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19350; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19687 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19351; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19688 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19352; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19689 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19353; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19690 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19354; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19691 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19355; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19692 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19476; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19693 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19477; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19694 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19478; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19695 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19479; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19696 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19480; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19697 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19481; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19698 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19482; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19699 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19483; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19700 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19132; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19701 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19133; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19702 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19134; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19703 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19135; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19704 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19136; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19705 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19137; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19706 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19138; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19707 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19139; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19708 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19364; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19709 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19365; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19710 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19366; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19711 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19367; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19712 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19368; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19713 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19369; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19714 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19370; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19715 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19371; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19716 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19492; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19717 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19493; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19718 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19494; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19719 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19495; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19720 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19496; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19721 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19497; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19722 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19498; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19723 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19499; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19724 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19156; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19725 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19157; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19726 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19158; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19727 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19159; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19728 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19160; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19729 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19161; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19730 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19162; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19731 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19163; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19732 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19380; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19733 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19381; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19734 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19382; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19735 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19383; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19736 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19384; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19737 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19385; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19738 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19386; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19739 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19387; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19740 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19508; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19741 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19509; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19742 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19510; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19743 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19511; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19744 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19512; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19745 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19513; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19746 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19514; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19747 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19515; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19748 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19180; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19749 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19181; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19750 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19182; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19751 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19183; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19752 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19184; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19753 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19185; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19754 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19186; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19755 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19187; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19756 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19396; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19757 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19397; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19758 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19398; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19759 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19399; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19760 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19400; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19761 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19401; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19762 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19402; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19763 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19403; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19764 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19524; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19765 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19525; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19766 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19526; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19767 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19527; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19768 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19528; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19769 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19529; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19770 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19530; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19771 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19531; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19772 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19204; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19773 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19205; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19774 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19206; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19775 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19207; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19776 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19208; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19777 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19209; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19778 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19210; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19779 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19211; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19780 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19412; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19781 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19413; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19782 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19414; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19783 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19415; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19784 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19416; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19785 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19417; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19786 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19418; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19787 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19419; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19788 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19540; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19789 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19541; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19790 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19542; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19791 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19543; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19792 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19544; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19793 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19545; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19794 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19546; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19795 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19547; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19796 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19228; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19797 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19229; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19798 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19230; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19799 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19231; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19800 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19232; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19801 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19233; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19802 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19234; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19803 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19235; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_19804 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19428; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19805 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19429; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19806 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19430; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19807 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19431; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19808 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19432; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19809 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19433; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19810 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19434; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19811 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19435; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_19812 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19556; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19813 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19557; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19814 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19558; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19815 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19559; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19816 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19560; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19817 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19561; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19818 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19562; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19819 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19563; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_19820 = 3'h0 == _T_1647 ? 1'h0 : _GEN_19252; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19821 = 3'h1 == _T_1647 ? 1'h0 : _GEN_19253; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19822 = 3'h2 == _T_1647 ? 1'h0 : _GEN_19254; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19823 = 3'h3 == _T_1647 ? 1'h0 : _GEN_19255; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19824 = 3'h4 == _T_1647 ? 1'h0 : _GEN_19256; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19825 = 3'h5 == _T_1647 ? 1'h0 : _GEN_19257; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19826 = 3'h6 == _T_1647 ? 1'h0 : _GEN_19258; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19827 = 3'h7 == _T_1647 ? 1'h0 : _GEN_19259; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_19836 = _GEN_36426 | e_0_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19837 = _GEN_36427 | e_1_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19838 = _GEN_36428 | e_2_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19839 = _GEN_36429 | e_3_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19840 = _GEN_36430 | e_4_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19841 = _GEN_36431 | e_5_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19842 = _GEN_36432 | e_6_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_19843 = _GEN_36433 | e_7_active_vsu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_19844 = 3'h0 == _T_1647 ? io_op_bits_fn_union : _GEN_19276; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19845 = 3'h1 == _T_1647 ? io_op_bits_fn_union : _GEN_19277; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19846 = 3'h2 == _T_1647 ? io_op_bits_fn_union : _GEN_19278; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19847 = 3'h3 == _T_1647 ? io_op_bits_fn_union : _GEN_19279; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19848 = 3'h4 == _T_1647 ? io_op_bits_fn_union : _GEN_19280; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19849 = 3'h5 == _T_1647 ? io_op_bits_fn_union : _GEN_19281; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19850 = 3'h6 == _T_1647 ? io_op_bits_fn_union : _GEN_19282; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_19851 = 3'h7 == _T_1647 ? io_op_bits_fn_union : _GEN_19283; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_19852 = 3'h0 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18556; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19853 = 3'h1 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18557; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19854 = 3'h2 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18558; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19855 = 3'h3 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18559; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19856 = 3'h4 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18560; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19857 = 3'h5 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18561; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19858 = 3'h6 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18562; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_19859 = 3'h7 == _T_1647 ? io_op_bits_base_vp_id : _GEN_18563; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19860 = 3'h0 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19580; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19861 = 3'h1 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19581; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19862 = 3'h2 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19582; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19863 = 3'h3 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19583; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19864 = 3'h4 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19584; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19865 = 3'h5 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19585; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19866 = 3'h6 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19586; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19867 = 3'h7 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_19587; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19868 = 3'h0 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18572; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19869 = 3'h1 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18573; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19870 = 3'h2 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18574; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19871 = 3'h3 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18575; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19872 = 3'h4 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18576; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19873 = 3'h5 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18577; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19874 = 3'h6 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18578; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19875 = 3'h7 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_18579; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19876 = 3'h0 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18580; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19877 = 3'h1 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18581; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19878 = 3'h2 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18582; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19879 = 3'h3 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18583; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19880 = 3'h4 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18584; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19881 = 3'h5 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18585; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19882 = 3'h6 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18586; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_19883 = 3'h7 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_18587; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_19884 = 3'h0 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18588; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19885 = 3'h1 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18589; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19886 = 3'h2 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18590; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19887 = 3'h3 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18591; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19888 = 3'h4 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18592; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19889 = 3'h5 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18593; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19890 = 3'h6 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18594; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_19891 = 3'h7 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_18595; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_19892 = io_op_bits_base_vp_valid ? _GEN_19852 : _GEN_18556; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19893 = io_op_bits_base_vp_valid ? _GEN_19853 : _GEN_18557; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19894 = io_op_bits_base_vp_valid ? _GEN_19854 : _GEN_18558; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19895 = io_op_bits_base_vp_valid ? _GEN_19855 : _GEN_18559; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19896 = io_op_bits_base_vp_valid ? _GEN_19856 : _GEN_18560; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19897 = io_op_bits_base_vp_valid ? _GEN_19857 : _GEN_18561; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19898 = io_op_bits_base_vp_valid ? _GEN_19858 : _GEN_18562; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_19899 = io_op_bits_base_vp_valid ? _GEN_19859 : _GEN_18563; // @[sequencer-master.scala 320:41]
  wire  _GEN_19900 = io_op_bits_base_vp_valid ? _GEN_19860 : _GEN_19580; // @[sequencer-master.scala 320:41]
  wire  _GEN_19901 = io_op_bits_base_vp_valid ? _GEN_19861 : _GEN_19581; // @[sequencer-master.scala 320:41]
  wire  _GEN_19902 = io_op_bits_base_vp_valid ? _GEN_19862 : _GEN_19582; // @[sequencer-master.scala 320:41]
  wire  _GEN_19903 = io_op_bits_base_vp_valid ? _GEN_19863 : _GEN_19583; // @[sequencer-master.scala 320:41]
  wire  _GEN_19904 = io_op_bits_base_vp_valid ? _GEN_19864 : _GEN_19584; // @[sequencer-master.scala 320:41]
  wire  _GEN_19905 = io_op_bits_base_vp_valid ? _GEN_19865 : _GEN_19585; // @[sequencer-master.scala 320:41]
  wire  _GEN_19906 = io_op_bits_base_vp_valid ? _GEN_19866 : _GEN_19586; // @[sequencer-master.scala 320:41]
  wire  _GEN_19907 = io_op_bits_base_vp_valid ? _GEN_19867 : _GEN_19587; // @[sequencer-master.scala 320:41]
  wire  _GEN_19908 = io_op_bits_base_vp_valid ? _GEN_19868 : _GEN_18572; // @[sequencer-master.scala 320:41]
  wire  _GEN_19909 = io_op_bits_base_vp_valid ? _GEN_19869 : _GEN_18573; // @[sequencer-master.scala 320:41]
  wire  _GEN_19910 = io_op_bits_base_vp_valid ? _GEN_19870 : _GEN_18574; // @[sequencer-master.scala 320:41]
  wire  _GEN_19911 = io_op_bits_base_vp_valid ? _GEN_19871 : _GEN_18575; // @[sequencer-master.scala 320:41]
  wire  _GEN_19912 = io_op_bits_base_vp_valid ? _GEN_19872 : _GEN_18576; // @[sequencer-master.scala 320:41]
  wire  _GEN_19913 = io_op_bits_base_vp_valid ? _GEN_19873 : _GEN_18577; // @[sequencer-master.scala 320:41]
  wire  _GEN_19914 = io_op_bits_base_vp_valid ? _GEN_19874 : _GEN_18578; // @[sequencer-master.scala 320:41]
  wire  _GEN_19915 = io_op_bits_base_vp_valid ? _GEN_19875 : _GEN_18579; // @[sequencer-master.scala 320:41]
  wire  _GEN_19916 = io_op_bits_base_vp_valid ? _GEN_19876 : _GEN_18580; // @[sequencer-master.scala 320:41]
  wire  _GEN_19917 = io_op_bits_base_vp_valid ? _GEN_19877 : _GEN_18581; // @[sequencer-master.scala 320:41]
  wire  _GEN_19918 = io_op_bits_base_vp_valid ? _GEN_19878 : _GEN_18582; // @[sequencer-master.scala 320:41]
  wire  _GEN_19919 = io_op_bits_base_vp_valid ? _GEN_19879 : _GEN_18583; // @[sequencer-master.scala 320:41]
  wire  _GEN_19920 = io_op_bits_base_vp_valid ? _GEN_19880 : _GEN_18584; // @[sequencer-master.scala 320:41]
  wire  _GEN_19921 = io_op_bits_base_vp_valid ? _GEN_19881 : _GEN_18585; // @[sequencer-master.scala 320:41]
  wire  _GEN_19922 = io_op_bits_base_vp_valid ? _GEN_19882 : _GEN_18586; // @[sequencer-master.scala 320:41]
  wire  _GEN_19923 = io_op_bits_base_vp_valid ? _GEN_19883 : _GEN_18587; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19924 = io_op_bits_base_vp_valid ? _GEN_19884 : _GEN_18588; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19925 = io_op_bits_base_vp_valid ? _GEN_19885 : _GEN_18589; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19926 = io_op_bits_base_vp_valid ? _GEN_19886 : _GEN_18590; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19927 = io_op_bits_base_vp_valid ? _GEN_19887 : _GEN_18591; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19928 = io_op_bits_base_vp_valid ? _GEN_19888 : _GEN_18592; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19929 = io_op_bits_base_vp_valid ? _GEN_19889 : _GEN_18593; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19930 = io_op_bits_base_vp_valid ? _GEN_19890 : _GEN_18594; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_19931 = io_op_bits_base_vp_valid ? _GEN_19891 : _GEN_18595; // @[sequencer-master.scala 320:41]
  wire  _GEN_19932 = _GEN_36426 | _GEN_19628; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19933 = _GEN_36427 | _GEN_19629; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19934 = _GEN_36428 | _GEN_19630; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19935 = _GEN_36429 | _GEN_19631; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19936 = _GEN_36430 | _GEN_19632; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19937 = _GEN_36431 | _GEN_19633; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19938 = _GEN_36432 | _GEN_19634; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19939 = _GEN_36433 | _GEN_19635; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19940 = _T_26 ? _GEN_19932 : _GEN_19628; // @[sequencer-master.scala 154:24]
  wire  _GEN_19941 = _T_26 ? _GEN_19933 : _GEN_19629; // @[sequencer-master.scala 154:24]
  wire  _GEN_19942 = _T_26 ? _GEN_19934 : _GEN_19630; // @[sequencer-master.scala 154:24]
  wire  _GEN_19943 = _T_26 ? _GEN_19935 : _GEN_19631; // @[sequencer-master.scala 154:24]
  wire  _GEN_19944 = _T_26 ? _GEN_19936 : _GEN_19632; // @[sequencer-master.scala 154:24]
  wire  _GEN_19945 = _T_26 ? _GEN_19937 : _GEN_19633; // @[sequencer-master.scala 154:24]
  wire  _GEN_19946 = _T_26 ? _GEN_19938 : _GEN_19634; // @[sequencer-master.scala 154:24]
  wire  _GEN_19947 = _T_26 ? _GEN_19939 : _GEN_19635; // @[sequencer-master.scala 154:24]
  wire  _GEN_19948 = _GEN_36426 | _GEN_19652; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19949 = _GEN_36427 | _GEN_19653; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19950 = _GEN_36428 | _GEN_19654; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19951 = _GEN_36429 | _GEN_19655; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19952 = _GEN_36430 | _GEN_19656; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19953 = _GEN_36431 | _GEN_19657; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19954 = _GEN_36432 | _GEN_19658; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19955 = _GEN_36433 | _GEN_19659; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19956 = _T_48 ? _GEN_19948 : _GEN_19652; // @[sequencer-master.scala 154:24]
  wire  _GEN_19957 = _T_48 ? _GEN_19949 : _GEN_19653; // @[sequencer-master.scala 154:24]
  wire  _GEN_19958 = _T_48 ? _GEN_19950 : _GEN_19654; // @[sequencer-master.scala 154:24]
  wire  _GEN_19959 = _T_48 ? _GEN_19951 : _GEN_19655; // @[sequencer-master.scala 154:24]
  wire  _GEN_19960 = _T_48 ? _GEN_19952 : _GEN_19656; // @[sequencer-master.scala 154:24]
  wire  _GEN_19961 = _T_48 ? _GEN_19953 : _GEN_19657; // @[sequencer-master.scala 154:24]
  wire  _GEN_19962 = _T_48 ? _GEN_19954 : _GEN_19658; // @[sequencer-master.scala 154:24]
  wire  _GEN_19963 = _T_48 ? _GEN_19955 : _GEN_19659; // @[sequencer-master.scala 154:24]
  wire  _GEN_19964 = _GEN_36426 | _GEN_19676; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19965 = _GEN_36427 | _GEN_19677; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19966 = _GEN_36428 | _GEN_19678; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19967 = _GEN_36429 | _GEN_19679; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19968 = _GEN_36430 | _GEN_19680; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19969 = _GEN_36431 | _GEN_19681; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19970 = _GEN_36432 | _GEN_19682; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19971 = _GEN_36433 | _GEN_19683; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19972 = _T_70 ? _GEN_19964 : _GEN_19676; // @[sequencer-master.scala 154:24]
  wire  _GEN_19973 = _T_70 ? _GEN_19965 : _GEN_19677; // @[sequencer-master.scala 154:24]
  wire  _GEN_19974 = _T_70 ? _GEN_19966 : _GEN_19678; // @[sequencer-master.scala 154:24]
  wire  _GEN_19975 = _T_70 ? _GEN_19967 : _GEN_19679; // @[sequencer-master.scala 154:24]
  wire  _GEN_19976 = _T_70 ? _GEN_19968 : _GEN_19680; // @[sequencer-master.scala 154:24]
  wire  _GEN_19977 = _T_70 ? _GEN_19969 : _GEN_19681; // @[sequencer-master.scala 154:24]
  wire  _GEN_19978 = _T_70 ? _GEN_19970 : _GEN_19682; // @[sequencer-master.scala 154:24]
  wire  _GEN_19979 = _T_70 ? _GEN_19971 : _GEN_19683; // @[sequencer-master.scala 154:24]
  wire  _GEN_19980 = _GEN_36426 | _GEN_19700; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19981 = _GEN_36427 | _GEN_19701; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19982 = _GEN_36428 | _GEN_19702; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19983 = _GEN_36429 | _GEN_19703; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19984 = _GEN_36430 | _GEN_19704; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19985 = _GEN_36431 | _GEN_19705; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19986 = _GEN_36432 | _GEN_19706; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19987 = _GEN_36433 | _GEN_19707; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19988 = _T_92 ? _GEN_19980 : _GEN_19700; // @[sequencer-master.scala 154:24]
  wire  _GEN_19989 = _T_92 ? _GEN_19981 : _GEN_19701; // @[sequencer-master.scala 154:24]
  wire  _GEN_19990 = _T_92 ? _GEN_19982 : _GEN_19702; // @[sequencer-master.scala 154:24]
  wire  _GEN_19991 = _T_92 ? _GEN_19983 : _GEN_19703; // @[sequencer-master.scala 154:24]
  wire  _GEN_19992 = _T_92 ? _GEN_19984 : _GEN_19704; // @[sequencer-master.scala 154:24]
  wire  _GEN_19993 = _T_92 ? _GEN_19985 : _GEN_19705; // @[sequencer-master.scala 154:24]
  wire  _GEN_19994 = _T_92 ? _GEN_19986 : _GEN_19706; // @[sequencer-master.scala 154:24]
  wire  _GEN_19995 = _T_92 ? _GEN_19987 : _GEN_19707; // @[sequencer-master.scala 154:24]
  wire  _GEN_19996 = _GEN_36426 | _GEN_19724; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19997 = _GEN_36427 | _GEN_19725; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19998 = _GEN_36428 | _GEN_19726; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_19999 = _GEN_36429 | _GEN_19727; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20000 = _GEN_36430 | _GEN_19728; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20001 = _GEN_36431 | _GEN_19729; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20002 = _GEN_36432 | _GEN_19730; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20003 = _GEN_36433 | _GEN_19731; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20004 = _T_114 ? _GEN_19996 : _GEN_19724; // @[sequencer-master.scala 154:24]
  wire  _GEN_20005 = _T_114 ? _GEN_19997 : _GEN_19725; // @[sequencer-master.scala 154:24]
  wire  _GEN_20006 = _T_114 ? _GEN_19998 : _GEN_19726; // @[sequencer-master.scala 154:24]
  wire  _GEN_20007 = _T_114 ? _GEN_19999 : _GEN_19727; // @[sequencer-master.scala 154:24]
  wire  _GEN_20008 = _T_114 ? _GEN_20000 : _GEN_19728; // @[sequencer-master.scala 154:24]
  wire  _GEN_20009 = _T_114 ? _GEN_20001 : _GEN_19729; // @[sequencer-master.scala 154:24]
  wire  _GEN_20010 = _T_114 ? _GEN_20002 : _GEN_19730; // @[sequencer-master.scala 154:24]
  wire  _GEN_20011 = _T_114 ? _GEN_20003 : _GEN_19731; // @[sequencer-master.scala 154:24]
  wire  _GEN_20012 = _GEN_36426 | _GEN_19748; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20013 = _GEN_36427 | _GEN_19749; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20014 = _GEN_36428 | _GEN_19750; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20015 = _GEN_36429 | _GEN_19751; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20016 = _GEN_36430 | _GEN_19752; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20017 = _GEN_36431 | _GEN_19753; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20018 = _GEN_36432 | _GEN_19754; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20019 = _GEN_36433 | _GEN_19755; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20020 = _T_136 ? _GEN_20012 : _GEN_19748; // @[sequencer-master.scala 154:24]
  wire  _GEN_20021 = _T_136 ? _GEN_20013 : _GEN_19749; // @[sequencer-master.scala 154:24]
  wire  _GEN_20022 = _T_136 ? _GEN_20014 : _GEN_19750; // @[sequencer-master.scala 154:24]
  wire  _GEN_20023 = _T_136 ? _GEN_20015 : _GEN_19751; // @[sequencer-master.scala 154:24]
  wire  _GEN_20024 = _T_136 ? _GEN_20016 : _GEN_19752; // @[sequencer-master.scala 154:24]
  wire  _GEN_20025 = _T_136 ? _GEN_20017 : _GEN_19753; // @[sequencer-master.scala 154:24]
  wire  _GEN_20026 = _T_136 ? _GEN_20018 : _GEN_19754; // @[sequencer-master.scala 154:24]
  wire  _GEN_20027 = _T_136 ? _GEN_20019 : _GEN_19755; // @[sequencer-master.scala 154:24]
  wire  _GEN_20028 = _GEN_36426 | _GEN_19772; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20029 = _GEN_36427 | _GEN_19773; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20030 = _GEN_36428 | _GEN_19774; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20031 = _GEN_36429 | _GEN_19775; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20032 = _GEN_36430 | _GEN_19776; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20033 = _GEN_36431 | _GEN_19777; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20034 = _GEN_36432 | _GEN_19778; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20035 = _GEN_36433 | _GEN_19779; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20036 = _T_158 ? _GEN_20028 : _GEN_19772; // @[sequencer-master.scala 154:24]
  wire  _GEN_20037 = _T_158 ? _GEN_20029 : _GEN_19773; // @[sequencer-master.scala 154:24]
  wire  _GEN_20038 = _T_158 ? _GEN_20030 : _GEN_19774; // @[sequencer-master.scala 154:24]
  wire  _GEN_20039 = _T_158 ? _GEN_20031 : _GEN_19775; // @[sequencer-master.scala 154:24]
  wire  _GEN_20040 = _T_158 ? _GEN_20032 : _GEN_19776; // @[sequencer-master.scala 154:24]
  wire  _GEN_20041 = _T_158 ? _GEN_20033 : _GEN_19777; // @[sequencer-master.scala 154:24]
  wire  _GEN_20042 = _T_158 ? _GEN_20034 : _GEN_19778; // @[sequencer-master.scala 154:24]
  wire  _GEN_20043 = _T_158 ? _GEN_20035 : _GEN_19779; // @[sequencer-master.scala 154:24]
  wire  _GEN_20044 = _GEN_36426 | _GEN_19796; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20045 = _GEN_36427 | _GEN_19797; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20046 = _GEN_36428 | _GEN_19798; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20047 = _GEN_36429 | _GEN_19799; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20048 = _GEN_36430 | _GEN_19800; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20049 = _GEN_36431 | _GEN_19801; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20050 = _GEN_36432 | _GEN_19802; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20051 = _GEN_36433 | _GEN_19803; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20052 = _T_180 ? _GEN_20044 : _GEN_19796; // @[sequencer-master.scala 154:24]
  wire  _GEN_20053 = _T_180 ? _GEN_20045 : _GEN_19797; // @[sequencer-master.scala 154:24]
  wire  _GEN_20054 = _T_180 ? _GEN_20046 : _GEN_19798; // @[sequencer-master.scala 154:24]
  wire  _GEN_20055 = _T_180 ? _GEN_20047 : _GEN_19799; // @[sequencer-master.scala 154:24]
  wire  _GEN_20056 = _T_180 ? _GEN_20048 : _GEN_19800; // @[sequencer-master.scala 154:24]
  wire  _GEN_20057 = _T_180 ? _GEN_20049 : _GEN_19801; // @[sequencer-master.scala 154:24]
  wire  _GEN_20058 = _T_180 ? _GEN_20050 : _GEN_19802; // @[sequencer-master.scala 154:24]
  wire  _GEN_20059 = _T_180 ? _GEN_20051 : _GEN_19803; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_20060 = 3'h0 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18788; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20061 = 3'h1 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18789; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20062 = 3'h2 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18790; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20063 = 3'h3 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18791; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20064 = 3'h4 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18792; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20065 = 3'h5 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18793; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20066 = 3'h6 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18794; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20067 = 3'h7 == _T_1647 ? io_op_bits_base_vs2_id : _GEN_18795; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20068 = 3'h0 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19588; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20069 = 3'h1 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19589; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20070 = 3'h2 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19590; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20071 = 3'h3 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19591; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20072 = 3'h4 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19592; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20073 = 3'h5 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19593; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20074 = 3'h6 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19594; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20075 = 3'h7 == _T_1647 ? io_op_bits_base_vs2_valid : _GEN_19595; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20076 = 3'h0 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18804; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20077 = 3'h1 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18805; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20078 = 3'h2 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18806; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20079 = 3'h3 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18807; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20080 = 3'h4 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18808; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20081 = 3'h5 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18809; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20082 = 3'h6 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18810; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20083 = 3'h7 == _T_1647 ? io_op_bits_base_vs2_scalar : _GEN_18811; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20084 = 3'h0 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18812; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20085 = 3'h1 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18813; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20086 = 3'h2 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18814; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20087 = 3'h3 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18815; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20088 = 3'h4 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18816; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20089 = 3'h5 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18817; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20090 = 3'h6 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18818; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_20091 = 3'h7 == _T_1647 ? io_op_bits_base_vs2_pred : _GEN_18819; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20092 = 3'h0 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18820; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20093 = 3'h1 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18821; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20094 = 3'h2 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18822; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20095 = 3'h3 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18823; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20096 = 3'h4 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18824; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20097 = 3'h5 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18825; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20098 = 3'h6 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18826; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_20099 = 3'h7 == _T_1647 ? io_op_bits_base_vs2_prec : _GEN_18827; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_20100 = 3'h0 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18828; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20101 = 3'h1 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18829; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20102 = 3'h2 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18830; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20103 = 3'h3 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18831; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20104 = 3'h4 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18832; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20105 = 3'h5 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18833; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20106 = 3'h6 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18834; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_20107 = 3'h7 == _T_1647 ? io_op_bits_reg_vs2_id : _GEN_18835; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_20108 = 3'h0 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18836; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20109 = 3'h1 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18837; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20110 = 3'h2 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18838; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20111 = 3'h3 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18839; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20112 = 3'h4 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18840; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20113 = 3'h5 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18841; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20114 = 3'h6 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18842; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20115 = 3'h7 == _T_1647 ? io_op_bits_sreg_ss2 : _GEN_18843; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_20116 = _T_366 ? _GEN_20108 : _GEN_18836; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20117 = _T_366 ? _GEN_20109 : _GEN_18837; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20118 = _T_366 ? _GEN_20110 : _GEN_18838; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20119 = _T_366 ? _GEN_20111 : _GEN_18839; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20120 = _T_366 ? _GEN_20112 : _GEN_18840; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20121 = _T_366 ? _GEN_20113 : _GEN_18841; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20122 = _T_366 ? _GEN_20114 : _GEN_18842; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_20123 = _T_366 ? _GEN_20115 : _GEN_18843; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_20124 = io_op_bits_base_vs2_valid ? _GEN_20060 : _GEN_18788; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20125 = io_op_bits_base_vs2_valid ? _GEN_20061 : _GEN_18789; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20126 = io_op_bits_base_vs2_valid ? _GEN_20062 : _GEN_18790; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20127 = io_op_bits_base_vs2_valid ? _GEN_20063 : _GEN_18791; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20128 = io_op_bits_base_vs2_valid ? _GEN_20064 : _GEN_18792; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20129 = io_op_bits_base_vs2_valid ? _GEN_20065 : _GEN_18793; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20130 = io_op_bits_base_vs2_valid ? _GEN_20066 : _GEN_18794; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20131 = io_op_bits_base_vs2_valid ? _GEN_20067 : _GEN_18795; // @[sequencer-master.scala 328:47]
  wire  _GEN_20132 = io_op_bits_base_vs2_valid ? _GEN_20068 : _GEN_19588; // @[sequencer-master.scala 328:47]
  wire  _GEN_20133 = io_op_bits_base_vs2_valid ? _GEN_20069 : _GEN_19589; // @[sequencer-master.scala 328:47]
  wire  _GEN_20134 = io_op_bits_base_vs2_valid ? _GEN_20070 : _GEN_19590; // @[sequencer-master.scala 328:47]
  wire  _GEN_20135 = io_op_bits_base_vs2_valid ? _GEN_20071 : _GEN_19591; // @[sequencer-master.scala 328:47]
  wire  _GEN_20136 = io_op_bits_base_vs2_valid ? _GEN_20072 : _GEN_19592; // @[sequencer-master.scala 328:47]
  wire  _GEN_20137 = io_op_bits_base_vs2_valid ? _GEN_20073 : _GEN_19593; // @[sequencer-master.scala 328:47]
  wire  _GEN_20138 = io_op_bits_base_vs2_valid ? _GEN_20074 : _GEN_19594; // @[sequencer-master.scala 328:47]
  wire  _GEN_20139 = io_op_bits_base_vs2_valid ? _GEN_20075 : _GEN_19595; // @[sequencer-master.scala 328:47]
  wire  _GEN_20140 = io_op_bits_base_vs2_valid ? _GEN_20076 : _GEN_18804; // @[sequencer-master.scala 328:47]
  wire  _GEN_20141 = io_op_bits_base_vs2_valid ? _GEN_20077 : _GEN_18805; // @[sequencer-master.scala 328:47]
  wire  _GEN_20142 = io_op_bits_base_vs2_valid ? _GEN_20078 : _GEN_18806; // @[sequencer-master.scala 328:47]
  wire  _GEN_20143 = io_op_bits_base_vs2_valid ? _GEN_20079 : _GEN_18807; // @[sequencer-master.scala 328:47]
  wire  _GEN_20144 = io_op_bits_base_vs2_valid ? _GEN_20080 : _GEN_18808; // @[sequencer-master.scala 328:47]
  wire  _GEN_20145 = io_op_bits_base_vs2_valid ? _GEN_20081 : _GEN_18809; // @[sequencer-master.scala 328:47]
  wire  _GEN_20146 = io_op_bits_base_vs2_valid ? _GEN_20082 : _GEN_18810; // @[sequencer-master.scala 328:47]
  wire  _GEN_20147 = io_op_bits_base_vs2_valid ? _GEN_20083 : _GEN_18811; // @[sequencer-master.scala 328:47]
  wire  _GEN_20148 = io_op_bits_base_vs2_valid ? _GEN_20084 : _GEN_18812; // @[sequencer-master.scala 328:47]
  wire  _GEN_20149 = io_op_bits_base_vs2_valid ? _GEN_20085 : _GEN_18813; // @[sequencer-master.scala 328:47]
  wire  _GEN_20150 = io_op_bits_base_vs2_valid ? _GEN_20086 : _GEN_18814; // @[sequencer-master.scala 328:47]
  wire  _GEN_20151 = io_op_bits_base_vs2_valid ? _GEN_20087 : _GEN_18815; // @[sequencer-master.scala 328:47]
  wire  _GEN_20152 = io_op_bits_base_vs2_valid ? _GEN_20088 : _GEN_18816; // @[sequencer-master.scala 328:47]
  wire  _GEN_20153 = io_op_bits_base_vs2_valid ? _GEN_20089 : _GEN_18817; // @[sequencer-master.scala 328:47]
  wire  _GEN_20154 = io_op_bits_base_vs2_valid ? _GEN_20090 : _GEN_18818; // @[sequencer-master.scala 328:47]
  wire  _GEN_20155 = io_op_bits_base_vs2_valid ? _GEN_20091 : _GEN_18819; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20156 = io_op_bits_base_vs2_valid ? _GEN_20092 : _GEN_18820; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20157 = io_op_bits_base_vs2_valid ? _GEN_20093 : _GEN_18821; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20158 = io_op_bits_base_vs2_valid ? _GEN_20094 : _GEN_18822; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20159 = io_op_bits_base_vs2_valid ? _GEN_20095 : _GEN_18823; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20160 = io_op_bits_base_vs2_valid ? _GEN_20096 : _GEN_18824; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20161 = io_op_bits_base_vs2_valid ? _GEN_20097 : _GEN_18825; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20162 = io_op_bits_base_vs2_valid ? _GEN_20098 : _GEN_18826; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_20163 = io_op_bits_base_vs2_valid ? _GEN_20099 : _GEN_18827; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20164 = io_op_bits_base_vs2_valid ? _GEN_20100 : _GEN_18828; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20165 = io_op_bits_base_vs2_valid ? _GEN_20101 : _GEN_18829; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20166 = io_op_bits_base_vs2_valid ? _GEN_20102 : _GEN_18830; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20167 = io_op_bits_base_vs2_valid ? _GEN_20103 : _GEN_18831; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20168 = io_op_bits_base_vs2_valid ? _GEN_20104 : _GEN_18832; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20169 = io_op_bits_base_vs2_valid ? _GEN_20105 : _GEN_18833; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20170 = io_op_bits_base_vs2_valid ? _GEN_20106 : _GEN_18834; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_20171 = io_op_bits_base_vs2_valid ? _GEN_20107 : _GEN_18835; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20172 = io_op_bits_base_vs2_valid ? _GEN_20116 : _GEN_18836; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20173 = io_op_bits_base_vs2_valid ? _GEN_20117 : _GEN_18837; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20174 = io_op_bits_base_vs2_valid ? _GEN_20118 : _GEN_18838; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20175 = io_op_bits_base_vs2_valid ? _GEN_20119 : _GEN_18839; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20176 = io_op_bits_base_vs2_valid ? _GEN_20120 : _GEN_18840; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20177 = io_op_bits_base_vs2_valid ? _GEN_20121 : _GEN_18841; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20178 = io_op_bits_base_vs2_valid ? _GEN_20122 : _GEN_18842; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_20179 = io_op_bits_base_vs2_valid ? _GEN_20123 : _GEN_18843; // @[sequencer-master.scala 328:47]
  wire  _GEN_20180 = _GEN_36426 | _GEN_19940; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20181 = _GEN_36427 | _GEN_19941; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20182 = _GEN_36428 | _GEN_19942; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20183 = _GEN_36429 | _GEN_19943; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20184 = _GEN_36430 | _GEN_19944; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20185 = _GEN_36431 | _GEN_19945; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20186 = _GEN_36432 | _GEN_19946; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20187 = _GEN_36433 | _GEN_19947; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20188 = _T_380 ? _GEN_20180 : _GEN_19940; // @[sequencer-master.scala 154:24]
  wire  _GEN_20189 = _T_380 ? _GEN_20181 : _GEN_19941; // @[sequencer-master.scala 154:24]
  wire  _GEN_20190 = _T_380 ? _GEN_20182 : _GEN_19942; // @[sequencer-master.scala 154:24]
  wire  _GEN_20191 = _T_380 ? _GEN_20183 : _GEN_19943; // @[sequencer-master.scala 154:24]
  wire  _GEN_20192 = _T_380 ? _GEN_20184 : _GEN_19944; // @[sequencer-master.scala 154:24]
  wire  _GEN_20193 = _T_380 ? _GEN_20185 : _GEN_19945; // @[sequencer-master.scala 154:24]
  wire  _GEN_20194 = _T_380 ? _GEN_20186 : _GEN_19946; // @[sequencer-master.scala 154:24]
  wire  _GEN_20195 = _T_380 ? _GEN_20187 : _GEN_19947; // @[sequencer-master.scala 154:24]
  wire  _GEN_20196 = _GEN_36426 | _GEN_19956; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20197 = _GEN_36427 | _GEN_19957; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20198 = _GEN_36428 | _GEN_19958; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20199 = _GEN_36429 | _GEN_19959; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20200 = _GEN_36430 | _GEN_19960; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20201 = _GEN_36431 | _GEN_19961; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20202 = _GEN_36432 | _GEN_19962; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20203 = _GEN_36433 | _GEN_19963; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20204 = _T_402 ? _GEN_20196 : _GEN_19956; // @[sequencer-master.scala 154:24]
  wire  _GEN_20205 = _T_402 ? _GEN_20197 : _GEN_19957; // @[sequencer-master.scala 154:24]
  wire  _GEN_20206 = _T_402 ? _GEN_20198 : _GEN_19958; // @[sequencer-master.scala 154:24]
  wire  _GEN_20207 = _T_402 ? _GEN_20199 : _GEN_19959; // @[sequencer-master.scala 154:24]
  wire  _GEN_20208 = _T_402 ? _GEN_20200 : _GEN_19960; // @[sequencer-master.scala 154:24]
  wire  _GEN_20209 = _T_402 ? _GEN_20201 : _GEN_19961; // @[sequencer-master.scala 154:24]
  wire  _GEN_20210 = _T_402 ? _GEN_20202 : _GEN_19962; // @[sequencer-master.scala 154:24]
  wire  _GEN_20211 = _T_402 ? _GEN_20203 : _GEN_19963; // @[sequencer-master.scala 154:24]
  wire  _GEN_20212 = _GEN_36426 | _GEN_19972; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20213 = _GEN_36427 | _GEN_19973; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20214 = _GEN_36428 | _GEN_19974; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20215 = _GEN_36429 | _GEN_19975; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20216 = _GEN_36430 | _GEN_19976; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20217 = _GEN_36431 | _GEN_19977; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20218 = _GEN_36432 | _GEN_19978; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20219 = _GEN_36433 | _GEN_19979; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20220 = _T_424 ? _GEN_20212 : _GEN_19972; // @[sequencer-master.scala 154:24]
  wire  _GEN_20221 = _T_424 ? _GEN_20213 : _GEN_19973; // @[sequencer-master.scala 154:24]
  wire  _GEN_20222 = _T_424 ? _GEN_20214 : _GEN_19974; // @[sequencer-master.scala 154:24]
  wire  _GEN_20223 = _T_424 ? _GEN_20215 : _GEN_19975; // @[sequencer-master.scala 154:24]
  wire  _GEN_20224 = _T_424 ? _GEN_20216 : _GEN_19976; // @[sequencer-master.scala 154:24]
  wire  _GEN_20225 = _T_424 ? _GEN_20217 : _GEN_19977; // @[sequencer-master.scala 154:24]
  wire  _GEN_20226 = _T_424 ? _GEN_20218 : _GEN_19978; // @[sequencer-master.scala 154:24]
  wire  _GEN_20227 = _T_424 ? _GEN_20219 : _GEN_19979; // @[sequencer-master.scala 154:24]
  wire  _GEN_20228 = _GEN_36426 | _GEN_19988; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20229 = _GEN_36427 | _GEN_19989; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20230 = _GEN_36428 | _GEN_19990; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20231 = _GEN_36429 | _GEN_19991; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20232 = _GEN_36430 | _GEN_19992; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20233 = _GEN_36431 | _GEN_19993; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20234 = _GEN_36432 | _GEN_19994; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20235 = _GEN_36433 | _GEN_19995; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20236 = _T_446 ? _GEN_20228 : _GEN_19988; // @[sequencer-master.scala 154:24]
  wire  _GEN_20237 = _T_446 ? _GEN_20229 : _GEN_19989; // @[sequencer-master.scala 154:24]
  wire  _GEN_20238 = _T_446 ? _GEN_20230 : _GEN_19990; // @[sequencer-master.scala 154:24]
  wire  _GEN_20239 = _T_446 ? _GEN_20231 : _GEN_19991; // @[sequencer-master.scala 154:24]
  wire  _GEN_20240 = _T_446 ? _GEN_20232 : _GEN_19992; // @[sequencer-master.scala 154:24]
  wire  _GEN_20241 = _T_446 ? _GEN_20233 : _GEN_19993; // @[sequencer-master.scala 154:24]
  wire  _GEN_20242 = _T_446 ? _GEN_20234 : _GEN_19994; // @[sequencer-master.scala 154:24]
  wire  _GEN_20243 = _T_446 ? _GEN_20235 : _GEN_19995; // @[sequencer-master.scala 154:24]
  wire  _GEN_20244 = _GEN_36426 | _GEN_20004; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20245 = _GEN_36427 | _GEN_20005; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20246 = _GEN_36428 | _GEN_20006; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20247 = _GEN_36429 | _GEN_20007; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20248 = _GEN_36430 | _GEN_20008; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20249 = _GEN_36431 | _GEN_20009; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20250 = _GEN_36432 | _GEN_20010; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20251 = _GEN_36433 | _GEN_20011; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20252 = _T_468 ? _GEN_20244 : _GEN_20004; // @[sequencer-master.scala 154:24]
  wire  _GEN_20253 = _T_468 ? _GEN_20245 : _GEN_20005; // @[sequencer-master.scala 154:24]
  wire  _GEN_20254 = _T_468 ? _GEN_20246 : _GEN_20006; // @[sequencer-master.scala 154:24]
  wire  _GEN_20255 = _T_468 ? _GEN_20247 : _GEN_20007; // @[sequencer-master.scala 154:24]
  wire  _GEN_20256 = _T_468 ? _GEN_20248 : _GEN_20008; // @[sequencer-master.scala 154:24]
  wire  _GEN_20257 = _T_468 ? _GEN_20249 : _GEN_20009; // @[sequencer-master.scala 154:24]
  wire  _GEN_20258 = _T_468 ? _GEN_20250 : _GEN_20010; // @[sequencer-master.scala 154:24]
  wire  _GEN_20259 = _T_468 ? _GEN_20251 : _GEN_20011; // @[sequencer-master.scala 154:24]
  wire  _GEN_20260 = _GEN_36426 | _GEN_20020; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20261 = _GEN_36427 | _GEN_20021; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20262 = _GEN_36428 | _GEN_20022; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20263 = _GEN_36429 | _GEN_20023; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20264 = _GEN_36430 | _GEN_20024; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20265 = _GEN_36431 | _GEN_20025; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20266 = _GEN_36432 | _GEN_20026; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20267 = _GEN_36433 | _GEN_20027; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20268 = _T_490 ? _GEN_20260 : _GEN_20020; // @[sequencer-master.scala 154:24]
  wire  _GEN_20269 = _T_490 ? _GEN_20261 : _GEN_20021; // @[sequencer-master.scala 154:24]
  wire  _GEN_20270 = _T_490 ? _GEN_20262 : _GEN_20022; // @[sequencer-master.scala 154:24]
  wire  _GEN_20271 = _T_490 ? _GEN_20263 : _GEN_20023; // @[sequencer-master.scala 154:24]
  wire  _GEN_20272 = _T_490 ? _GEN_20264 : _GEN_20024; // @[sequencer-master.scala 154:24]
  wire  _GEN_20273 = _T_490 ? _GEN_20265 : _GEN_20025; // @[sequencer-master.scala 154:24]
  wire  _GEN_20274 = _T_490 ? _GEN_20266 : _GEN_20026; // @[sequencer-master.scala 154:24]
  wire  _GEN_20275 = _T_490 ? _GEN_20267 : _GEN_20027; // @[sequencer-master.scala 154:24]
  wire  _GEN_20276 = _GEN_36426 | _GEN_20036; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20277 = _GEN_36427 | _GEN_20037; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20278 = _GEN_36428 | _GEN_20038; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20279 = _GEN_36429 | _GEN_20039; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20280 = _GEN_36430 | _GEN_20040; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20281 = _GEN_36431 | _GEN_20041; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20282 = _GEN_36432 | _GEN_20042; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20283 = _GEN_36433 | _GEN_20043; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20284 = _T_512 ? _GEN_20276 : _GEN_20036; // @[sequencer-master.scala 154:24]
  wire  _GEN_20285 = _T_512 ? _GEN_20277 : _GEN_20037; // @[sequencer-master.scala 154:24]
  wire  _GEN_20286 = _T_512 ? _GEN_20278 : _GEN_20038; // @[sequencer-master.scala 154:24]
  wire  _GEN_20287 = _T_512 ? _GEN_20279 : _GEN_20039; // @[sequencer-master.scala 154:24]
  wire  _GEN_20288 = _T_512 ? _GEN_20280 : _GEN_20040; // @[sequencer-master.scala 154:24]
  wire  _GEN_20289 = _T_512 ? _GEN_20281 : _GEN_20041; // @[sequencer-master.scala 154:24]
  wire  _GEN_20290 = _T_512 ? _GEN_20282 : _GEN_20042; // @[sequencer-master.scala 154:24]
  wire  _GEN_20291 = _T_512 ? _GEN_20283 : _GEN_20043; // @[sequencer-master.scala 154:24]
  wire  _GEN_20292 = _GEN_36426 | _GEN_20052; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20293 = _GEN_36427 | _GEN_20053; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20294 = _GEN_36428 | _GEN_20054; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20295 = _GEN_36429 | _GEN_20055; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20296 = _GEN_36430 | _GEN_20056; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20297 = _GEN_36431 | _GEN_20057; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20298 = _GEN_36432 | _GEN_20058; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20299 = _GEN_36433 | _GEN_20059; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20300 = _T_534 ? _GEN_20292 : _GEN_20052; // @[sequencer-master.scala 154:24]
  wire  _GEN_20301 = _T_534 ? _GEN_20293 : _GEN_20053; // @[sequencer-master.scala 154:24]
  wire  _GEN_20302 = _T_534 ? _GEN_20294 : _GEN_20054; // @[sequencer-master.scala 154:24]
  wire  _GEN_20303 = _T_534 ? _GEN_20295 : _GEN_20055; // @[sequencer-master.scala 154:24]
  wire  _GEN_20304 = _T_534 ? _GEN_20296 : _GEN_20056; // @[sequencer-master.scala 154:24]
  wire  _GEN_20305 = _T_534 ? _GEN_20297 : _GEN_20057; // @[sequencer-master.scala 154:24]
  wire  _GEN_20306 = _T_534 ? _GEN_20298 : _GEN_20058; // @[sequencer-master.scala 154:24]
  wire  _GEN_20307 = _T_534 ? _GEN_20299 : _GEN_20059; // @[sequencer-master.scala 154:24]
  wire [1:0] _e_T_1647_rports = {{1'd0}, _T_1631}; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20308 = 3'h0 == _T_1647 ? _e_T_1647_rports : _GEN_19284; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20309 = 3'h1 == _T_1647 ? _e_T_1647_rports : _GEN_19285; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20310 = 3'h2 == _T_1647 ? _e_T_1647_rports : _GEN_19286; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20311 = 3'h3 == _T_1647 ? _e_T_1647_rports : _GEN_19287; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20312 = 3'h4 == _T_1647 ? _e_T_1647_rports : _GEN_19288; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20313 = 3'h5 == _T_1647 ? _e_T_1647_rports : _GEN_19289; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20314 = 3'h6 == _T_1647 ? _e_T_1647_rports : _GEN_19290; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_20315 = 3'h7 == _T_1647 ? _e_T_1647_rports : _GEN_19291; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_20316 = 3'h0 == _T_1647 ? 4'h0 : _GEN_19292; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20317 = 3'h1 == _T_1647 ? 4'h0 : _GEN_19293; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20318 = 3'h2 == _T_1647 ? 4'h0 : _GEN_19294; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20319 = 3'h3 == _T_1647 ? 4'h0 : _GEN_19295; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20320 = 3'h4 == _T_1647 ? 4'h0 : _GEN_19296; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20321 = 3'h5 == _T_1647 ? 4'h0 : _GEN_19297; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20322 = 3'h6 == _T_1647 ? 4'h0 : _GEN_19298; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_20323 = 3'h7 == _T_1647 ? 4'h0 : _GEN_19299; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_20324 = 3'h0 == _T_1647 ? 3'h0 : _GEN_19300; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20325 = 3'h1 == _T_1647 ? 3'h0 : _GEN_19301; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20326 = 3'h2 == _T_1647 ? 3'h0 : _GEN_19302; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20327 = 3'h3 == _T_1647 ? 3'h0 : _GEN_19303; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20328 = 3'h4 == _T_1647 ? 3'h0 : _GEN_19304; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20329 = 3'h5 == _T_1647 ? 3'h0 : _GEN_19305; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20330 = 3'h6 == _T_1647 ? 3'h0 : _GEN_19306; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_20331 = 3'h7 == _T_1647 ? 3'h0 : _GEN_19307; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_20332 = _GEN_36426 & _GEN_34121 | _GEN_20188; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20333 = _GEN_36426 & _GEN_34122 | _GEN_20204; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20334 = _GEN_36426 & _GEN_34123 | _GEN_20220; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20335 = _GEN_36426 & _GEN_34124 | _GEN_20236; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20336 = _GEN_36426 & _GEN_34125 | _GEN_20252; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20337 = _GEN_36426 & _GEN_34126 | _GEN_20268; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20338 = _GEN_36426 & _GEN_34127 | _GEN_20284; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20339 = _GEN_36426 & _GEN_34128 | _GEN_20300; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20340 = _GEN_36427 & _GEN_34121 | _GEN_20189; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20341 = _GEN_36427 & _GEN_34122 | _GEN_20205; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20342 = _GEN_36427 & _GEN_34123 | _GEN_20221; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20343 = _GEN_36427 & _GEN_34124 | _GEN_20237; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20344 = _GEN_36427 & _GEN_34125 | _GEN_20253; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20345 = _GEN_36427 & _GEN_34126 | _GEN_20269; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20346 = _GEN_36427 & _GEN_34127 | _GEN_20285; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20347 = _GEN_36427 & _GEN_34128 | _GEN_20301; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20348 = _GEN_36428 & _GEN_34121 | _GEN_20190; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20349 = _GEN_36428 & _GEN_34122 | _GEN_20206; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20350 = _GEN_36428 & _GEN_34123 | _GEN_20222; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20351 = _GEN_36428 & _GEN_34124 | _GEN_20238; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20352 = _GEN_36428 & _GEN_34125 | _GEN_20254; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20353 = _GEN_36428 & _GEN_34126 | _GEN_20270; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20354 = _GEN_36428 & _GEN_34127 | _GEN_20286; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20355 = _GEN_36428 & _GEN_34128 | _GEN_20302; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20356 = _GEN_36429 & _GEN_34121 | _GEN_20191; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20357 = _GEN_36429 & _GEN_34122 | _GEN_20207; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20358 = _GEN_36429 & _GEN_34123 | _GEN_20223; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20359 = _GEN_36429 & _GEN_34124 | _GEN_20239; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20360 = _GEN_36429 & _GEN_34125 | _GEN_20255; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20361 = _GEN_36429 & _GEN_34126 | _GEN_20271; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20362 = _GEN_36429 & _GEN_34127 | _GEN_20287; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20363 = _GEN_36429 & _GEN_34128 | _GEN_20303; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20364 = _GEN_36430 & _GEN_34121 | _GEN_20192; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20365 = _GEN_36430 & _GEN_34122 | _GEN_20208; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20366 = _GEN_36430 & _GEN_34123 | _GEN_20224; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20367 = _GEN_36430 & _GEN_34124 | _GEN_20240; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20368 = _GEN_36430 & _GEN_34125 | _GEN_20256; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20369 = _GEN_36430 & _GEN_34126 | _GEN_20272; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20370 = _GEN_36430 & _GEN_34127 | _GEN_20288; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20371 = _GEN_36430 & _GEN_34128 | _GEN_20304; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20372 = _GEN_36431 & _GEN_34121 | _GEN_20193; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20373 = _GEN_36431 & _GEN_34122 | _GEN_20209; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20374 = _GEN_36431 & _GEN_34123 | _GEN_20225; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20375 = _GEN_36431 & _GEN_34124 | _GEN_20241; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20376 = _GEN_36431 & _GEN_34125 | _GEN_20257; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20377 = _GEN_36431 & _GEN_34126 | _GEN_20273; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20378 = _GEN_36431 & _GEN_34127 | _GEN_20289; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20379 = _GEN_36431 & _GEN_34128 | _GEN_20305; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20380 = _GEN_36432 & _GEN_34121 | _GEN_20194; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20381 = _GEN_36432 & _GEN_34122 | _GEN_20210; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20382 = _GEN_36432 & _GEN_34123 | _GEN_20226; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20383 = _GEN_36432 & _GEN_34124 | _GEN_20242; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20384 = _GEN_36432 & _GEN_34125 | _GEN_20258; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20385 = _GEN_36432 & _GEN_34126 | _GEN_20274; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20386 = _GEN_36432 & _GEN_34127 | _GEN_20290; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20387 = _GEN_36432 & _GEN_34128 | _GEN_20306; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20388 = _GEN_36433 & _GEN_34121 | _GEN_20195; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20389 = _GEN_36433 & _GEN_34122 | _GEN_20211; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20390 = _GEN_36433 & _GEN_34123 | _GEN_20227; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20391 = _GEN_36433 & _GEN_34124 | _GEN_20243; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20392 = _GEN_36433 & _GEN_34125 | _GEN_20259; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20393 = _GEN_36433 & _GEN_34126 | _GEN_20275; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20394 = _GEN_36433 & _GEN_34127 | _GEN_20291; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_20395 = _GEN_36433 & _GEN_34128 | _GEN_20307; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_36778 = 3'h0 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20396 = 3'h0 == _T_1649 | (3'h0 == _T_1647 | (3'h0 == _T_1645 | (_GEN_32729 | _GEN_17834))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36779 = 3'h1 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20397 = 3'h1 == _T_1649 | (3'h1 == _T_1647 | (3'h1 == _T_1645 | (_GEN_32730 | _GEN_17835))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36780 = 3'h2 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20398 = 3'h2 == _T_1649 | (3'h2 == _T_1647 | (3'h2 == _T_1645 | (_GEN_32731 | _GEN_17836))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36781 = 3'h3 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20399 = 3'h3 == _T_1649 | (3'h3 == _T_1647 | (3'h3 == _T_1645 | (_GEN_32732 | _GEN_17837))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36782 = 3'h4 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20400 = 3'h4 == _T_1649 | (3'h4 == _T_1647 | (3'h4 == _T_1645 | (_GEN_32733 | _GEN_17838))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36783 = 3'h5 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20401 = 3'h5 == _T_1649 | (3'h5 == _T_1647 | (3'h5 == _T_1645 | (_GEN_32734 | _GEN_17839))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36784 = 3'h6 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20402 = 3'h6 == _T_1649 | (3'h6 == _T_1647 | (3'h6 == _T_1645 | (_GEN_32735 | _GEN_17840))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_36785 = 3'h7 == _T_1649; // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20403 = 3'h7 == _T_1649 | (3'h7 == _T_1647 | (3'h7 == _T_1645 | (_GEN_32736 | _GEN_17841))); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_20412 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19900; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20413 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19901; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20414 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19902; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20415 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19903; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20416 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19904; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20417 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19905; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20418 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19906; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20419 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19907; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_20420 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20132; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20421 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20133; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20422 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20134; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20423 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20135; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20424 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20136; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20425 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20137; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20426 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20138; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20427 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20139; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_20428 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19596; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20429 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19597; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20430 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19598; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20431 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19599; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20432 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19600; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20433 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19601; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20434 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19602; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20435 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19603; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_20436 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19604; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20437 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19605; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20438 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19606; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20439 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19607; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20440 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19608; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20441 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19609; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20442 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19610; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20443 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19611; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_20444 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19612; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20445 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19613; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20446 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19614; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20447 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19615; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20448 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19616; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20449 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19617; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20450 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19618; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20451 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19619; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_20452 = _GEN_36778 | (_GEN_36426 | (_GEN_34121 | (_GEN_32729 | _GEN_17890))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20453 = _GEN_36779 | (_GEN_36427 | (_GEN_34122 | (_GEN_32730 | _GEN_17891))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20454 = _GEN_36780 | (_GEN_36428 | (_GEN_34123 | (_GEN_32731 | _GEN_17892))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20455 = _GEN_36781 | (_GEN_36429 | (_GEN_34124 | (_GEN_32732 | _GEN_17893))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20456 = _GEN_36782 | (_GEN_36430 | (_GEN_34125 | (_GEN_32733 | _GEN_17894))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20457 = _GEN_36783 | (_GEN_36431 | (_GEN_34126 | (_GEN_32734 | _GEN_17895))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20458 = _GEN_36784 | (_GEN_36432 | (_GEN_34127 | (_GEN_32735 | _GEN_17896))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20459 = _GEN_36785 | (_GEN_36433 | (_GEN_34128 | (_GEN_32736 | _GEN_17897))); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_20460 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20332; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20461 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20340; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20462 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20348; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20463 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20356; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20464 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20364; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20465 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20372; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20466 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20380; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20467 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20388; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20468 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19636; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20469 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19637; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20470 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19638; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20471 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19639; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20472 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19640; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20473 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19641; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20474 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19642; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20475 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19643; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20476 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19644; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20477 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19645; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20478 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19646; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20479 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19647; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20480 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19648; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20481 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19649; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20482 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19650; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20483 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19651; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20484 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20333; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20485 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20341; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20486 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20349; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20487 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20357; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20488 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20365; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20489 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20373; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20490 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20381; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20491 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20389; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20492 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19660; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20493 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19661; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20494 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19662; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20495 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19663; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20496 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19664; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20497 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19665; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20498 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19666; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20499 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19667; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20500 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19668; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20501 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19669; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20502 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19670; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20503 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19671; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20504 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19672; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20505 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19673; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20506 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19674; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20507 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19675; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20508 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20334; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20509 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20342; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20510 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20350; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20511 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20358; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20512 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20366; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20513 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20374; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20514 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20382; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20515 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20390; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20516 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19684; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20517 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19685; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20518 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19686; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20519 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19687; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20520 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19688; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20521 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19689; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20522 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19690; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20523 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19691; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20524 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19692; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20525 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19693; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20526 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19694; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20527 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19695; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20528 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19696; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20529 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19697; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20530 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19698; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20531 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19699; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20532 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20335; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20533 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20343; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20534 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20351; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20535 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20359; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20536 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20367; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20537 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20375; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20538 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20383; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20539 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20391; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20540 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19708; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20541 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19709; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20542 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19710; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20543 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19711; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20544 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19712; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20545 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19713; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20546 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19714; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20547 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19715; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20548 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19716; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20549 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19717; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20550 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19718; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20551 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19719; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20552 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19720; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20553 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19721; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20554 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19722; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20555 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19723; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20556 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20336; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20557 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20344; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20558 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20352; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20559 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20360; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20560 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20368; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20561 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20376; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20562 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20384; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20563 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20392; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20564 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19732; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20565 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19733; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20566 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19734; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20567 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19735; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20568 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19736; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20569 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19737; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20570 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19738; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20571 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19739; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20572 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19740; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20573 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19741; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20574 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19742; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20575 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19743; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20576 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19744; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20577 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19745; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20578 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19746; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20579 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19747; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20580 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20337; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20581 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20345; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20582 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20353; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20583 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20361; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20584 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20369; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20585 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20377; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20586 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20385; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20587 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20393; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20588 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19756; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20589 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19757; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20590 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19758; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20591 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19759; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20592 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19760; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20593 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19761; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20594 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19762; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20595 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19763; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20596 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19764; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20597 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19765; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20598 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19766; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20599 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19767; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20600 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19768; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20601 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19769; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20602 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19770; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20603 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19771; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20604 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20338; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20605 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20346; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20606 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20354; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20607 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20362; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20608 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20370; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20609 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20378; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20610 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20386; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20611 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20394; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20612 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19780; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20613 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19781; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20614 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19782; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20615 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19783; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20616 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19784; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20617 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19785; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20618 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19786; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20619 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19787; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20620 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19788; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20621 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19789; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20622 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19790; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20623 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19791; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20624 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19792; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20625 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19793; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20626 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19794; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20627 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19795; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20628 = 3'h0 == _T_1649 ? 1'h0 : _GEN_20339; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20629 = 3'h1 == _T_1649 ? 1'h0 : _GEN_20347; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20630 = 3'h2 == _T_1649 ? 1'h0 : _GEN_20355; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20631 = 3'h3 == _T_1649 ? 1'h0 : _GEN_20363; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20632 = 3'h4 == _T_1649 ? 1'h0 : _GEN_20371; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20633 = 3'h5 == _T_1649 ? 1'h0 : _GEN_20379; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20634 = 3'h6 == _T_1649 ? 1'h0 : _GEN_20387; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20635 = 3'h7 == _T_1649 ? 1'h0 : _GEN_20395; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_20636 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19804; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20637 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19805; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20638 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19806; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20639 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19807; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20640 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19808; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20641 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19809; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20642 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19810; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20643 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19811; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_20644 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19812; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20645 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19813; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20646 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19814; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20647 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19815; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20648 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19816; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20649 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19817; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20650 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19818; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20651 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19819; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_20652 = 3'h0 == _T_1649 ? 1'h0 : _GEN_19820; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20653 = 3'h1 == _T_1649 ? 1'h0 : _GEN_19821; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20654 = 3'h2 == _T_1649 ? 1'h0 : _GEN_19822; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20655 = 3'h3 == _T_1649 ? 1'h0 : _GEN_19823; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20656 = 3'h4 == _T_1649 ? 1'h0 : _GEN_19824; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20657 = 3'h5 == _T_1649 ? 1'h0 : _GEN_19825; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20658 = 3'h6 == _T_1649 ? 1'h0 : _GEN_19826; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20659 = 3'h7 == _T_1649 ? 1'h0 : _GEN_19827; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_20668 = _GEN_36778 | e_0_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20669 = _GEN_36779 | e_1_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20670 = _GEN_36780 | e_2_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20671 = _GEN_36781 | e_3_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20672 = _GEN_36782 | e_4_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20673 = _GEN_36783 | e_5_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20674 = _GEN_36784 | e_6_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_20675 = _GEN_36785 | e_7_active_vlu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_20676 = 3'h0 == _T_1649 ? io_op_bits_fn_union : _GEN_19844; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20677 = 3'h1 == _T_1649 ? io_op_bits_fn_union : _GEN_19845; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20678 = 3'h2 == _T_1649 ? io_op_bits_fn_union : _GEN_19846; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20679 = 3'h3 == _T_1649 ? io_op_bits_fn_union : _GEN_19847; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20680 = 3'h4 == _T_1649 ? io_op_bits_fn_union : _GEN_19848; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20681 = 3'h5 == _T_1649 ? io_op_bits_fn_union : _GEN_19849; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20682 = 3'h6 == _T_1649 ? io_op_bits_fn_union : _GEN_19850; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_20683 = 3'h7 == _T_1649 ? io_op_bits_fn_union : _GEN_19851; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [7:0] _GEN_20684 = 3'h0 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16134; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20685 = 3'h1 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16135; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20686 = 3'h2 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16136; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20687 = 3'h3 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16137; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20688 = 3'h4 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16138; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20689 = 3'h5 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16139; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20690 = 3'h6 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16140; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20691 = 3'h7 == _T_1649 ? io_op_bits_base_vd_id : _GEN_16141; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20692 = 3'h0 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20444; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20693 = 3'h1 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20445; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20694 = 3'h2 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20446; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20695 = 3'h3 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20447; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20696 = 3'h4 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20448; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20697 = 3'h5 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20449; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20698 = 3'h6 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20450; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20699 = 3'h7 == _T_1649 ? io_op_bits_base_vd_valid : _GEN_20451; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20700 = 3'h0 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16142; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20701 = 3'h1 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16143; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20702 = 3'h2 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16144; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20703 = 3'h3 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16145; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20704 = 3'h4 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16146; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20705 = 3'h5 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16147; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20706 = 3'h6 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16148; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20707 = 3'h7 == _T_1649 ? io_op_bits_base_vd_scalar : _GEN_16149; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20708 = 3'h0 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16150; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20709 = 3'h1 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16151; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20710 = 3'h2 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16152; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20711 = 3'h3 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16153; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20712 = 3'h4 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16154; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20713 = 3'h5 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16155; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20714 = 3'h6 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16156; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_20715 = 3'h7 == _T_1649 ? io_op_bits_base_vd_pred : _GEN_16157; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20716 = 3'h0 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16158; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20717 = 3'h1 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16159; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20718 = 3'h2 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16160; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20719 = 3'h3 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16161; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20720 = 3'h4 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16162; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20721 = 3'h5 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16163; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20722 = 3'h6 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16164; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_20723 = 3'h7 == _T_1649 ? io_op_bits_base_vd_prec : _GEN_16165; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_20724 = 3'h0 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16166; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20725 = 3'h1 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16167; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20726 = 3'h2 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16168; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20727 = 3'h3 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16169; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20728 = 3'h4 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16170; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20729 = 3'h5 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16171; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20730 = 3'h6 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16172; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20731 = 3'h7 == _T_1649 ? io_op_bits_reg_vd_id : _GEN_16173; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_20732 = io_op_bits_base_vd_valid ? _GEN_20684 : _GEN_16134; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20733 = io_op_bits_base_vd_valid ? _GEN_20685 : _GEN_16135; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20734 = io_op_bits_base_vd_valid ? _GEN_20686 : _GEN_16136; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20735 = io_op_bits_base_vd_valid ? _GEN_20687 : _GEN_16137; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20736 = io_op_bits_base_vd_valid ? _GEN_20688 : _GEN_16138; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20737 = io_op_bits_base_vd_valid ? _GEN_20689 : _GEN_16139; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20738 = io_op_bits_base_vd_valid ? _GEN_20690 : _GEN_16140; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20739 = io_op_bits_base_vd_valid ? _GEN_20691 : _GEN_16141; // @[sequencer-master.scala 362:41]
  wire  _GEN_20740 = io_op_bits_base_vd_valid ? _GEN_20692 : _GEN_20444; // @[sequencer-master.scala 362:41]
  wire  _GEN_20741 = io_op_bits_base_vd_valid ? _GEN_20693 : _GEN_20445; // @[sequencer-master.scala 362:41]
  wire  _GEN_20742 = io_op_bits_base_vd_valid ? _GEN_20694 : _GEN_20446; // @[sequencer-master.scala 362:41]
  wire  _GEN_20743 = io_op_bits_base_vd_valid ? _GEN_20695 : _GEN_20447; // @[sequencer-master.scala 362:41]
  wire  _GEN_20744 = io_op_bits_base_vd_valid ? _GEN_20696 : _GEN_20448; // @[sequencer-master.scala 362:41]
  wire  _GEN_20745 = io_op_bits_base_vd_valid ? _GEN_20697 : _GEN_20449; // @[sequencer-master.scala 362:41]
  wire  _GEN_20746 = io_op_bits_base_vd_valid ? _GEN_20698 : _GEN_20450; // @[sequencer-master.scala 362:41]
  wire  _GEN_20747 = io_op_bits_base_vd_valid ? _GEN_20699 : _GEN_20451; // @[sequencer-master.scala 362:41]
  wire  _GEN_20748 = io_op_bits_base_vd_valid ? _GEN_20700 : _GEN_16142; // @[sequencer-master.scala 362:41]
  wire  _GEN_20749 = io_op_bits_base_vd_valid ? _GEN_20701 : _GEN_16143; // @[sequencer-master.scala 362:41]
  wire  _GEN_20750 = io_op_bits_base_vd_valid ? _GEN_20702 : _GEN_16144; // @[sequencer-master.scala 362:41]
  wire  _GEN_20751 = io_op_bits_base_vd_valid ? _GEN_20703 : _GEN_16145; // @[sequencer-master.scala 362:41]
  wire  _GEN_20752 = io_op_bits_base_vd_valid ? _GEN_20704 : _GEN_16146; // @[sequencer-master.scala 362:41]
  wire  _GEN_20753 = io_op_bits_base_vd_valid ? _GEN_20705 : _GEN_16147; // @[sequencer-master.scala 362:41]
  wire  _GEN_20754 = io_op_bits_base_vd_valid ? _GEN_20706 : _GEN_16148; // @[sequencer-master.scala 362:41]
  wire  _GEN_20755 = io_op_bits_base_vd_valid ? _GEN_20707 : _GEN_16149; // @[sequencer-master.scala 362:41]
  wire  _GEN_20756 = io_op_bits_base_vd_valid ? _GEN_20708 : _GEN_16150; // @[sequencer-master.scala 362:41]
  wire  _GEN_20757 = io_op_bits_base_vd_valid ? _GEN_20709 : _GEN_16151; // @[sequencer-master.scala 362:41]
  wire  _GEN_20758 = io_op_bits_base_vd_valid ? _GEN_20710 : _GEN_16152; // @[sequencer-master.scala 362:41]
  wire  _GEN_20759 = io_op_bits_base_vd_valid ? _GEN_20711 : _GEN_16153; // @[sequencer-master.scala 362:41]
  wire  _GEN_20760 = io_op_bits_base_vd_valid ? _GEN_20712 : _GEN_16154; // @[sequencer-master.scala 362:41]
  wire  _GEN_20761 = io_op_bits_base_vd_valid ? _GEN_20713 : _GEN_16155; // @[sequencer-master.scala 362:41]
  wire  _GEN_20762 = io_op_bits_base_vd_valid ? _GEN_20714 : _GEN_16156; // @[sequencer-master.scala 362:41]
  wire  _GEN_20763 = io_op_bits_base_vd_valid ? _GEN_20715 : _GEN_16157; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20764 = io_op_bits_base_vd_valid ? _GEN_20716 : _GEN_16158; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20765 = io_op_bits_base_vd_valid ? _GEN_20717 : _GEN_16159; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20766 = io_op_bits_base_vd_valid ? _GEN_20718 : _GEN_16160; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20767 = io_op_bits_base_vd_valid ? _GEN_20719 : _GEN_16161; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20768 = io_op_bits_base_vd_valid ? _GEN_20720 : _GEN_16162; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20769 = io_op_bits_base_vd_valid ? _GEN_20721 : _GEN_16163; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20770 = io_op_bits_base_vd_valid ? _GEN_20722 : _GEN_16164; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_20771 = io_op_bits_base_vd_valid ? _GEN_20723 : _GEN_16165; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20772 = io_op_bits_base_vd_valid ? _GEN_20724 : _GEN_16166; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20773 = io_op_bits_base_vd_valid ? _GEN_20725 : _GEN_16167; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20774 = io_op_bits_base_vd_valid ? _GEN_20726 : _GEN_16168; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20775 = io_op_bits_base_vd_valid ? _GEN_20727 : _GEN_16169; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20776 = io_op_bits_base_vd_valid ? _GEN_20728 : _GEN_16170; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20777 = io_op_bits_base_vd_valid ? _GEN_20729 : _GEN_16171; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20778 = io_op_bits_base_vd_valid ? _GEN_20730 : _GEN_16172; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_20779 = io_op_bits_base_vd_valid ? _GEN_20731 : _GEN_16173; // @[sequencer-master.scala 362:41]
  wire  _GEN_20780 = _GEN_36778 | _GEN_20468; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20781 = _GEN_36779 | _GEN_20469; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20782 = _GEN_36780 | _GEN_20470; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20783 = _GEN_36781 | _GEN_20471; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20784 = _GEN_36782 | _GEN_20472; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20785 = _GEN_36783 | _GEN_20473; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20786 = _GEN_36784 | _GEN_20474; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20787 = _GEN_36785 | _GEN_20475; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20788 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20780 : _GEN_20468; // @[sequencer-master.scala 161:86]
  wire  _GEN_20789 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20781 : _GEN_20469; // @[sequencer-master.scala 161:86]
  wire  _GEN_20790 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20782 : _GEN_20470; // @[sequencer-master.scala 161:86]
  wire  _GEN_20791 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20783 : _GEN_20471; // @[sequencer-master.scala 161:86]
  wire  _GEN_20792 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20784 : _GEN_20472; // @[sequencer-master.scala 161:86]
  wire  _GEN_20793 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20785 : _GEN_20473; // @[sequencer-master.scala 161:86]
  wire  _GEN_20794 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20786 : _GEN_20474; // @[sequencer-master.scala 161:86]
  wire  _GEN_20795 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_20787 : _GEN_20475; // @[sequencer-master.scala 161:86]
  wire  _GEN_20796 = _GEN_36778 | _GEN_20492; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20797 = _GEN_36779 | _GEN_20493; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20798 = _GEN_36780 | _GEN_20494; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20799 = _GEN_36781 | _GEN_20495; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20800 = _GEN_36782 | _GEN_20496; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20801 = _GEN_36783 | _GEN_20497; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20802 = _GEN_36784 | _GEN_20498; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20803 = _GEN_36785 | _GEN_20499; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20804 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20796 : _GEN_20492; // @[sequencer-master.scala 161:86]
  wire  _GEN_20805 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20797 : _GEN_20493; // @[sequencer-master.scala 161:86]
  wire  _GEN_20806 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20798 : _GEN_20494; // @[sequencer-master.scala 161:86]
  wire  _GEN_20807 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20799 : _GEN_20495; // @[sequencer-master.scala 161:86]
  wire  _GEN_20808 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20800 : _GEN_20496; // @[sequencer-master.scala 161:86]
  wire  _GEN_20809 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20801 : _GEN_20497; // @[sequencer-master.scala 161:86]
  wire  _GEN_20810 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20802 : _GEN_20498; // @[sequencer-master.scala 161:86]
  wire  _GEN_20811 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_20803 : _GEN_20499; // @[sequencer-master.scala 161:86]
  wire  _GEN_20812 = _GEN_36778 | _GEN_20516; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20813 = _GEN_36779 | _GEN_20517; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20814 = _GEN_36780 | _GEN_20518; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20815 = _GEN_36781 | _GEN_20519; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20816 = _GEN_36782 | _GEN_20520; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20817 = _GEN_36783 | _GEN_20521; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20818 = _GEN_36784 | _GEN_20522; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20819 = _GEN_36785 | _GEN_20523; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20820 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20812 : _GEN_20516; // @[sequencer-master.scala 161:86]
  wire  _GEN_20821 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20813 : _GEN_20517; // @[sequencer-master.scala 161:86]
  wire  _GEN_20822 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20814 : _GEN_20518; // @[sequencer-master.scala 161:86]
  wire  _GEN_20823 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20815 : _GEN_20519; // @[sequencer-master.scala 161:86]
  wire  _GEN_20824 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20816 : _GEN_20520; // @[sequencer-master.scala 161:86]
  wire  _GEN_20825 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20817 : _GEN_20521; // @[sequencer-master.scala 161:86]
  wire  _GEN_20826 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20818 : _GEN_20522; // @[sequencer-master.scala 161:86]
  wire  _GEN_20827 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_20819 : _GEN_20523; // @[sequencer-master.scala 161:86]
  wire  _GEN_20828 = _GEN_36778 | _GEN_20540; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20829 = _GEN_36779 | _GEN_20541; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20830 = _GEN_36780 | _GEN_20542; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20831 = _GEN_36781 | _GEN_20543; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20832 = _GEN_36782 | _GEN_20544; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20833 = _GEN_36783 | _GEN_20545; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20834 = _GEN_36784 | _GEN_20546; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20835 = _GEN_36785 | _GEN_20547; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20836 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20828 : _GEN_20540; // @[sequencer-master.scala 161:86]
  wire  _GEN_20837 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20829 : _GEN_20541; // @[sequencer-master.scala 161:86]
  wire  _GEN_20838 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20830 : _GEN_20542; // @[sequencer-master.scala 161:86]
  wire  _GEN_20839 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20831 : _GEN_20543; // @[sequencer-master.scala 161:86]
  wire  _GEN_20840 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20832 : _GEN_20544; // @[sequencer-master.scala 161:86]
  wire  _GEN_20841 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20833 : _GEN_20545; // @[sequencer-master.scala 161:86]
  wire  _GEN_20842 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20834 : _GEN_20546; // @[sequencer-master.scala 161:86]
  wire  _GEN_20843 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_20835 : _GEN_20547; // @[sequencer-master.scala 161:86]
  wire  _GEN_20844 = _GEN_36778 | _GEN_20564; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20845 = _GEN_36779 | _GEN_20565; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20846 = _GEN_36780 | _GEN_20566; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20847 = _GEN_36781 | _GEN_20567; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20848 = _GEN_36782 | _GEN_20568; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20849 = _GEN_36783 | _GEN_20569; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20850 = _GEN_36784 | _GEN_20570; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20851 = _GEN_36785 | _GEN_20571; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20852 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20844 : _GEN_20564; // @[sequencer-master.scala 161:86]
  wire  _GEN_20853 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20845 : _GEN_20565; // @[sequencer-master.scala 161:86]
  wire  _GEN_20854 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20846 : _GEN_20566; // @[sequencer-master.scala 161:86]
  wire  _GEN_20855 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20847 : _GEN_20567; // @[sequencer-master.scala 161:86]
  wire  _GEN_20856 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20848 : _GEN_20568; // @[sequencer-master.scala 161:86]
  wire  _GEN_20857 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20849 : _GEN_20569; // @[sequencer-master.scala 161:86]
  wire  _GEN_20858 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20850 : _GEN_20570; // @[sequencer-master.scala 161:86]
  wire  _GEN_20859 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_20851 : _GEN_20571; // @[sequencer-master.scala 161:86]
  wire  _GEN_20860 = _GEN_36778 | _GEN_20588; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20861 = _GEN_36779 | _GEN_20589; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20862 = _GEN_36780 | _GEN_20590; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20863 = _GEN_36781 | _GEN_20591; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20864 = _GEN_36782 | _GEN_20592; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20865 = _GEN_36783 | _GEN_20593; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20866 = _GEN_36784 | _GEN_20594; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20867 = _GEN_36785 | _GEN_20595; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20868 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20860 : _GEN_20588; // @[sequencer-master.scala 161:86]
  wire  _GEN_20869 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20861 : _GEN_20589; // @[sequencer-master.scala 161:86]
  wire  _GEN_20870 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20862 : _GEN_20590; // @[sequencer-master.scala 161:86]
  wire  _GEN_20871 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20863 : _GEN_20591; // @[sequencer-master.scala 161:86]
  wire  _GEN_20872 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20864 : _GEN_20592; // @[sequencer-master.scala 161:86]
  wire  _GEN_20873 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20865 : _GEN_20593; // @[sequencer-master.scala 161:86]
  wire  _GEN_20874 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20866 : _GEN_20594; // @[sequencer-master.scala 161:86]
  wire  _GEN_20875 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_20867 : _GEN_20595; // @[sequencer-master.scala 161:86]
  wire  _GEN_20876 = _GEN_36778 | _GEN_20612; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20877 = _GEN_36779 | _GEN_20613; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20878 = _GEN_36780 | _GEN_20614; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20879 = _GEN_36781 | _GEN_20615; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20880 = _GEN_36782 | _GEN_20616; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20881 = _GEN_36783 | _GEN_20617; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20882 = _GEN_36784 | _GEN_20618; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20883 = _GEN_36785 | _GEN_20619; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20884 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20876 : _GEN_20612; // @[sequencer-master.scala 161:86]
  wire  _GEN_20885 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20877 : _GEN_20613; // @[sequencer-master.scala 161:86]
  wire  _GEN_20886 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20878 : _GEN_20614; // @[sequencer-master.scala 161:86]
  wire  _GEN_20887 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20879 : _GEN_20615; // @[sequencer-master.scala 161:86]
  wire  _GEN_20888 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20880 : _GEN_20616; // @[sequencer-master.scala 161:86]
  wire  _GEN_20889 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20881 : _GEN_20617; // @[sequencer-master.scala 161:86]
  wire  _GEN_20890 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20882 : _GEN_20618; // @[sequencer-master.scala 161:86]
  wire  _GEN_20891 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_20883 : _GEN_20619; // @[sequencer-master.scala 161:86]
  wire  _GEN_20892 = _GEN_36778 | _GEN_20636; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20893 = _GEN_36779 | _GEN_20637; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20894 = _GEN_36780 | _GEN_20638; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20895 = _GEN_36781 | _GEN_20639; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20896 = _GEN_36782 | _GEN_20640; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20897 = _GEN_36783 | _GEN_20641; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20898 = _GEN_36784 | _GEN_20642; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20899 = _GEN_36785 | _GEN_20643; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_20900 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20892 : _GEN_20636; // @[sequencer-master.scala 161:86]
  wire  _GEN_20901 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20893 : _GEN_20637; // @[sequencer-master.scala 161:86]
  wire  _GEN_20902 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20894 : _GEN_20638; // @[sequencer-master.scala 161:86]
  wire  _GEN_20903 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20895 : _GEN_20639; // @[sequencer-master.scala 161:86]
  wire  _GEN_20904 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20896 : _GEN_20640; // @[sequencer-master.scala 161:86]
  wire  _GEN_20905 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20897 : _GEN_20641; // @[sequencer-master.scala 161:86]
  wire  _GEN_20906 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20898 : _GEN_20642; // @[sequencer-master.scala 161:86]
  wire  _GEN_20907 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_20899 : _GEN_20643; // @[sequencer-master.scala 161:86]
  wire  _GEN_20908 = _GEN_36778 | _GEN_20476; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20909 = _GEN_36779 | _GEN_20477; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20910 = _GEN_36780 | _GEN_20478; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20911 = _GEN_36781 | _GEN_20479; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20912 = _GEN_36782 | _GEN_20480; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20913 = _GEN_36783 | _GEN_20481; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20914 = _GEN_36784 | _GEN_20482; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20915 = _GEN_36785 | _GEN_20483; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20916 = _T_1442 ? _GEN_20908 : _GEN_20476; // @[sequencer-master.scala 168:32]
  wire  _GEN_20917 = _T_1442 ? _GEN_20909 : _GEN_20477; // @[sequencer-master.scala 168:32]
  wire  _GEN_20918 = _T_1442 ? _GEN_20910 : _GEN_20478; // @[sequencer-master.scala 168:32]
  wire  _GEN_20919 = _T_1442 ? _GEN_20911 : _GEN_20479; // @[sequencer-master.scala 168:32]
  wire  _GEN_20920 = _T_1442 ? _GEN_20912 : _GEN_20480; // @[sequencer-master.scala 168:32]
  wire  _GEN_20921 = _T_1442 ? _GEN_20913 : _GEN_20481; // @[sequencer-master.scala 168:32]
  wire  _GEN_20922 = _T_1442 ? _GEN_20914 : _GEN_20482; // @[sequencer-master.scala 168:32]
  wire  _GEN_20923 = _T_1442 ? _GEN_20915 : _GEN_20483; // @[sequencer-master.scala 168:32]
  wire  _GEN_20924 = _GEN_36778 | _GEN_20500; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20925 = _GEN_36779 | _GEN_20501; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20926 = _GEN_36780 | _GEN_20502; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20927 = _GEN_36781 | _GEN_20503; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20928 = _GEN_36782 | _GEN_20504; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20929 = _GEN_36783 | _GEN_20505; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20930 = _GEN_36784 | _GEN_20506; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20931 = _GEN_36785 | _GEN_20507; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20932 = _T_1464 ? _GEN_20924 : _GEN_20500; // @[sequencer-master.scala 168:32]
  wire  _GEN_20933 = _T_1464 ? _GEN_20925 : _GEN_20501; // @[sequencer-master.scala 168:32]
  wire  _GEN_20934 = _T_1464 ? _GEN_20926 : _GEN_20502; // @[sequencer-master.scala 168:32]
  wire  _GEN_20935 = _T_1464 ? _GEN_20927 : _GEN_20503; // @[sequencer-master.scala 168:32]
  wire  _GEN_20936 = _T_1464 ? _GEN_20928 : _GEN_20504; // @[sequencer-master.scala 168:32]
  wire  _GEN_20937 = _T_1464 ? _GEN_20929 : _GEN_20505; // @[sequencer-master.scala 168:32]
  wire  _GEN_20938 = _T_1464 ? _GEN_20930 : _GEN_20506; // @[sequencer-master.scala 168:32]
  wire  _GEN_20939 = _T_1464 ? _GEN_20931 : _GEN_20507; // @[sequencer-master.scala 168:32]
  wire  _GEN_20940 = _GEN_36778 | _GEN_20524; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20941 = _GEN_36779 | _GEN_20525; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20942 = _GEN_36780 | _GEN_20526; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20943 = _GEN_36781 | _GEN_20527; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20944 = _GEN_36782 | _GEN_20528; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20945 = _GEN_36783 | _GEN_20529; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20946 = _GEN_36784 | _GEN_20530; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20947 = _GEN_36785 | _GEN_20531; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20948 = _T_1486 ? _GEN_20940 : _GEN_20524; // @[sequencer-master.scala 168:32]
  wire  _GEN_20949 = _T_1486 ? _GEN_20941 : _GEN_20525; // @[sequencer-master.scala 168:32]
  wire  _GEN_20950 = _T_1486 ? _GEN_20942 : _GEN_20526; // @[sequencer-master.scala 168:32]
  wire  _GEN_20951 = _T_1486 ? _GEN_20943 : _GEN_20527; // @[sequencer-master.scala 168:32]
  wire  _GEN_20952 = _T_1486 ? _GEN_20944 : _GEN_20528; // @[sequencer-master.scala 168:32]
  wire  _GEN_20953 = _T_1486 ? _GEN_20945 : _GEN_20529; // @[sequencer-master.scala 168:32]
  wire  _GEN_20954 = _T_1486 ? _GEN_20946 : _GEN_20530; // @[sequencer-master.scala 168:32]
  wire  _GEN_20955 = _T_1486 ? _GEN_20947 : _GEN_20531; // @[sequencer-master.scala 168:32]
  wire  _GEN_20956 = _GEN_36778 | _GEN_20548; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20957 = _GEN_36779 | _GEN_20549; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20958 = _GEN_36780 | _GEN_20550; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20959 = _GEN_36781 | _GEN_20551; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20960 = _GEN_36782 | _GEN_20552; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20961 = _GEN_36783 | _GEN_20553; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20962 = _GEN_36784 | _GEN_20554; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20963 = _GEN_36785 | _GEN_20555; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20964 = _T_1508 ? _GEN_20956 : _GEN_20548; // @[sequencer-master.scala 168:32]
  wire  _GEN_20965 = _T_1508 ? _GEN_20957 : _GEN_20549; // @[sequencer-master.scala 168:32]
  wire  _GEN_20966 = _T_1508 ? _GEN_20958 : _GEN_20550; // @[sequencer-master.scala 168:32]
  wire  _GEN_20967 = _T_1508 ? _GEN_20959 : _GEN_20551; // @[sequencer-master.scala 168:32]
  wire  _GEN_20968 = _T_1508 ? _GEN_20960 : _GEN_20552; // @[sequencer-master.scala 168:32]
  wire  _GEN_20969 = _T_1508 ? _GEN_20961 : _GEN_20553; // @[sequencer-master.scala 168:32]
  wire  _GEN_20970 = _T_1508 ? _GEN_20962 : _GEN_20554; // @[sequencer-master.scala 168:32]
  wire  _GEN_20971 = _T_1508 ? _GEN_20963 : _GEN_20555; // @[sequencer-master.scala 168:32]
  wire  _GEN_20972 = _GEN_36778 | _GEN_20572; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20973 = _GEN_36779 | _GEN_20573; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20974 = _GEN_36780 | _GEN_20574; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20975 = _GEN_36781 | _GEN_20575; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20976 = _GEN_36782 | _GEN_20576; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20977 = _GEN_36783 | _GEN_20577; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20978 = _GEN_36784 | _GEN_20578; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20979 = _GEN_36785 | _GEN_20579; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20980 = _T_1530 ? _GEN_20972 : _GEN_20572; // @[sequencer-master.scala 168:32]
  wire  _GEN_20981 = _T_1530 ? _GEN_20973 : _GEN_20573; // @[sequencer-master.scala 168:32]
  wire  _GEN_20982 = _T_1530 ? _GEN_20974 : _GEN_20574; // @[sequencer-master.scala 168:32]
  wire  _GEN_20983 = _T_1530 ? _GEN_20975 : _GEN_20575; // @[sequencer-master.scala 168:32]
  wire  _GEN_20984 = _T_1530 ? _GEN_20976 : _GEN_20576; // @[sequencer-master.scala 168:32]
  wire  _GEN_20985 = _T_1530 ? _GEN_20977 : _GEN_20577; // @[sequencer-master.scala 168:32]
  wire  _GEN_20986 = _T_1530 ? _GEN_20978 : _GEN_20578; // @[sequencer-master.scala 168:32]
  wire  _GEN_20987 = _T_1530 ? _GEN_20979 : _GEN_20579; // @[sequencer-master.scala 168:32]
  wire  _GEN_20988 = _GEN_36778 | _GEN_20596; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20989 = _GEN_36779 | _GEN_20597; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20990 = _GEN_36780 | _GEN_20598; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20991 = _GEN_36781 | _GEN_20599; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20992 = _GEN_36782 | _GEN_20600; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20993 = _GEN_36783 | _GEN_20601; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20994 = _GEN_36784 | _GEN_20602; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20995 = _GEN_36785 | _GEN_20603; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_20996 = _T_1552 ? _GEN_20988 : _GEN_20596; // @[sequencer-master.scala 168:32]
  wire  _GEN_20997 = _T_1552 ? _GEN_20989 : _GEN_20597; // @[sequencer-master.scala 168:32]
  wire  _GEN_20998 = _T_1552 ? _GEN_20990 : _GEN_20598; // @[sequencer-master.scala 168:32]
  wire  _GEN_20999 = _T_1552 ? _GEN_20991 : _GEN_20599; // @[sequencer-master.scala 168:32]
  wire  _GEN_21000 = _T_1552 ? _GEN_20992 : _GEN_20600; // @[sequencer-master.scala 168:32]
  wire  _GEN_21001 = _T_1552 ? _GEN_20993 : _GEN_20601; // @[sequencer-master.scala 168:32]
  wire  _GEN_21002 = _T_1552 ? _GEN_20994 : _GEN_20602; // @[sequencer-master.scala 168:32]
  wire  _GEN_21003 = _T_1552 ? _GEN_20995 : _GEN_20603; // @[sequencer-master.scala 168:32]
  wire  _GEN_21004 = _GEN_36778 | _GEN_20620; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21005 = _GEN_36779 | _GEN_20621; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21006 = _GEN_36780 | _GEN_20622; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21007 = _GEN_36781 | _GEN_20623; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21008 = _GEN_36782 | _GEN_20624; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21009 = _GEN_36783 | _GEN_20625; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21010 = _GEN_36784 | _GEN_20626; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21011 = _GEN_36785 | _GEN_20627; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21012 = _T_1574 ? _GEN_21004 : _GEN_20620; // @[sequencer-master.scala 168:32]
  wire  _GEN_21013 = _T_1574 ? _GEN_21005 : _GEN_20621; // @[sequencer-master.scala 168:32]
  wire  _GEN_21014 = _T_1574 ? _GEN_21006 : _GEN_20622; // @[sequencer-master.scala 168:32]
  wire  _GEN_21015 = _T_1574 ? _GEN_21007 : _GEN_20623; // @[sequencer-master.scala 168:32]
  wire  _GEN_21016 = _T_1574 ? _GEN_21008 : _GEN_20624; // @[sequencer-master.scala 168:32]
  wire  _GEN_21017 = _T_1574 ? _GEN_21009 : _GEN_20625; // @[sequencer-master.scala 168:32]
  wire  _GEN_21018 = _T_1574 ? _GEN_21010 : _GEN_20626; // @[sequencer-master.scala 168:32]
  wire  _GEN_21019 = _T_1574 ? _GEN_21011 : _GEN_20627; // @[sequencer-master.scala 168:32]
  wire  _GEN_21020 = _GEN_36778 | _GEN_20644; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21021 = _GEN_36779 | _GEN_20645; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21022 = _GEN_36780 | _GEN_20646; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21023 = _GEN_36781 | _GEN_20647; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21024 = _GEN_36782 | _GEN_20648; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21025 = _GEN_36783 | _GEN_20649; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21026 = _GEN_36784 | _GEN_20650; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21027 = _GEN_36785 | _GEN_20651; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_21028 = _T_1596 ? _GEN_21020 : _GEN_20644; // @[sequencer-master.scala 168:32]
  wire  _GEN_21029 = _T_1596 ? _GEN_21021 : _GEN_20645; // @[sequencer-master.scala 168:32]
  wire  _GEN_21030 = _T_1596 ? _GEN_21022 : _GEN_20646; // @[sequencer-master.scala 168:32]
  wire  _GEN_21031 = _T_1596 ? _GEN_21023 : _GEN_20647; // @[sequencer-master.scala 168:32]
  wire  _GEN_21032 = _T_1596 ? _GEN_21024 : _GEN_20648; // @[sequencer-master.scala 168:32]
  wire  _GEN_21033 = _T_1596 ? _GEN_21025 : _GEN_20649; // @[sequencer-master.scala 168:32]
  wire  _GEN_21034 = _T_1596 ? _GEN_21026 : _GEN_20650; // @[sequencer-master.scala 168:32]
  wire  _GEN_21035 = _T_1596 ? _GEN_21027 : _GEN_20651; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_21036 = 3'h0 == _T_1649 ? 2'h0 : _GEN_20308; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21037 = 3'h1 == _T_1649 ? 2'h0 : _GEN_20309; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21038 = 3'h2 == _T_1649 ? 2'h0 : _GEN_20310; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21039 = 3'h3 == _T_1649 ? 2'h0 : _GEN_20311; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21040 = 3'h4 == _T_1649 ? 2'h0 : _GEN_20312; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21041 = 3'h5 == _T_1649 ? 2'h0 : _GEN_20313; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21042 = 3'h6 == _T_1649 ? 2'h0 : _GEN_20314; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_21043 = 3'h7 == _T_1649 ? 2'h0 : _GEN_20315; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_21044 = 3'h0 == _T_1649 ? 4'h0 : _GEN_20316; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21045 = 3'h1 == _T_1649 ? 4'h0 : _GEN_20317; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21046 = 3'h2 == _T_1649 ? 4'h0 : _GEN_20318; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21047 = 3'h3 == _T_1649 ? 4'h0 : _GEN_20319; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21048 = 3'h4 == _T_1649 ? 4'h0 : _GEN_20320; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21049 = 3'h5 == _T_1649 ? 4'h0 : _GEN_20321; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21050 = 3'h6 == _T_1649 ? 4'h0 : _GEN_20322; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_21051 = 3'h7 == _T_1649 ? 4'h0 : _GEN_20323; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_21052 = 3'h0 == _T_1649 ? 3'h0 : _GEN_20324; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21053 = 3'h1 == _T_1649 ? 3'h0 : _GEN_20325; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21054 = 3'h2 == _T_1649 ? 3'h0 : _GEN_20326; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21055 = 3'h3 == _T_1649 ? 3'h0 : _GEN_20327; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21056 = 3'h4 == _T_1649 ? 3'h0 : _GEN_20328; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21057 = 3'h5 == _T_1649 ? 3'h0 : _GEN_20329; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21058 = 3'h6 == _T_1649 ? 3'h0 : _GEN_20330; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_21059 = 3'h7 == _T_1649 ? 3'h0 : _GEN_20331; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_21060 = io_op_bits_active_vamo ? _GEN_20396 : _GEN_17834; // @[sequencer-master.scala 650:39]
  wire  _GEN_21061 = io_op_bits_active_vamo ? _GEN_20397 : _GEN_17835; // @[sequencer-master.scala 650:39]
  wire  _GEN_21062 = io_op_bits_active_vamo ? _GEN_20398 : _GEN_17836; // @[sequencer-master.scala 650:39]
  wire  _GEN_21063 = io_op_bits_active_vamo ? _GEN_20399 : _GEN_17837; // @[sequencer-master.scala 650:39]
  wire  _GEN_21064 = io_op_bits_active_vamo ? _GEN_20400 : _GEN_17838; // @[sequencer-master.scala 650:39]
  wire  _GEN_21065 = io_op_bits_active_vamo ? _GEN_20401 : _GEN_17839; // @[sequencer-master.scala 650:39]
  wire  _GEN_21066 = io_op_bits_active_vamo ? _GEN_20402 : _GEN_17840; // @[sequencer-master.scala 650:39]
  wire  _GEN_21067 = io_op_bits_active_vamo ? _GEN_20403 : _GEN_17841; // @[sequencer-master.scala 650:39]
  wire  _GEN_21076 = io_op_bits_active_vamo ? _GEN_20412 : _GEN_17850; // @[sequencer-master.scala 650:39]
  wire  _GEN_21077 = io_op_bits_active_vamo ? _GEN_20413 : _GEN_17851; // @[sequencer-master.scala 650:39]
  wire  _GEN_21078 = io_op_bits_active_vamo ? _GEN_20414 : _GEN_17852; // @[sequencer-master.scala 650:39]
  wire  _GEN_21079 = io_op_bits_active_vamo ? _GEN_20415 : _GEN_17853; // @[sequencer-master.scala 650:39]
  wire  _GEN_21080 = io_op_bits_active_vamo ? _GEN_20416 : _GEN_17854; // @[sequencer-master.scala 650:39]
  wire  _GEN_21081 = io_op_bits_active_vamo ? _GEN_20417 : _GEN_17855; // @[sequencer-master.scala 650:39]
  wire  _GEN_21082 = io_op_bits_active_vamo ? _GEN_20418 : _GEN_17856; // @[sequencer-master.scala 650:39]
  wire  _GEN_21083 = io_op_bits_active_vamo ? _GEN_20419 : _GEN_17857; // @[sequencer-master.scala 650:39]
  wire  _GEN_21084 = io_op_bits_active_vamo ? _GEN_20420 : _GEN_17858; // @[sequencer-master.scala 650:39]
  wire  _GEN_21085 = io_op_bits_active_vamo ? _GEN_20421 : _GEN_17859; // @[sequencer-master.scala 650:39]
  wire  _GEN_21086 = io_op_bits_active_vamo ? _GEN_20422 : _GEN_17860; // @[sequencer-master.scala 650:39]
  wire  _GEN_21087 = io_op_bits_active_vamo ? _GEN_20423 : _GEN_17861; // @[sequencer-master.scala 650:39]
  wire  _GEN_21088 = io_op_bits_active_vamo ? _GEN_20424 : _GEN_17862; // @[sequencer-master.scala 650:39]
  wire  _GEN_21089 = io_op_bits_active_vamo ? _GEN_20425 : _GEN_17863; // @[sequencer-master.scala 650:39]
  wire  _GEN_21090 = io_op_bits_active_vamo ? _GEN_20426 : _GEN_17864; // @[sequencer-master.scala 650:39]
  wire  _GEN_21091 = io_op_bits_active_vamo ? _GEN_20427 : _GEN_17865; // @[sequencer-master.scala 650:39]
  wire  _GEN_21092 = io_op_bits_active_vamo ? _GEN_20428 : _GEN_17866; // @[sequencer-master.scala 650:39]
  wire  _GEN_21093 = io_op_bits_active_vamo ? _GEN_20429 : _GEN_17867; // @[sequencer-master.scala 650:39]
  wire  _GEN_21094 = io_op_bits_active_vamo ? _GEN_20430 : _GEN_17868; // @[sequencer-master.scala 650:39]
  wire  _GEN_21095 = io_op_bits_active_vamo ? _GEN_20431 : _GEN_17869; // @[sequencer-master.scala 650:39]
  wire  _GEN_21096 = io_op_bits_active_vamo ? _GEN_20432 : _GEN_17870; // @[sequencer-master.scala 650:39]
  wire  _GEN_21097 = io_op_bits_active_vamo ? _GEN_20433 : _GEN_17871; // @[sequencer-master.scala 650:39]
  wire  _GEN_21098 = io_op_bits_active_vamo ? _GEN_20434 : _GEN_17872; // @[sequencer-master.scala 650:39]
  wire  _GEN_21099 = io_op_bits_active_vamo ? _GEN_20435 : _GEN_17873; // @[sequencer-master.scala 650:39]
  wire  _GEN_21100 = io_op_bits_active_vamo ? _GEN_20436 : _GEN_17874; // @[sequencer-master.scala 650:39]
  wire  _GEN_21101 = io_op_bits_active_vamo ? _GEN_20437 : _GEN_17875; // @[sequencer-master.scala 650:39]
  wire  _GEN_21102 = io_op_bits_active_vamo ? _GEN_20438 : _GEN_17876; // @[sequencer-master.scala 650:39]
  wire  _GEN_21103 = io_op_bits_active_vamo ? _GEN_20439 : _GEN_17877; // @[sequencer-master.scala 650:39]
  wire  _GEN_21104 = io_op_bits_active_vamo ? _GEN_20440 : _GEN_17878; // @[sequencer-master.scala 650:39]
  wire  _GEN_21105 = io_op_bits_active_vamo ? _GEN_20441 : _GEN_17879; // @[sequencer-master.scala 650:39]
  wire  _GEN_21106 = io_op_bits_active_vamo ? _GEN_20442 : _GEN_17880; // @[sequencer-master.scala 650:39]
  wire  _GEN_21107 = io_op_bits_active_vamo ? _GEN_20443 : _GEN_17881; // @[sequencer-master.scala 650:39]
  wire  _GEN_21108 = io_op_bits_active_vamo ? _GEN_20740 : _GEN_17882; // @[sequencer-master.scala 650:39]
  wire  _GEN_21109 = io_op_bits_active_vamo ? _GEN_20741 : _GEN_17883; // @[sequencer-master.scala 650:39]
  wire  _GEN_21110 = io_op_bits_active_vamo ? _GEN_20742 : _GEN_17884; // @[sequencer-master.scala 650:39]
  wire  _GEN_21111 = io_op_bits_active_vamo ? _GEN_20743 : _GEN_17885; // @[sequencer-master.scala 650:39]
  wire  _GEN_21112 = io_op_bits_active_vamo ? _GEN_20744 : _GEN_17886; // @[sequencer-master.scala 650:39]
  wire  _GEN_21113 = io_op_bits_active_vamo ? _GEN_20745 : _GEN_17887; // @[sequencer-master.scala 650:39]
  wire  _GEN_21114 = io_op_bits_active_vamo ? _GEN_20746 : _GEN_17888; // @[sequencer-master.scala 650:39]
  wire  _GEN_21115 = io_op_bits_active_vamo ? _GEN_20747 : _GEN_17889; // @[sequencer-master.scala 650:39]
  wire  _GEN_21116 = io_op_bits_active_vamo ? _GEN_20452 : _GEN_17890; // @[sequencer-master.scala 650:39]
  wire  _GEN_21117 = io_op_bits_active_vamo ? _GEN_20453 : _GEN_17891; // @[sequencer-master.scala 650:39]
  wire  _GEN_21118 = io_op_bits_active_vamo ? _GEN_20454 : _GEN_17892; // @[sequencer-master.scala 650:39]
  wire  _GEN_21119 = io_op_bits_active_vamo ? _GEN_20455 : _GEN_17893; // @[sequencer-master.scala 650:39]
  wire  _GEN_21120 = io_op_bits_active_vamo ? _GEN_20456 : _GEN_17894; // @[sequencer-master.scala 650:39]
  wire  _GEN_21121 = io_op_bits_active_vamo ? _GEN_20457 : _GEN_17895; // @[sequencer-master.scala 650:39]
  wire  _GEN_21122 = io_op_bits_active_vamo ? _GEN_20458 : _GEN_17896; // @[sequencer-master.scala 650:39]
  wire  _GEN_21123 = io_op_bits_active_vamo ? _GEN_20459 : _GEN_17897; // @[sequencer-master.scala 650:39]
  wire  _GEN_21124 = io_op_bits_active_vamo ? _GEN_20460 : _GEN_17898; // @[sequencer-master.scala 650:39]
  wire  _GEN_21125 = io_op_bits_active_vamo ? _GEN_20461 : _GEN_17899; // @[sequencer-master.scala 650:39]
  wire  _GEN_21126 = io_op_bits_active_vamo ? _GEN_20462 : _GEN_17900; // @[sequencer-master.scala 650:39]
  wire  _GEN_21127 = io_op_bits_active_vamo ? _GEN_20463 : _GEN_17901; // @[sequencer-master.scala 650:39]
  wire  _GEN_21128 = io_op_bits_active_vamo ? _GEN_20464 : _GEN_17902; // @[sequencer-master.scala 650:39]
  wire  _GEN_21129 = io_op_bits_active_vamo ? _GEN_20465 : _GEN_17903; // @[sequencer-master.scala 650:39]
  wire  _GEN_21130 = io_op_bits_active_vamo ? _GEN_20466 : _GEN_17904; // @[sequencer-master.scala 650:39]
  wire  _GEN_21131 = io_op_bits_active_vamo ? _GEN_20467 : _GEN_17905; // @[sequencer-master.scala 650:39]
  wire  _GEN_21132 = io_op_bits_active_vamo ? _GEN_20788 : _GEN_17906; // @[sequencer-master.scala 650:39]
  wire  _GEN_21133 = io_op_bits_active_vamo ? _GEN_20789 : _GEN_17907; // @[sequencer-master.scala 650:39]
  wire  _GEN_21134 = io_op_bits_active_vamo ? _GEN_20790 : _GEN_17908; // @[sequencer-master.scala 650:39]
  wire  _GEN_21135 = io_op_bits_active_vamo ? _GEN_20791 : _GEN_17909; // @[sequencer-master.scala 650:39]
  wire  _GEN_21136 = io_op_bits_active_vamo ? _GEN_20792 : _GEN_17910; // @[sequencer-master.scala 650:39]
  wire  _GEN_21137 = io_op_bits_active_vamo ? _GEN_20793 : _GEN_17911; // @[sequencer-master.scala 650:39]
  wire  _GEN_21138 = io_op_bits_active_vamo ? _GEN_20794 : _GEN_17912; // @[sequencer-master.scala 650:39]
  wire  _GEN_21139 = io_op_bits_active_vamo ? _GEN_20795 : _GEN_17913; // @[sequencer-master.scala 650:39]
  wire  _GEN_21140 = io_op_bits_active_vamo ? _GEN_20916 : _GEN_17914; // @[sequencer-master.scala 650:39]
  wire  _GEN_21141 = io_op_bits_active_vamo ? _GEN_20917 : _GEN_17915; // @[sequencer-master.scala 650:39]
  wire  _GEN_21142 = io_op_bits_active_vamo ? _GEN_20918 : _GEN_17916; // @[sequencer-master.scala 650:39]
  wire  _GEN_21143 = io_op_bits_active_vamo ? _GEN_20919 : _GEN_17917; // @[sequencer-master.scala 650:39]
  wire  _GEN_21144 = io_op_bits_active_vamo ? _GEN_20920 : _GEN_17918; // @[sequencer-master.scala 650:39]
  wire  _GEN_21145 = io_op_bits_active_vamo ? _GEN_20921 : _GEN_17919; // @[sequencer-master.scala 650:39]
  wire  _GEN_21146 = io_op_bits_active_vamo ? _GEN_20922 : _GEN_17920; // @[sequencer-master.scala 650:39]
  wire  _GEN_21147 = io_op_bits_active_vamo ? _GEN_20923 : _GEN_17921; // @[sequencer-master.scala 650:39]
  wire  _GEN_21148 = io_op_bits_active_vamo ? _GEN_20484 : _GEN_17922; // @[sequencer-master.scala 650:39]
  wire  _GEN_21149 = io_op_bits_active_vamo ? _GEN_20485 : _GEN_17923; // @[sequencer-master.scala 650:39]
  wire  _GEN_21150 = io_op_bits_active_vamo ? _GEN_20486 : _GEN_17924; // @[sequencer-master.scala 650:39]
  wire  _GEN_21151 = io_op_bits_active_vamo ? _GEN_20487 : _GEN_17925; // @[sequencer-master.scala 650:39]
  wire  _GEN_21152 = io_op_bits_active_vamo ? _GEN_20488 : _GEN_17926; // @[sequencer-master.scala 650:39]
  wire  _GEN_21153 = io_op_bits_active_vamo ? _GEN_20489 : _GEN_17927; // @[sequencer-master.scala 650:39]
  wire  _GEN_21154 = io_op_bits_active_vamo ? _GEN_20490 : _GEN_17928; // @[sequencer-master.scala 650:39]
  wire  _GEN_21155 = io_op_bits_active_vamo ? _GEN_20491 : _GEN_17929; // @[sequencer-master.scala 650:39]
  wire  _GEN_21156 = io_op_bits_active_vamo ? _GEN_20804 : _GEN_17930; // @[sequencer-master.scala 650:39]
  wire  _GEN_21157 = io_op_bits_active_vamo ? _GEN_20805 : _GEN_17931; // @[sequencer-master.scala 650:39]
  wire  _GEN_21158 = io_op_bits_active_vamo ? _GEN_20806 : _GEN_17932; // @[sequencer-master.scala 650:39]
  wire  _GEN_21159 = io_op_bits_active_vamo ? _GEN_20807 : _GEN_17933; // @[sequencer-master.scala 650:39]
  wire  _GEN_21160 = io_op_bits_active_vamo ? _GEN_20808 : _GEN_17934; // @[sequencer-master.scala 650:39]
  wire  _GEN_21161 = io_op_bits_active_vamo ? _GEN_20809 : _GEN_17935; // @[sequencer-master.scala 650:39]
  wire  _GEN_21162 = io_op_bits_active_vamo ? _GEN_20810 : _GEN_17936; // @[sequencer-master.scala 650:39]
  wire  _GEN_21163 = io_op_bits_active_vamo ? _GEN_20811 : _GEN_17937; // @[sequencer-master.scala 650:39]
  wire  _GEN_21164 = io_op_bits_active_vamo ? _GEN_20932 : _GEN_17938; // @[sequencer-master.scala 650:39]
  wire  _GEN_21165 = io_op_bits_active_vamo ? _GEN_20933 : _GEN_17939; // @[sequencer-master.scala 650:39]
  wire  _GEN_21166 = io_op_bits_active_vamo ? _GEN_20934 : _GEN_17940; // @[sequencer-master.scala 650:39]
  wire  _GEN_21167 = io_op_bits_active_vamo ? _GEN_20935 : _GEN_17941; // @[sequencer-master.scala 650:39]
  wire  _GEN_21168 = io_op_bits_active_vamo ? _GEN_20936 : _GEN_17942; // @[sequencer-master.scala 650:39]
  wire  _GEN_21169 = io_op_bits_active_vamo ? _GEN_20937 : _GEN_17943; // @[sequencer-master.scala 650:39]
  wire  _GEN_21170 = io_op_bits_active_vamo ? _GEN_20938 : _GEN_17944; // @[sequencer-master.scala 650:39]
  wire  _GEN_21171 = io_op_bits_active_vamo ? _GEN_20939 : _GEN_17945; // @[sequencer-master.scala 650:39]
  wire  _GEN_21172 = io_op_bits_active_vamo ? _GEN_20508 : _GEN_17946; // @[sequencer-master.scala 650:39]
  wire  _GEN_21173 = io_op_bits_active_vamo ? _GEN_20509 : _GEN_17947; // @[sequencer-master.scala 650:39]
  wire  _GEN_21174 = io_op_bits_active_vamo ? _GEN_20510 : _GEN_17948; // @[sequencer-master.scala 650:39]
  wire  _GEN_21175 = io_op_bits_active_vamo ? _GEN_20511 : _GEN_17949; // @[sequencer-master.scala 650:39]
  wire  _GEN_21176 = io_op_bits_active_vamo ? _GEN_20512 : _GEN_17950; // @[sequencer-master.scala 650:39]
  wire  _GEN_21177 = io_op_bits_active_vamo ? _GEN_20513 : _GEN_17951; // @[sequencer-master.scala 650:39]
  wire  _GEN_21178 = io_op_bits_active_vamo ? _GEN_20514 : _GEN_17952; // @[sequencer-master.scala 650:39]
  wire  _GEN_21179 = io_op_bits_active_vamo ? _GEN_20515 : _GEN_17953; // @[sequencer-master.scala 650:39]
  wire  _GEN_21180 = io_op_bits_active_vamo ? _GEN_20820 : _GEN_17954; // @[sequencer-master.scala 650:39]
  wire  _GEN_21181 = io_op_bits_active_vamo ? _GEN_20821 : _GEN_17955; // @[sequencer-master.scala 650:39]
  wire  _GEN_21182 = io_op_bits_active_vamo ? _GEN_20822 : _GEN_17956; // @[sequencer-master.scala 650:39]
  wire  _GEN_21183 = io_op_bits_active_vamo ? _GEN_20823 : _GEN_17957; // @[sequencer-master.scala 650:39]
  wire  _GEN_21184 = io_op_bits_active_vamo ? _GEN_20824 : _GEN_17958; // @[sequencer-master.scala 650:39]
  wire  _GEN_21185 = io_op_bits_active_vamo ? _GEN_20825 : _GEN_17959; // @[sequencer-master.scala 650:39]
  wire  _GEN_21186 = io_op_bits_active_vamo ? _GEN_20826 : _GEN_17960; // @[sequencer-master.scala 650:39]
  wire  _GEN_21187 = io_op_bits_active_vamo ? _GEN_20827 : _GEN_17961; // @[sequencer-master.scala 650:39]
  wire  _GEN_21188 = io_op_bits_active_vamo ? _GEN_20948 : _GEN_17962; // @[sequencer-master.scala 650:39]
  wire  _GEN_21189 = io_op_bits_active_vamo ? _GEN_20949 : _GEN_17963; // @[sequencer-master.scala 650:39]
  wire  _GEN_21190 = io_op_bits_active_vamo ? _GEN_20950 : _GEN_17964; // @[sequencer-master.scala 650:39]
  wire  _GEN_21191 = io_op_bits_active_vamo ? _GEN_20951 : _GEN_17965; // @[sequencer-master.scala 650:39]
  wire  _GEN_21192 = io_op_bits_active_vamo ? _GEN_20952 : _GEN_17966; // @[sequencer-master.scala 650:39]
  wire  _GEN_21193 = io_op_bits_active_vamo ? _GEN_20953 : _GEN_17967; // @[sequencer-master.scala 650:39]
  wire  _GEN_21194 = io_op_bits_active_vamo ? _GEN_20954 : _GEN_17968; // @[sequencer-master.scala 650:39]
  wire  _GEN_21195 = io_op_bits_active_vamo ? _GEN_20955 : _GEN_17969; // @[sequencer-master.scala 650:39]
  wire  _GEN_21196 = io_op_bits_active_vamo ? _GEN_20532 : _GEN_17970; // @[sequencer-master.scala 650:39]
  wire  _GEN_21197 = io_op_bits_active_vamo ? _GEN_20533 : _GEN_17971; // @[sequencer-master.scala 650:39]
  wire  _GEN_21198 = io_op_bits_active_vamo ? _GEN_20534 : _GEN_17972; // @[sequencer-master.scala 650:39]
  wire  _GEN_21199 = io_op_bits_active_vamo ? _GEN_20535 : _GEN_17973; // @[sequencer-master.scala 650:39]
  wire  _GEN_21200 = io_op_bits_active_vamo ? _GEN_20536 : _GEN_17974; // @[sequencer-master.scala 650:39]
  wire  _GEN_21201 = io_op_bits_active_vamo ? _GEN_20537 : _GEN_17975; // @[sequencer-master.scala 650:39]
  wire  _GEN_21202 = io_op_bits_active_vamo ? _GEN_20538 : _GEN_17976; // @[sequencer-master.scala 650:39]
  wire  _GEN_21203 = io_op_bits_active_vamo ? _GEN_20539 : _GEN_17977; // @[sequencer-master.scala 650:39]
  wire  _GEN_21204 = io_op_bits_active_vamo ? _GEN_20836 : _GEN_17978; // @[sequencer-master.scala 650:39]
  wire  _GEN_21205 = io_op_bits_active_vamo ? _GEN_20837 : _GEN_17979; // @[sequencer-master.scala 650:39]
  wire  _GEN_21206 = io_op_bits_active_vamo ? _GEN_20838 : _GEN_17980; // @[sequencer-master.scala 650:39]
  wire  _GEN_21207 = io_op_bits_active_vamo ? _GEN_20839 : _GEN_17981; // @[sequencer-master.scala 650:39]
  wire  _GEN_21208 = io_op_bits_active_vamo ? _GEN_20840 : _GEN_17982; // @[sequencer-master.scala 650:39]
  wire  _GEN_21209 = io_op_bits_active_vamo ? _GEN_20841 : _GEN_17983; // @[sequencer-master.scala 650:39]
  wire  _GEN_21210 = io_op_bits_active_vamo ? _GEN_20842 : _GEN_17984; // @[sequencer-master.scala 650:39]
  wire  _GEN_21211 = io_op_bits_active_vamo ? _GEN_20843 : _GEN_17985; // @[sequencer-master.scala 650:39]
  wire  _GEN_21212 = io_op_bits_active_vamo ? _GEN_20964 : _GEN_17986; // @[sequencer-master.scala 650:39]
  wire  _GEN_21213 = io_op_bits_active_vamo ? _GEN_20965 : _GEN_17987; // @[sequencer-master.scala 650:39]
  wire  _GEN_21214 = io_op_bits_active_vamo ? _GEN_20966 : _GEN_17988; // @[sequencer-master.scala 650:39]
  wire  _GEN_21215 = io_op_bits_active_vamo ? _GEN_20967 : _GEN_17989; // @[sequencer-master.scala 650:39]
  wire  _GEN_21216 = io_op_bits_active_vamo ? _GEN_20968 : _GEN_17990; // @[sequencer-master.scala 650:39]
  wire  _GEN_21217 = io_op_bits_active_vamo ? _GEN_20969 : _GEN_17991; // @[sequencer-master.scala 650:39]
  wire  _GEN_21218 = io_op_bits_active_vamo ? _GEN_20970 : _GEN_17992; // @[sequencer-master.scala 650:39]
  wire  _GEN_21219 = io_op_bits_active_vamo ? _GEN_20971 : _GEN_17993; // @[sequencer-master.scala 650:39]
  wire  _GEN_21220 = io_op_bits_active_vamo ? _GEN_20556 : _GEN_17994; // @[sequencer-master.scala 650:39]
  wire  _GEN_21221 = io_op_bits_active_vamo ? _GEN_20557 : _GEN_17995; // @[sequencer-master.scala 650:39]
  wire  _GEN_21222 = io_op_bits_active_vamo ? _GEN_20558 : _GEN_17996; // @[sequencer-master.scala 650:39]
  wire  _GEN_21223 = io_op_bits_active_vamo ? _GEN_20559 : _GEN_17997; // @[sequencer-master.scala 650:39]
  wire  _GEN_21224 = io_op_bits_active_vamo ? _GEN_20560 : _GEN_17998; // @[sequencer-master.scala 650:39]
  wire  _GEN_21225 = io_op_bits_active_vamo ? _GEN_20561 : _GEN_17999; // @[sequencer-master.scala 650:39]
  wire  _GEN_21226 = io_op_bits_active_vamo ? _GEN_20562 : _GEN_18000; // @[sequencer-master.scala 650:39]
  wire  _GEN_21227 = io_op_bits_active_vamo ? _GEN_20563 : _GEN_18001; // @[sequencer-master.scala 650:39]
  wire  _GEN_21228 = io_op_bits_active_vamo ? _GEN_20852 : _GEN_18002; // @[sequencer-master.scala 650:39]
  wire  _GEN_21229 = io_op_bits_active_vamo ? _GEN_20853 : _GEN_18003; // @[sequencer-master.scala 650:39]
  wire  _GEN_21230 = io_op_bits_active_vamo ? _GEN_20854 : _GEN_18004; // @[sequencer-master.scala 650:39]
  wire  _GEN_21231 = io_op_bits_active_vamo ? _GEN_20855 : _GEN_18005; // @[sequencer-master.scala 650:39]
  wire  _GEN_21232 = io_op_bits_active_vamo ? _GEN_20856 : _GEN_18006; // @[sequencer-master.scala 650:39]
  wire  _GEN_21233 = io_op_bits_active_vamo ? _GEN_20857 : _GEN_18007; // @[sequencer-master.scala 650:39]
  wire  _GEN_21234 = io_op_bits_active_vamo ? _GEN_20858 : _GEN_18008; // @[sequencer-master.scala 650:39]
  wire  _GEN_21235 = io_op_bits_active_vamo ? _GEN_20859 : _GEN_18009; // @[sequencer-master.scala 650:39]
  wire  _GEN_21236 = io_op_bits_active_vamo ? _GEN_20980 : _GEN_18010; // @[sequencer-master.scala 650:39]
  wire  _GEN_21237 = io_op_bits_active_vamo ? _GEN_20981 : _GEN_18011; // @[sequencer-master.scala 650:39]
  wire  _GEN_21238 = io_op_bits_active_vamo ? _GEN_20982 : _GEN_18012; // @[sequencer-master.scala 650:39]
  wire  _GEN_21239 = io_op_bits_active_vamo ? _GEN_20983 : _GEN_18013; // @[sequencer-master.scala 650:39]
  wire  _GEN_21240 = io_op_bits_active_vamo ? _GEN_20984 : _GEN_18014; // @[sequencer-master.scala 650:39]
  wire  _GEN_21241 = io_op_bits_active_vamo ? _GEN_20985 : _GEN_18015; // @[sequencer-master.scala 650:39]
  wire  _GEN_21242 = io_op_bits_active_vamo ? _GEN_20986 : _GEN_18016; // @[sequencer-master.scala 650:39]
  wire  _GEN_21243 = io_op_bits_active_vamo ? _GEN_20987 : _GEN_18017; // @[sequencer-master.scala 650:39]
  wire  _GEN_21244 = io_op_bits_active_vamo ? _GEN_20580 : _GEN_18018; // @[sequencer-master.scala 650:39]
  wire  _GEN_21245 = io_op_bits_active_vamo ? _GEN_20581 : _GEN_18019; // @[sequencer-master.scala 650:39]
  wire  _GEN_21246 = io_op_bits_active_vamo ? _GEN_20582 : _GEN_18020; // @[sequencer-master.scala 650:39]
  wire  _GEN_21247 = io_op_bits_active_vamo ? _GEN_20583 : _GEN_18021; // @[sequencer-master.scala 650:39]
  wire  _GEN_21248 = io_op_bits_active_vamo ? _GEN_20584 : _GEN_18022; // @[sequencer-master.scala 650:39]
  wire  _GEN_21249 = io_op_bits_active_vamo ? _GEN_20585 : _GEN_18023; // @[sequencer-master.scala 650:39]
  wire  _GEN_21250 = io_op_bits_active_vamo ? _GEN_20586 : _GEN_18024; // @[sequencer-master.scala 650:39]
  wire  _GEN_21251 = io_op_bits_active_vamo ? _GEN_20587 : _GEN_18025; // @[sequencer-master.scala 650:39]
  wire  _GEN_21252 = io_op_bits_active_vamo ? _GEN_20868 : _GEN_18026; // @[sequencer-master.scala 650:39]
  wire  _GEN_21253 = io_op_bits_active_vamo ? _GEN_20869 : _GEN_18027; // @[sequencer-master.scala 650:39]
  wire  _GEN_21254 = io_op_bits_active_vamo ? _GEN_20870 : _GEN_18028; // @[sequencer-master.scala 650:39]
  wire  _GEN_21255 = io_op_bits_active_vamo ? _GEN_20871 : _GEN_18029; // @[sequencer-master.scala 650:39]
  wire  _GEN_21256 = io_op_bits_active_vamo ? _GEN_20872 : _GEN_18030; // @[sequencer-master.scala 650:39]
  wire  _GEN_21257 = io_op_bits_active_vamo ? _GEN_20873 : _GEN_18031; // @[sequencer-master.scala 650:39]
  wire  _GEN_21258 = io_op_bits_active_vamo ? _GEN_20874 : _GEN_18032; // @[sequencer-master.scala 650:39]
  wire  _GEN_21259 = io_op_bits_active_vamo ? _GEN_20875 : _GEN_18033; // @[sequencer-master.scala 650:39]
  wire  _GEN_21260 = io_op_bits_active_vamo ? _GEN_20996 : _GEN_18034; // @[sequencer-master.scala 650:39]
  wire  _GEN_21261 = io_op_bits_active_vamo ? _GEN_20997 : _GEN_18035; // @[sequencer-master.scala 650:39]
  wire  _GEN_21262 = io_op_bits_active_vamo ? _GEN_20998 : _GEN_18036; // @[sequencer-master.scala 650:39]
  wire  _GEN_21263 = io_op_bits_active_vamo ? _GEN_20999 : _GEN_18037; // @[sequencer-master.scala 650:39]
  wire  _GEN_21264 = io_op_bits_active_vamo ? _GEN_21000 : _GEN_18038; // @[sequencer-master.scala 650:39]
  wire  _GEN_21265 = io_op_bits_active_vamo ? _GEN_21001 : _GEN_18039; // @[sequencer-master.scala 650:39]
  wire  _GEN_21266 = io_op_bits_active_vamo ? _GEN_21002 : _GEN_18040; // @[sequencer-master.scala 650:39]
  wire  _GEN_21267 = io_op_bits_active_vamo ? _GEN_21003 : _GEN_18041; // @[sequencer-master.scala 650:39]
  wire  _GEN_21268 = io_op_bits_active_vamo ? _GEN_20604 : _GEN_18042; // @[sequencer-master.scala 650:39]
  wire  _GEN_21269 = io_op_bits_active_vamo ? _GEN_20605 : _GEN_18043; // @[sequencer-master.scala 650:39]
  wire  _GEN_21270 = io_op_bits_active_vamo ? _GEN_20606 : _GEN_18044; // @[sequencer-master.scala 650:39]
  wire  _GEN_21271 = io_op_bits_active_vamo ? _GEN_20607 : _GEN_18045; // @[sequencer-master.scala 650:39]
  wire  _GEN_21272 = io_op_bits_active_vamo ? _GEN_20608 : _GEN_18046; // @[sequencer-master.scala 650:39]
  wire  _GEN_21273 = io_op_bits_active_vamo ? _GEN_20609 : _GEN_18047; // @[sequencer-master.scala 650:39]
  wire  _GEN_21274 = io_op_bits_active_vamo ? _GEN_20610 : _GEN_18048; // @[sequencer-master.scala 650:39]
  wire  _GEN_21275 = io_op_bits_active_vamo ? _GEN_20611 : _GEN_18049; // @[sequencer-master.scala 650:39]
  wire  _GEN_21276 = io_op_bits_active_vamo ? _GEN_20884 : _GEN_18050; // @[sequencer-master.scala 650:39]
  wire  _GEN_21277 = io_op_bits_active_vamo ? _GEN_20885 : _GEN_18051; // @[sequencer-master.scala 650:39]
  wire  _GEN_21278 = io_op_bits_active_vamo ? _GEN_20886 : _GEN_18052; // @[sequencer-master.scala 650:39]
  wire  _GEN_21279 = io_op_bits_active_vamo ? _GEN_20887 : _GEN_18053; // @[sequencer-master.scala 650:39]
  wire  _GEN_21280 = io_op_bits_active_vamo ? _GEN_20888 : _GEN_18054; // @[sequencer-master.scala 650:39]
  wire  _GEN_21281 = io_op_bits_active_vamo ? _GEN_20889 : _GEN_18055; // @[sequencer-master.scala 650:39]
  wire  _GEN_21282 = io_op_bits_active_vamo ? _GEN_20890 : _GEN_18056; // @[sequencer-master.scala 650:39]
  wire  _GEN_21283 = io_op_bits_active_vamo ? _GEN_20891 : _GEN_18057; // @[sequencer-master.scala 650:39]
  wire  _GEN_21284 = io_op_bits_active_vamo ? _GEN_21012 : _GEN_18058; // @[sequencer-master.scala 650:39]
  wire  _GEN_21285 = io_op_bits_active_vamo ? _GEN_21013 : _GEN_18059; // @[sequencer-master.scala 650:39]
  wire  _GEN_21286 = io_op_bits_active_vamo ? _GEN_21014 : _GEN_18060; // @[sequencer-master.scala 650:39]
  wire  _GEN_21287 = io_op_bits_active_vamo ? _GEN_21015 : _GEN_18061; // @[sequencer-master.scala 650:39]
  wire  _GEN_21288 = io_op_bits_active_vamo ? _GEN_21016 : _GEN_18062; // @[sequencer-master.scala 650:39]
  wire  _GEN_21289 = io_op_bits_active_vamo ? _GEN_21017 : _GEN_18063; // @[sequencer-master.scala 650:39]
  wire  _GEN_21290 = io_op_bits_active_vamo ? _GEN_21018 : _GEN_18064; // @[sequencer-master.scala 650:39]
  wire  _GEN_21291 = io_op_bits_active_vamo ? _GEN_21019 : _GEN_18065; // @[sequencer-master.scala 650:39]
  wire  _GEN_21292 = io_op_bits_active_vamo ? _GEN_20628 : _GEN_18066; // @[sequencer-master.scala 650:39]
  wire  _GEN_21293 = io_op_bits_active_vamo ? _GEN_20629 : _GEN_18067; // @[sequencer-master.scala 650:39]
  wire  _GEN_21294 = io_op_bits_active_vamo ? _GEN_20630 : _GEN_18068; // @[sequencer-master.scala 650:39]
  wire  _GEN_21295 = io_op_bits_active_vamo ? _GEN_20631 : _GEN_18069; // @[sequencer-master.scala 650:39]
  wire  _GEN_21296 = io_op_bits_active_vamo ? _GEN_20632 : _GEN_18070; // @[sequencer-master.scala 650:39]
  wire  _GEN_21297 = io_op_bits_active_vamo ? _GEN_20633 : _GEN_18071; // @[sequencer-master.scala 650:39]
  wire  _GEN_21298 = io_op_bits_active_vamo ? _GEN_20634 : _GEN_18072; // @[sequencer-master.scala 650:39]
  wire  _GEN_21299 = io_op_bits_active_vamo ? _GEN_20635 : _GEN_18073; // @[sequencer-master.scala 650:39]
  wire  _GEN_21300 = io_op_bits_active_vamo ? _GEN_20900 : _GEN_18074; // @[sequencer-master.scala 650:39]
  wire  _GEN_21301 = io_op_bits_active_vamo ? _GEN_20901 : _GEN_18075; // @[sequencer-master.scala 650:39]
  wire  _GEN_21302 = io_op_bits_active_vamo ? _GEN_20902 : _GEN_18076; // @[sequencer-master.scala 650:39]
  wire  _GEN_21303 = io_op_bits_active_vamo ? _GEN_20903 : _GEN_18077; // @[sequencer-master.scala 650:39]
  wire  _GEN_21304 = io_op_bits_active_vamo ? _GEN_20904 : _GEN_18078; // @[sequencer-master.scala 650:39]
  wire  _GEN_21305 = io_op_bits_active_vamo ? _GEN_20905 : _GEN_18079; // @[sequencer-master.scala 650:39]
  wire  _GEN_21306 = io_op_bits_active_vamo ? _GEN_20906 : _GEN_18080; // @[sequencer-master.scala 650:39]
  wire  _GEN_21307 = io_op_bits_active_vamo ? _GEN_20907 : _GEN_18081; // @[sequencer-master.scala 650:39]
  wire  _GEN_21308 = io_op_bits_active_vamo ? _GEN_21028 : _GEN_18082; // @[sequencer-master.scala 650:39]
  wire  _GEN_21309 = io_op_bits_active_vamo ? _GEN_21029 : _GEN_18083; // @[sequencer-master.scala 650:39]
  wire  _GEN_21310 = io_op_bits_active_vamo ? _GEN_21030 : _GEN_18084; // @[sequencer-master.scala 650:39]
  wire  _GEN_21311 = io_op_bits_active_vamo ? _GEN_21031 : _GEN_18085; // @[sequencer-master.scala 650:39]
  wire  _GEN_21312 = io_op_bits_active_vamo ? _GEN_21032 : _GEN_18086; // @[sequencer-master.scala 650:39]
  wire  _GEN_21313 = io_op_bits_active_vamo ? _GEN_21033 : _GEN_18087; // @[sequencer-master.scala 650:39]
  wire  _GEN_21314 = io_op_bits_active_vamo ? _GEN_21034 : _GEN_18088; // @[sequencer-master.scala 650:39]
  wire  _GEN_21315 = io_op_bits_active_vamo ? _GEN_21035 : _GEN_18089; // @[sequencer-master.scala 650:39]
  wire  _GEN_21316 = io_op_bits_active_vamo ? _GEN_20652 : _GEN_18090; // @[sequencer-master.scala 650:39]
  wire  _GEN_21317 = io_op_bits_active_vamo ? _GEN_20653 : _GEN_18091; // @[sequencer-master.scala 650:39]
  wire  _GEN_21318 = io_op_bits_active_vamo ? _GEN_20654 : _GEN_18092; // @[sequencer-master.scala 650:39]
  wire  _GEN_21319 = io_op_bits_active_vamo ? _GEN_20655 : _GEN_18093; // @[sequencer-master.scala 650:39]
  wire  _GEN_21320 = io_op_bits_active_vamo ? _GEN_20656 : _GEN_18094; // @[sequencer-master.scala 650:39]
  wire  _GEN_21321 = io_op_bits_active_vamo ? _GEN_20657 : _GEN_18095; // @[sequencer-master.scala 650:39]
  wire  _GEN_21322 = io_op_bits_active_vamo ? _GEN_20658 : _GEN_18096; // @[sequencer-master.scala 650:39]
  wire  _GEN_21323 = io_op_bits_active_vamo ? _GEN_20659 : _GEN_18097; // @[sequencer-master.scala 650:39]
  wire  _GEN_21332 = io_op_bits_active_vamo ? _GEN_18500 : e_0_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21333 = io_op_bits_active_vamo ? _GEN_18501 : e_1_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21334 = io_op_bits_active_vamo ? _GEN_18502 : e_2_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21335 = io_op_bits_active_vamo ? _GEN_18503 : e_3_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21336 = io_op_bits_active_vamo ? _GEN_18504 : e_4_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21337 = io_op_bits_active_vamo ? _GEN_18505 : e_5_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21338 = io_op_bits_active_vamo ? _GEN_18506 : e_6_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21339 = io_op_bits_active_vamo ? _GEN_18507 : e_7_active_vgu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire [9:0] _GEN_21340 = io_op_bits_active_vamo ? _GEN_20676 : _GEN_18114; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21341 = io_op_bits_active_vamo ? _GEN_20677 : _GEN_18115; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21342 = io_op_bits_active_vamo ? _GEN_20678 : _GEN_18116; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21343 = io_op_bits_active_vamo ? _GEN_20679 : _GEN_18117; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21344 = io_op_bits_active_vamo ? _GEN_20680 : _GEN_18118; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21345 = io_op_bits_active_vamo ? _GEN_20681 : _GEN_18119; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21346 = io_op_bits_active_vamo ? _GEN_20682 : _GEN_18120; // @[sequencer-master.scala 650:39]
  wire [9:0] _GEN_21347 = io_op_bits_active_vamo ? _GEN_20683 : _GEN_18121; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21348 = io_op_bits_active_vamo ? _GEN_19892 : _GEN_18122; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21349 = io_op_bits_active_vamo ? _GEN_19893 : _GEN_18123; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21350 = io_op_bits_active_vamo ? _GEN_19894 : _GEN_18124; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21351 = io_op_bits_active_vamo ? _GEN_19895 : _GEN_18125; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21352 = io_op_bits_active_vamo ? _GEN_19896 : _GEN_18126; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21353 = io_op_bits_active_vamo ? _GEN_19897 : _GEN_18127; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21354 = io_op_bits_active_vamo ? _GEN_19898 : _GEN_18128; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21355 = io_op_bits_active_vamo ? _GEN_19899 : _GEN_18129; // @[sequencer-master.scala 650:39]
  wire  _GEN_21356 = io_op_bits_active_vamo ? _GEN_19908 : _GEN_18130; // @[sequencer-master.scala 650:39]
  wire  _GEN_21357 = io_op_bits_active_vamo ? _GEN_19909 : _GEN_18131; // @[sequencer-master.scala 650:39]
  wire  _GEN_21358 = io_op_bits_active_vamo ? _GEN_19910 : _GEN_18132; // @[sequencer-master.scala 650:39]
  wire  _GEN_21359 = io_op_bits_active_vamo ? _GEN_19911 : _GEN_18133; // @[sequencer-master.scala 650:39]
  wire  _GEN_21360 = io_op_bits_active_vamo ? _GEN_19912 : _GEN_18134; // @[sequencer-master.scala 650:39]
  wire  _GEN_21361 = io_op_bits_active_vamo ? _GEN_19913 : _GEN_18135; // @[sequencer-master.scala 650:39]
  wire  _GEN_21362 = io_op_bits_active_vamo ? _GEN_19914 : _GEN_18136; // @[sequencer-master.scala 650:39]
  wire  _GEN_21363 = io_op_bits_active_vamo ? _GEN_19915 : _GEN_18137; // @[sequencer-master.scala 650:39]
  wire  _GEN_21364 = io_op_bits_active_vamo ? _GEN_19916 : _GEN_18138; // @[sequencer-master.scala 650:39]
  wire  _GEN_21365 = io_op_bits_active_vamo ? _GEN_19917 : _GEN_18139; // @[sequencer-master.scala 650:39]
  wire  _GEN_21366 = io_op_bits_active_vamo ? _GEN_19918 : _GEN_18140; // @[sequencer-master.scala 650:39]
  wire  _GEN_21367 = io_op_bits_active_vamo ? _GEN_19919 : _GEN_18141; // @[sequencer-master.scala 650:39]
  wire  _GEN_21368 = io_op_bits_active_vamo ? _GEN_19920 : _GEN_18142; // @[sequencer-master.scala 650:39]
  wire  _GEN_21369 = io_op_bits_active_vamo ? _GEN_19921 : _GEN_18143; // @[sequencer-master.scala 650:39]
  wire  _GEN_21370 = io_op_bits_active_vamo ? _GEN_19922 : _GEN_18144; // @[sequencer-master.scala 650:39]
  wire  _GEN_21371 = io_op_bits_active_vamo ? _GEN_19923 : _GEN_18145; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21372 = io_op_bits_active_vamo ? _GEN_19924 : _GEN_18146; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21373 = io_op_bits_active_vamo ? _GEN_19925 : _GEN_18147; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21374 = io_op_bits_active_vamo ? _GEN_19926 : _GEN_18148; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21375 = io_op_bits_active_vamo ? _GEN_19927 : _GEN_18149; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21376 = io_op_bits_active_vamo ? _GEN_19928 : _GEN_18150; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21377 = io_op_bits_active_vamo ? _GEN_19929 : _GEN_18151; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21378 = io_op_bits_active_vamo ? _GEN_19930 : _GEN_18152; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21379 = io_op_bits_active_vamo ? _GEN_19931 : _GEN_18153; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21380 = io_op_bits_active_vamo ? _GEN_20124 : _GEN_18154; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21381 = io_op_bits_active_vamo ? _GEN_20125 : _GEN_18155; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21382 = io_op_bits_active_vamo ? _GEN_20126 : _GEN_18156; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21383 = io_op_bits_active_vamo ? _GEN_20127 : _GEN_18157; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21384 = io_op_bits_active_vamo ? _GEN_20128 : _GEN_18158; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21385 = io_op_bits_active_vamo ? _GEN_20129 : _GEN_18159; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21386 = io_op_bits_active_vamo ? _GEN_20130 : _GEN_18160; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21387 = io_op_bits_active_vamo ? _GEN_20131 : _GEN_18161; // @[sequencer-master.scala 650:39]
  wire  _GEN_21388 = io_op_bits_active_vamo ? _GEN_20140 : _GEN_18162; // @[sequencer-master.scala 650:39]
  wire  _GEN_21389 = io_op_bits_active_vamo ? _GEN_20141 : _GEN_18163; // @[sequencer-master.scala 650:39]
  wire  _GEN_21390 = io_op_bits_active_vamo ? _GEN_20142 : _GEN_18164; // @[sequencer-master.scala 650:39]
  wire  _GEN_21391 = io_op_bits_active_vamo ? _GEN_20143 : _GEN_18165; // @[sequencer-master.scala 650:39]
  wire  _GEN_21392 = io_op_bits_active_vamo ? _GEN_20144 : _GEN_18166; // @[sequencer-master.scala 650:39]
  wire  _GEN_21393 = io_op_bits_active_vamo ? _GEN_20145 : _GEN_18167; // @[sequencer-master.scala 650:39]
  wire  _GEN_21394 = io_op_bits_active_vamo ? _GEN_20146 : _GEN_18168; // @[sequencer-master.scala 650:39]
  wire  _GEN_21395 = io_op_bits_active_vamo ? _GEN_20147 : _GEN_18169; // @[sequencer-master.scala 650:39]
  wire  _GEN_21396 = io_op_bits_active_vamo ? _GEN_20148 : _GEN_18170; // @[sequencer-master.scala 650:39]
  wire  _GEN_21397 = io_op_bits_active_vamo ? _GEN_20149 : _GEN_18171; // @[sequencer-master.scala 650:39]
  wire  _GEN_21398 = io_op_bits_active_vamo ? _GEN_20150 : _GEN_18172; // @[sequencer-master.scala 650:39]
  wire  _GEN_21399 = io_op_bits_active_vamo ? _GEN_20151 : _GEN_18173; // @[sequencer-master.scala 650:39]
  wire  _GEN_21400 = io_op_bits_active_vamo ? _GEN_20152 : _GEN_18174; // @[sequencer-master.scala 650:39]
  wire  _GEN_21401 = io_op_bits_active_vamo ? _GEN_20153 : _GEN_18175; // @[sequencer-master.scala 650:39]
  wire  _GEN_21402 = io_op_bits_active_vamo ? _GEN_20154 : _GEN_18176; // @[sequencer-master.scala 650:39]
  wire  _GEN_21403 = io_op_bits_active_vamo ? _GEN_20155 : _GEN_18177; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21404 = io_op_bits_active_vamo ? _GEN_20156 : _GEN_18178; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21405 = io_op_bits_active_vamo ? _GEN_20157 : _GEN_18179; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21406 = io_op_bits_active_vamo ? _GEN_20158 : _GEN_18180; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21407 = io_op_bits_active_vamo ? _GEN_20159 : _GEN_18181; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21408 = io_op_bits_active_vamo ? _GEN_20160 : _GEN_18182; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21409 = io_op_bits_active_vamo ? _GEN_20161 : _GEN_18183; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21410 = io_op_bits_active_vamo ? _GEN_20162 : _GEN_18184; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21411 = io_op_bits_active_vamo ? _GEN_20163 : _GEN_18185; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21412 = io_op_bits_active_vamo ? _GEN_20164 : _GEN_18186; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21413 = io_op_bits_active_vamo ? _GEN_20165 : _GEN_18187; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21414 = io_op_bits_active_vamo ? _GEN_20166 : _GEN_18188; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21415 = io_op_bits_active_vamo ? _GEN_20167 : _GEN_18189; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21416 = io_op_bits_active_vamo ? _GEN_20168 : _GEN_18190; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21417 = io_op_bits_active_vamo ? _GEN_20169 : _GEN_18191; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21418 = io_op_bits_active_vamo ? _GEN_20170 : _GEN_18192; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21419 = io_op_bits_active_vamo ? _GEN_20171 : _GEN_18193; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21420 = io_op_bits_active_vamo ? _GEN_20172 : _GEN_18194; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21421 = io_op_bits_active_vamo ? _GEN_20173 : _GEN_18195; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21422 = io_op_bits_active_vamo ? _GEN_20174 : _GEN_18196; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21423 = io_op_bits_active_vamo ? _GEN_20175 : _GEN_18197; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21424 = io_op_bits_active_vamo ? _GEN_20176 : _GEN_18198; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21425 = io_op_bits_active_vamo ? _GEN_20177 : _GEN_18199; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21426 = io_op_bits_active_vamo ? _GEN_20178 : _GEN_18200; // @[sequencer-master.scala 650:39]
  wire [63:0] _GEN_21427 = io_op_bits_active_vamo ? _GEN_20179 : _GEN_18201; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21428 = io_op_bits_active_vamo ? _GEN_21036 : _GEN_18202; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21429 = io_op_bits_active_vamo ? _GEN_21037 : _GEN_18203; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21430 = io_op_bits_active_vamo ? _GEN_21038 : _GEN_18204; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21431 = io_op_bits_active_vamo ? _GEN_21039 : _GEN_18205; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21432 = io_op_bits_active_vamo ? _GEN_21040 : _GEN_18206; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21433 = io_op_bits_active_vamo ? _GEN_21041 : _GEN_18207; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21434 = io_op_bits_active_vamo ? _GEN_21042 : _GEN_18208; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21435 = io_op_bits_active_vamo ? _GEN_21043 : _GEN_18209; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21436 = io_op_bits_active_vamo ? _GEN_21044 : _GEN_18210; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21437 = io_op_bits_active_vamo ? _GEN_21045 : _GEN_18211; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21438 = io_op_bits_active_vamo ? _GEN_21046 : _GEN_18212; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21439 = io_op_bits_active_vamo ? _GEN_21047 : _GEN_18213; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21440 = io_op_bits_active_vamo ? _GEN_21048 : _GEN_18214; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21441 = io_op_bits_active_vamo ? _GEN_21049 : _GEN_18215; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21442 = io_op_bits_active_vamo ? _GEN_21050 : _GEN_18216; // @[sequencer-master.scala 650:39]
  wire [3:0] _GEN_21443 = io_op_bits_active_vamo ? _GEN_21051 : _GEN_18217; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21444 = io_op_bits_active_vamo ? _GEN_21052 : _GEN_18218; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21445 = io_op_bits_active_vamo ? _GEN_21053 : _GEN_18219; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21446 = io_op_bits_active_vamo ? _GEN_21054 : _GEN_18220; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21447 = io_op_bits_active_vamo ? _GEN_21055 : _GEN_18221; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21448 = io_op_bits_active_vamo ? _GEN_21056 : _GEN_18222; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21449 = io_op_bits_active_vamo ? _GEN_21057 : _GEN_18223; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21450 = io_op_bits_active_vamo ? _GEN_21058 : _GEN_18224; // @[sequencer-master.scala 650:39]
  wire [2:0] _GEN_21451 = io_op_bits_active_vamo ? _GEN_21059 : _GEN_18225; // @[sequencer-master.scala 650:39]
  wire  _GEN_21452 = io_op_bits_active_vamo ? _GEN_19268 : e_0_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21453 = io_op_bits_active_vamo ? _GEN_19269 : e_1_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21454 = io_op_bits_active_vamo ? _GEN_19270 : e_2_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21455 = io_op_bits_active_vamo ? _GEN_19271 : e_3_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21456 = io_op_bits_active_vamo ? _GEN_19272 : e_4_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21457 = io_op_bits_active_vamo ? _GEN_19273 : e_5_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21458 = io_op_bits_active_vamo ? _GEN_19274 : e_6_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21459 = io_op_bits_active_vamo ? _GEN_19275 : e_7_active_vcu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21460 = io_op_bits_active_vamo ? _GEN_19836 : e_0_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21461 = io_op_bits_active_vamo ? _GEN_19837 : e_1_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21462 = io_op_bits_active_vamo ? _GEN_19838 : e_2_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21463 = io_op_bits_active_vamo ? _GEN_19839 : e_3_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21464 = io_op_bits_active_vamo ? _GEN_19840 : e_4_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21465 = io_op_bits_active_vamo ? _GEN_19841 : e_5_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21466 = io_op_bits_active_vamo ? _GEN_19842 : e_6_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21467 = io_op_bits_active_vamo ? _GEN_19843 : e_7_active_vsu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21468 = io_op_bits_active_vamo ? _GEN_20668 : e_0_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21469 = io_op_bits_active_vamo ? _GEN_20669 : e_1_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21470 = io_op_bits_active_vamo ? _GEN_20670 : e_2_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21471 = io_op_bits_active_vamo ? _GEN_20671 : e_3_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21472 = io_op_bits_active_vamo ? _GEN_20672 : e_4_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21473 = io_op_bits_active_vamo ? _GEN_20673 : e_5_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21474 = io_op_bits_active_vamo ? _GEN_20674 : e_6_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire  _GEN_21475 = io_op_bits_active_vamo ? _GEN_20675 : e_7_active_vlu; // @[sequencer-master.scala 650:39 sequencer-master.scala 109:14]
  wire [7:0] _GEN_21476 = io_op_bits_active_vamo ? _GEN_20732 : _GEN_16134; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21477 = io_op_bits_active_vamo ? _GEN_20733 : _GEN_16135; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21478 = io_op_bits_active_vamo ? _GEN_20734 : _GEN_16136; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21479 = io_op_bits_active_vamo ? _GEN_20735 : _GEN_16137; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21480 = io_op_bits_active_vamo ? _GEN_20736 : _GEN_16138; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21481 = io_op_bits_active_vamo ? _GEN_20737 : _GEN_16139; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21482 = io_op_bits_active_vamo ? _GEN_20738 : _GEN_16140; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21483 = io_op_bits_active_vamo ? _GEN_20739 : _GEN_16141; // @[sequencer-master.scala 650:39]
  wire  _GEN_21484 = io_op_bits_active_vamo ? _GEN_20748 : _GEN_16142; // @[sequencer-master.scala 650:39]
  wire  _GEN_21485 = io_op_bits_active_vamo ? _GEN_20749 : _GEN_16143; // @[sequencer-master.scala 650:39]
  wire  _GEN_21486 = io_op_bits_active_vamo ? _GEN_20750 : _GEN_16144; // @[sequencer-master.scala 650:39]
  wire  _GEN_21487 = io_op_bits_active_vamo ? _GEN_20751 : _GEN_16145; // @[sequencer-master.scala 650:39]
  wire  _GEN_21488 = io_op_bits_active_vamo ? _GEN_20752 : _GEN_16146; // @[sequencer-master.scala 650:39]
  wire  _GEN_21489 = io_op_bits_active_vamo ? _GEN_20753 : _GEN_16147; // @[sequencer-master.scala 650:39]
  wire  _GEN_21490 = io_op_bits_active_vamo ? _GEN_20754 : _GEN_16148; // @[sequencer-master.scala 650:39]
  wire  _GEN_21491 = io_op_bits_active_vamo ? _GEN_20755 : _GEN_16149; // @[sequencer-master.scala 650:39]
  wire  _GEN_21492 = io_op_bits_active_vamo ? _GEN_20756 : _GEN_16150; // @[sequencer-master.scala 650:39]
  wire  _GEN_21493 = io_op_bits_active_vamo ? _GEN_20757 : _GEN_16151; // @[sequencer-master.scala 650:39]
  wire  _GEN_21494 = io_op_bits_active_vamo ? _GEN_20758 : _GEN_16152; // @[sequencer-master.scala 650:39]
  wire  _GEN_21495 = io_op_bits_active_vamo ? _GEN_20759 : _GEN_16153; // @[sequencer-master.scala 650:39]
  wire  _GEN_21496 = io_op_bits_active_vamo ? _GEN_20760 : _GEN_16154; // @[sequencer-master.scala 650:39]
  wire  _GEN_21497 = io_op_bits_active_vamo ? _GEN_20761 : _GEN_16155; // @[sequencer-master.scala 650:39]
  wire  _GEN_21498 = io_op_bits_active_vamo ? _GEN_20762 : _GEN_16156; // @[sequencer-master.scala 650:39]
  wire  _GEN_21499 = io_op_bits_active_vamo ? _GEN_20763 : _GEN_16157; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21500 = io_op_bits_active_vamo ? _GEN_20764 : _GEN_16158; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21501 = io_op_bits_active_vamo ? _GEN_20765 : _GEN_16159; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21502 = io_op_bits_active_vamo ? _GEN_20766 : _GEN_16160; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21503 = io_op_bits_active_vamo ? _GEN_20767 : _GEN_16161; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21504 = io_op_bits_active_vamo ? _GEN_20768 : _GEN_16162; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21505 = io_op_bits_active_vamo ? _GEN_20769 : _GEN_16163; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21506 = io_op_bits_active_vamo ? _GEN_20770 : _GEN_16164; // @[sequencer-master.scala 650:39]
  wire [1:0] _GEN_21507 = io_op_bits_active_vamo ? _GEN_20771 : _GEN_16165; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21508 = io_op_bits_active_vamo ? _GEN_20772 : _GEN_16166; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21509 = io_op_bits_active_vamo ? _GEN_20773 : _GEN_16167; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21510 = io_op_bits_active_vamo ? _GEN_20774 : _GEN_16168; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21511 = io_op_bits_active_vamo ? _GEN_20775 : _GEN_16169; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21512 = io_op_bits_active_vamo ? _GEN_20776 : _GEN_16170; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21513 = io_op_bits_active_vamo ? _GEN_20777 : _GEN_16171; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21514 = io_op_bits_active_vamo ? _GEN_20778 : _GEN_16172; // @[sequencer-master.scala 650:39]
  wire [7:0] _GEN_21515 = io_op_bits_active_vamo ? _GEN_20779 : _GEN_16173; // @[sequencer-master.scala 650:39]
  wire  _GEN_21516 = io_op_bits_active_vamo | _GEN_18226; // @[sequencer-master.scala 650:39 sequencer-master.scala 265:41]
  wire [2:0] _GEN_21517 = io_op_bits_active_vamo ? _T_1651 : _GEN_18227; // @[sequencer-master.scala 650:39 sequencer-master.scala 265:66]
  wire  _GEN_21534 = 3'h0 == tail ? 1'h0 : _GEN_21076; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21535 = 3'h1 == tail ? 1'h0 : _GEN_21077; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21536 = 3'h2 == tail ? 1'h0 : _GEN_21078; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21537 = 3'h3 == tail ? 1'h0 : _GEN_21079; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21538 = 3'h4 == tail ? 1'h0 : _GEN_21080; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21539 = 3'h5 == tail ? 1'h0 : _GEN_21081; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21540 = 3'h6 == tail ? 1'h0 : _GEN_21082; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21541 = 3'h7 == tail ? 1'h0 : _GEN_21083; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_21542 = 3'h0 == tail ? 1'h0 : _GEN_21084; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21543 = 3'h1 == tail ? 1'h0 : _GEN_21085; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21544 = 3'h2 == tail ? 1'h0 : _GEN_21086; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21545 = 3'h3 == tail ? 1'h0 : _GEN_21087; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21546 = 3'h4 == tail ? 1'h0 : _GEN_21088; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21547 = 3'h5 == tail ? 1'h0 : _GEN_21089; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21548 = 3'h6 == tail ? 1'h0 : _GEN_21090; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21549 = 3'h7 == tail ? 1'h0 : _GEN_21091; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_21550 = 3'h0 == tail ? 1'h0 : _GEN_21092; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21551 = 3'h1 == tail ? 1'h0 : _GEN_21093; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21552 = 3'h2 == tail ? 1'h0 : _GEN_21094; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21553 = 3'h3 == tail ? 1'h0 : _GEN_21095; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21554 = 3'h4 == tail ? 1'h0 : _GEN_21096; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21555 = 3'h5 == tail ? 1'h0 : _GEN_21097; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21556 = 3'h6 == tail ? 1'h0 : _GEN_21098; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21557 = 3'h7 == tail ? 1'h0 : _GEN_21099; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_21558 = 3'h0 == tail ? 1'h0 : _GEN_21100; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21559 = 3'h1 == tail ? 1'h0 : _GEN_21101; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21560 = 3'h2 == tail ? 1'h0 : _GEN_21102; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21561 = 3'h3 == tail ? 1'h0 : _GEN_21103; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21562 = 3'h4 == tail ? 1'h0 : _GEN_21104; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21563 = 3'h5 == tail ? 1'h0 : _GEN_21105; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21564 = 3'h6 == tail ? 1'h0 : _GEN_21106; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21565 = 3'h7 == tail ? 1'h0 : _GEN_21107; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_21566 = 3'h0 == tail ? 1'h0 : _GEN_21108; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21567 = 3'h1 == tail ? 1'h0 : _GEN_21109; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21568 = 3'h2 == tail ? 1'h0 : _GEN_21110; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21569 = 3'h3 == tail ? 1'h0 : _GEN_21111; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21570 = 3'h4 == tail ? 1'h0 : _GEN_21112; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21571 = 3'h5 == tail ? 1'h0 : _GEN_21113; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21572 = 3'h6 == tail ? 1'h0 : _GEN_21114; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21573 = 3'h7 == tail ? 1'h0 : _GEN_21115; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_21582 = 3'h0 == tail ? 1'h0 : _GEN_21124; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21583 = 3'h1 == tail ? 1'h0 : _GEN_21125; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21584 = 3'h2 == tail ? 1'h0 : _GEN_21126; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21585 = 3'h3 == tail ? 1'h0 : _GEN_21127; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21586 = 3'h4 == tail ? 1'h0 : _GEN_21128; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21587 = 3'h5 == tail ? 1'h0 : _GEN_21129; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21588 = 3'h6 == tail ? 1'h0 : _GEN_21130; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21589 = 3'h7 == tail ? 1'h0 : _GEN_21131; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21590 = 3'h0 == tail ? 1'h0 : _GEN_21132; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21591 = 3'h1 == tail ? 1'h0 : _GEN_21133; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21592 = 3'h2 == tail ? 1'h0 : _GEN_21134; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21593 = 3'h3 == tail ? 1'h0 : _GEN_21135; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21594 = 3'h4 == tail ? 1'h0 : _GEN_21136; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21595 = 3'h5 == tail ? 1'h0 : _GEN_21137; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21596 = 3'h6 == tail ? 1'h0 : _GEN_21138; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21597 = 3'h7 == tail ? 1'h0 : _GEN_21139; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21598 = 3'h0 == tail ? 1'h0 : _GEN_21140; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21599 = 3'h1 == tail ? 1'h0 : _GEN_21141; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21600 = 3'h2 == tail ? 1'h0 : _GEN_21142; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21601 = 3'h3 == tail ? 1'h0 : _GEN_21143; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21602 = 3'h4 == tail ? 1'h0 : _GEN_21144; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21603 = 3'h5 == tail ? 1'h0 : _GEN_21145; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21604 = 3'h6 == tail ? 1'h0 : _GEN_21146; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21605 = 3'h7 == tail ? 1'h0 : _GEN_21147; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21606 = 3'h0 == tail ? 1'h0 : _GEN_21148; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21607 = 3'h1 == tail ? 1'h0 : _GEN_21149; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21608 = 3'h2 == tail ? 1'h0 : _GEN_21150; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21609 = 3'h3 == tail ? 1'h0 : _GEN_21151; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21610 = 3'h4 == tail ? 1'h0 : _GEN_21152; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21611 = 3'h5 == tail ? 1'h0 : _GEN_21153; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21612 = 3'h6 == tail ? 1'h0 : _GEN_21154; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21613 = 3'h7 == tail ? 1'h0 : _GEN_21155; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21614 = 3'h0 == tail ? 1'h0 : _GEN_21156; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21615 = 3'h1 == tail ? 1'h0 : _GEN_21157; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21616 = 3'h2 == tail ? 1'h0 : _GEN_21158; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21617 = 3'h3 == tail ? 1'h0 : _GEN_21159; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21618 = 3'h4 == tail ? 1'h0 : _GEN_21160; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21619 = 3'h5 == tail ? 1'h0 : _GEN_21161; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21620 = 3'h6 == tail ? 1'h0 : _GEN_21162; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21621 = 3'h7 == tail ? 1'h0 : _GEN_21163; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21622 = 3'h0 == tail ? 1'h0 : _GEN_21164; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21623 = 3'h1 == tail ? 1'h0 : _GEN_21165; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21624 = 3'h2 == tail ? 1'h0 : _GEN_21166; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21625 = 3'h3 == tail ? 1'h0 : _GEN_21167; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21626 = 3'h4 == tail ? 1'h0 : _GEN_21168; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21627 = 3'h5 == tail ? 1'h0 : _GEN_21169; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21628 = 3'h6 == tail ? 1'h0 : _GEN_21170; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21629 = 3'h7 == tail ? 1'h0 : _GEN_21171; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21630 = 3'h0 == tail ? 1'h0 : _GEN_21172; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21631 = 3'h1 == tail ? 1'h0 : _GEN_21173; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21632 = 3'h2 == tail ? 1'h0 : _GEN_21174; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21633 = 3'h3 == tail ? 1'h0 : _GEN_21175; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21634 = 3'h4 == tail ? 1'h0 : _GEN_21176; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21635 = 3'h5 == tail ? 1'h0 : _GEN_21177; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21636 = 3'h6 == tail ? 1'h0 : _GEN_21178; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21637 = 3'h7 == tail ? 1'h0 : _GEN_21179; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21638 = 3'h0 == tail ? 1'h0 : _GEN_21180; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21639 = 3'h1 == tail ? 1'h0 : _GEN_21181; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21640 = 3'h2 == tail ? 1'h0 : _GEN_21182; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21641 = 3'h3 == tail ? 1'h0 : _GEN_21183; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21642 = 3'h4 == tail ? 1'h0 : _GEN_21184; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21643 = 3'h5 == tail ? 1'h0 : _GEN_21185; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21644 = 3'h6 == tail ? 1'h0 : _GEN_21186; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21645 = 3'h7 == tail ? 1'h0 : _GEN_21187; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21646 = 3'h0 == tail ? 1'h0 : _GEN_21188; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21647 = 3'h1 == tail ? 1'h0 : _GEN_21189; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21648 = 3'h2 == tail ? 1'h0 : _GEN_21190; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21649 = 3'h3 == tail ? 1'h0 : _GEN_21191; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21650 = 3'h4 == tail ? 1'h0 : _GEN_21192; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21651 = 3'h5 == tail ? 1'h0 : _GEN_21193; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21652 = 3'h6 == tail ? 1'h0 : _GEN_21194; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21653 = 3'h7 == tail ? 1'h0 : _GEN_21195; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21654 = 3'h0 == tail ? 1'h0 : _GEN_21196; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21655 = 3'h1 == tail ? 1'h0 : _GEN_21197; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21656 = 3'h2 == tail ? 1'h0 : _GEN_21198; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21657 = 3'h3 == tail ? 1'h0 : _GEN_21199; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21658 = 3'h4 == tail ? 1'h0 : _GEN_21200; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21659 = 3'h5 == tail ? 1'h0 : _GEN_21201; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21660 = 3'h6 == tail ? 1'h0 : _GEN_21202; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21661 = 3'h7 == tail ? 1'h0 : _GEN_21203; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21662 = 3'h0 == tail ? 1'h0 : _GEN_21204; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21663 = 3'h1 == tail ? 1'h0 : _GEN_21205; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21664 = 3'h2 == tail ? 1'h0 : _GEN_21206; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21665 = 3'h3 == tail ? 1'h0 : _GEN_21207; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21666 = 3'h4 == tail ? 1'h0 : _GEN_21208; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21667 = 3'h5 == tail ? 1'h0 : _GEN_21209; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21668 = 3'h6 == tail ? 1'h0 : _GEN_21210; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21669 = 3'h7 == tail ? 1'h0 : _GEN_21211; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21670 = 3'h0 == tail ? 1'h0 : _GEN_21212; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21671 = 3'h1 == tail ? 1'h0 : _GEN_21213; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21672 = 3'h2 == tail ? 1'h0 : _GEN_21214; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21673 = 3'h3 == tail ? 1'h0 : _GEN_21215; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21674 = 3'h4 == tail ? 1'h0 : _GEN_21216; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21675 = 3'h5 == tail ? 1'h0 : _GEN_21217; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21676 = 3'h6 == tail ? 1'h0 : _GEN_21218; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21677 = 3'h7 == tail ? 1'h0 : _GEN_21219; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21678 = 3'h0 == tail ? 1'h0 : _GEN_21220; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21679 = 3'h1 == tail ? 1'h0 : _GEN_21221; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21680 = 3'h2 == tail ? 1'h0 : _GEN_21222; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21681 = 3'h3 == tail ? 1'h0 : _GEN_21223; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21682 = 3'h4 == tail ? 1'h0 : _GEN_21224; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21683 = 3'h5 == tail ? 1'h0 : _GEN_21225; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21684 = 3'h6 == tail ? 1'h0 : _GEN_21226; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21685 = 3'h7 == tail ? 1'h0 : _GEN_21227; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21686 = 3'h0 == tail ? 1'h0 : _GEN_21228; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21687 = 3'h1 == tail ? 1'h0 : _GEN_21229; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21688 = 3'h2 == tail ? 1'h0 : _GEN_21230; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21689 = 3'h3 == tail ? 1'h0 : _GEN_21231; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21690 = 3'h4 == tail ? 1'h0 : _GEN_21232; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21691 = 3'h5 == tail ? 1'h0 : _GEN_21233; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21692 = 3'h6 == tail ? 1'h0 : _GEN_21234; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21693 = 3'h7 == tail ? 1'h0 : _GEN_21235; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21694 = 3'h0 == tail ? 1'h0 : _GEN_21236; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21695 = 3'h1 == tail ? 1'h0 : _GEN_21237; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21696 = 3'h2 == tail ? 1'h0 : _GEN_21238; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21697 = 3'h3 == tail ? 1'h0 : _GEN_21239; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21698 = 3'h4 == tail ? 1'h0 : _GEN_21240; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21699 = 3'h5 == tail ? 1'h0 : _GEN_21241; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21700 = 3'h6 == tail ? 1'h0 : _GEN_21242; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21701 = 3'h7 == tail ? 1'h0 : _GEN_21243; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21702 = 3'h0 == tail ? 1'h0 : _GEN_21244; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21703 = 3'h1 == tail ? 1'h0 : _GEN_21245; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21704 = 3'h2 == tail ? 1'h0 : _GEN_21246; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21705 = 3'h3 == tail ? 1'h0 : _GEN_21247; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21706 = 3'h4 == tail ? 1'h0 : _GEN_21248; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21707 = 3'h5 == tail ? 1'h0 : _GEN_21249; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21708 = 3'h6 == tail ? 1'h0 : _GEN_21250; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21709 = 3'h7 == tail ? 1'h0 : _GEN_21251; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21710 = 3'h0 == tail ? 1'h0 : _GEN_21252; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21711 = 3'h1 == tail ? 1'h0 : _GEN_21253; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21712 = 3'h2 == tail ? 1'h0 : _GEN_21254; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21713 = 3'h3 == tail ? 1'h0 : _GEN_21255; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21714 = 3'h4 == tail ? 1'h0 : _GEN_21256; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21715 = 3'h5 == tail ? 1'h0 : _GEN_21257; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21716 = 3'h6 == tail ? 1'h0 : _GEN_21258; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21717 = 3'h7 == tail ? 1'h0 : _GEN_21259; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21718 = 3'h0 == tail ? 1'h0 : _GEN_21260; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21719 = 3'h1 == tail ? 1'h0 : _GEN_21261; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21720 = 3'h2 == tail ? 1'h0 : _GEN_21262; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21721 = 3'h3 == tail ? 1'h0 : _GEN_21263; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21722 = 3'h4 == tail ? 1'h0 : _GEN_21264; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21723 = 3'h5 == tail ? 1'h0 : _GEN_21265; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21724 = 3'h6 == tail ? 1'h0 : _GEN_21266; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21725 = 3'h7 == tail ? 1'h0 : _GEN_21267; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21726 = 3'h0 == tail ? 1'h0 : _GEN_21268; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21727 = 3'h1 == tail ? 1'h0 : _GEN_21269; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21728 = 3'h2 == tail ? 1'h0 : _GEN_21270; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21729 = 3'h3 == tail ? 1'h0 : _GEN_21271; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21730 = 3'h4 == tail ? 1'h0 : _GEN_21272; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21731 = 3'h5 == tail ? 1'h0 : _GEN_21273; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21732 = 3'h6 == tail ? 1'h0 : _GEN_21274; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21733 = 3'h7 == tail ? 1'h0 : _GEN_21275; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21734 = 3'h0 == tail ? 1'h0 : _GEN_21276; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21735 = 3'h1 == tail ? 1'h0 : _GEN_21277; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21736 = 3'h2 == tail ? 1'h0 : _GEN_21278; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21737 = 3'h3 == tail ? 1'h0 : _GEN_21279; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21738 = 3'h4 == tail ? 1'h0 : _GEN_21280; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21739 = 3'h5 == tail ? 1'h0 : _GEN_21281; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21740 = 3'h6 == tail ? 1'h0 : _GEN_21282; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21741 = 3'h7 == tail ? 1'h0 : _GEN_21283; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21742 = 3'h0 == tail ? 1'h0 : _GEN_21284; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21743 = 3'h1 == tail ? 1'h0 : _GEN_21285; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21744 = 3'h2 == tail ? 1'h0 : _GEN_21286; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21745 = 3'h3 == tail ? 1'h0 : _GEN_21287; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21746 = 3'h4 == tail ? 1'h0 : _GEN_21288; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21747 = 3'h5 == tail ? 1'h0 : _GEN_21289; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21748 = 3'h6 == tail ? 1'h0 : _GEN_21290; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21749 = 3'h7 == tail ? 1'h0 : _GEN_21291; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21750 = 3'h0 == tail ? 1'h0 : _GEN_21292; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21751 = 3'h1 == tail ? 1'h0 : _GEN_21293; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21752 = 3'h2 == tail ? 1'h0 : _GEN_21294; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21753 = 3'h3 == tail ? 1'h0 : _GEN_21295; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21754 = 3'h4 == tail ? 1'h0 : _GEN_21296; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21755 = 3'h5 == tail ? 1'h0 : _GEN_21297; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21756 = 3'h6 == tail ? 1'h0 : _GEN_21298; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21757 = 3'h7 == tail ? 1'h0 : _GEN_21299; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_21758 = 3'h0 == tail ? 1'h0 : _GEN_21300; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21759 = 3'h1 == tail ? 1'h0 : _GEN_21301; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21760 = 3'h2 == tail ? 1'h0 : _GEN_21302; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21761 = 3'h3 == tail ? 1'h0 : _GEN_21303; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21762 = 3'h4 == tail ? 1'h0 : _GEN_21304; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21763 = 3'h5 == tail ? 1'h0 : _GEN_21305; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21764 = 3'h6 == tail ? 1'h0 : _GEN_21306; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21765 = 3'h7 == tail ? 1'h0 : _GEN_21307; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_21766 = 3'h0 == tail ? 1'h0 : _GEN_21308; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21767 = 3'h1 == tail ? 1'h0 : _GEN_21309; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21768 = 3'h2 == tail ? 1'h0 : _GEN_21310; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21769 = 3'h3 == tail ? 1'h0 : _GEN_21311; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21770 = 3'h4 == tail ? 1'h0 : _GEN_21312; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21771 = 3'h5 == tail ? 1'h0 : _GEN_21313; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21772 = 3'h6 == tail ? 1'h0 : _GEN_21314; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21773 = 3'h7 == tail ? 1'h0 : _GEN_21315; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_21774 = 3'h0 == tail ? 1'h0 : _GEN_21316; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21775 = 3'h1 == tail ? 1'h0 : _GEN_21317; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21776 = 3'h2 == tail ? 1'h0 : _GEN_21318; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21777 = 3'h3 == tail ? 1'h0 : _GEN_21319; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21778 = 3'h4 == tail ? 1'h0 : _GEN_21320; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21779 = 3'h5 == tail ? 1'h0 : _GEN_21321; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21780 = 3'h6 == tail ? 1'h0 : _GEN_21322; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21781 = 3'h7 == tail ? 1'h0 : _GEN_21323; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_21790 = _GEN_32729 | _GEN_21332; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21791 = _GEN_32730 | _GEN_21333; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21792 = _GEN_32731 | _GEN_21334; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21793 = _GEN_32732 | _GEN_21335; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21794 = _GEN_32733 | _GEN_21336; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21795 = _GEN_32734 | _GEN_21337; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21796 = _GEN_32735 | _GEN_21338; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_21797 = _GEN_32736 | _GEN_21339; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_21798 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_21340; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21799 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_21341; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21800 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_21342; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21801 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_21343; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21802 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_21344; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21803 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_21345; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21804 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_21346; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_21805 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_21347; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_21806 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_21348; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21807 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_21349; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21808 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_21350; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21809 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_21351; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21810 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_21352; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21811 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_21353; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21812 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_21354; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_21813 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_21355; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21814 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_21534; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21815 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_21535; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21816 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_21536; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21817 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_21537; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21818 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_21538; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21819 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_21539; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21820 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_21540; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21821 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_21541; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21822 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_21356; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21823 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_21357; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21824 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_21358; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21825 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_21359; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21826 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_21360; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21827 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_21361; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21828 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_21362; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21829 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_21363; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21830 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_21364; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21831 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_21365; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21832 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_21366; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21833 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_21367; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21834 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_21368; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21835 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_21369; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21836 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_21370; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_21837 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_21371; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_21838 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_21372; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21839 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_21373; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21840 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_21374; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21841 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_21375; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21842 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_21376; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21843 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_21377; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21844 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_21378; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_21845 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_21379; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_21846 = io_op_bits_base_vp_valid ? _GEN_21806 : _GEN_21348; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21847 = io_op_bits_base_vp_valid ? _GEN_21807 : _GEN_21349; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21848 = io_op_bits_base_vp_valid ? _GEN_21808 : _GEN_21350; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21849 = io_op_bits_base_vp_valid ? _GEN_21809 : _GEN_21351; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21850 = io_op_bits_base_vp_valid ? _GEN_21810 : _GEN_21352; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21851 = io_op_bits_base_vp_valid ? _GEN_21811 : _GEN_21353; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21852 = io_op_bits_base_vp_valid ? _GEN_21812 : _GEN_21354; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_21853 = io_op_bits_base_vp_valid ? _GEN_21813 : _GEN_21355; // @[sequencer-master.scala 320:41]
  wire  _GEN_21854 = io_op_bits_base_vp_valid ? _GEN_21814 : _GEN_21534; // @[sequencer-master.scala 320:41]
  wire  _GEN_21855 = io_op_bits_base_vp_valid ? _GEN_21815 : _GEN_21535; // @[sequencer-master.scala 320:41]
  wire  _GEN_21856 = io_op_bits_base_vp_valid ? _GEN_21816 : _GEN_21536; // @[sequencer-master.scala 320:41]
  wire  _GEN_21857 = io_op_bits_base_vp_valid ? _GEN_21817 : _GEN_21537; // @[sequencer-master.scala 320:41]
  wire  _GEN_21858 = io_op_bits_base_vp_valid ? _GEN_21818 : _GEN_21538; // @[sequencer-master.scala 320:41]
  wire  _GEN_21859 = io_op_bits_base_vp_valid ? _GEN_21819 : _GEN_21539; // @[sequencer-master.scala 320:41]
  wire  _GEN_21860 = io_op_bits_base_vp_valid ? _GEN_21820 : _GEN_21540; // @[sequencer-master.scala 320:41]
  wire  _GEN_21861 = io_op_bits_base_vp_valid ? _GEN_21821 : _GEN_21541; // @[sequencer-master.scala 320:41]
  wire  _GEN_21862 = io_op_bits_base_vp_valid ? _GEN_21822 : _GEN_21356; // @[sequencer-master.scala 320:41]
  wire  _GEN_21863 = io_op_bits_base_vp_valid ? _GEN_21823 : _GEN_21357; // @[sequencer-master.scala 320:41]
  wire  _GEN_21864 = io_op_bits_base_vp_valid ? _GEN_21824 : _GEN_21358; // @[sequencer-master.scala 320:41]
  wire  _GEN_21865 = io_op_bits_base_vp_valid ? _GEN_21825 : _GEN_21359; // @[sequencer-master.scala 320:41]
  wire  _GEN_21866 = io_op_bits_base_vp_valid ? _GEN_21826 : _GEN_21360; // @[sequencer-master.scala 320:41]
  wire  _GEN_21867 = io_op_bits_base_vp_valid ? _GEN_21827 : _GEN_21361; // @[sequencer-master.scala 320:41]
  wire  _GEN_21868 = io_op_bits_base_vp_valid ? _GEN_21828 : _GEN_21362; // @[sequencer-master.scala 320:41]
  wire  _GEN_21869 = io_op_bits_base_vp_valid ? _GEN_21829 : _GEN_21363; // @[sequencer-master.scala 320:41]
  wire  _GEN_21870 = io_op_bits_base_vp_valid ? _GEN_21830 : _GEN_21364; // @[sequencer-master.scala 320:41]
  wire  _GEN_21871 = io_op_bits_base_vp_valid ? _GEN_21831 : _GEN_21365; // @[sequencer-master.scala 320:41]
  wire  _GEN_21872 = io_op_bits_base_vp_valid ? _GEN_21832 : _GEN_21366; // @[sequencer-master.scala 320:41]
  wire  _GEN_21873 = io_op_bits_base_vp_valid ? _GEN_21833 : _GEN_21367; // @[sequencer-master.scala 320:41]
  wire  _GEN_21874 = io_op_bits_base_vp_valid ? _GEN_21834 : _GEN_21368; // @[sequencer-master.scala 320:41]
  wire  _GEN_21875 = io_op_bits_base_vp_valid ? _GEN_21835 : _GEN_21369; // @[sequencer-master.scala 320:41]
  wire  _GEN_21876 = io_op_bits_base_vp_valid ? _GEN_21836 : _GEN_21370; // @[sequencer-master.scala 320:41]
  wire  _GEN_21877 = io_op_bits_base_vp_valid ? _GEN_21837 : _GEN_21371; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21878 = io_op_bits_base_vp_valid ? _GEN_21838 : _GEN_21372; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21879 = io_op_bits_base_vp_valid ? _GEN_21839 : _GEN_21373; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21880 = io_op_bits_base_vp_valid ? _GEN_21840 : _GEN_21374; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21881 = io_op_bits_base_vp_valid ? _GEN_21841 : _GEN_21375; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21882 = io_op_bits_base_vp_valid ? _GEN_21842 : _GEN_21376; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21883 = io_op_bits_base_vp_valid ? _GEN_21843 : _GEN_21377; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21884 = io_op_bits_base_vp_valid ? _GEN_21844 : _GEN_21378; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_21885 = io_op_bits_base_vp_valid ? _GEN_21845 : _GEN_21379; // @[sequencer-master.scala 320:41]
  wire  _GEN_21886 = _GEN_32729 | _GEN_21582; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21887 = _GEN_32730 | _GEN_21583; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21888 = _GEN_32731 | _GEN_21584; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21889 = _GEN_32732 | _GEN_21585; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21890 = _GEN_32733 | _GEN_21586; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21891 = _GEN_32734 | _GEN_21587; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21892 = _GEN_32735 | _GEN_21588; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21893 = _GEN_32736 | _GEN_21589; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21894 = _T_26 ? _GEN_21886 : _GEN_21582; // @[sequencer-master.scala 154:24]
  wire  _GEN_21895 = _T_26 ? _GEN_21887 : _GEN_21583; // @[sequencer-master.scala 154:24]
  wire  _GEN_21896 = _T_26 ? _GEN_21888 : _GEN_21584; // @[sequencer-master.scala 154:24]
  wire  _GEN_21897 = _T_26 ? _GEN_21889 : _GEN_21585; // @[sequencer-master.scala 154:24]
  wire  _GEN_21898 = _T_26 ? _GEN_21890 : _GEN_21586; // @[sequencer-master.scala 154:24]
  wire  _GEN_21899 = _T_26 ? _GEN_21891 : _GEN_21587; // @[sequencer-master.scala 154:24]
  wire  _GEN_21900 = _T_26 ? _GEN_21892 : _GEN_21588; // @[sequencer-master.scala 154:24]
  wire  _GEN_21901 = _T_26 ? _GEN_21893 : _GEN_21589; // @[sequencer-master.scala 154:24]
  wire  _GEN_21902 = _GEN_32729 | _GEN_21606; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21903 = _GEN_32730 | _GEN_21607; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21904 = _GEN_32731 | _GEN_21608; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21905 = _GEN_32732 | _GEN_21609; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21906 = _GEN_32733 | _GEN_21610; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21907 = _GEN_32734 | _GEN_21611; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21908 = _GEN_32735 | _GEN_21612; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21909 = _GEN_32736 | _GEN_21613; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21910 = _T_48 ? _GEN_21902 : _GEN_21606; // @[sequencer-master.scala 154:24]
  wire  _GEN_21911 = _T_48 ? _GEN_21903 : _GEN_21607; // @[sequencer-master.scala 154:24]
  wire  _GEN_21912 = _T_48 ? _GEN_21904 : _GEN_21608; // @[sequencer-master.scala 154:24]
  wire  _GEN_21913 = _T_48 ? _GEN_21905 : _GEN_21609; // @[sequencer-master.scala 154:24]
  wire  _GEN_21914 = _T_48 ? _GEN_21906 : _GEN_21610; // @[sequencer-master.scala 154:24]
  wire  _GEN_21915 = _T_48 ? _GEN_21907 : _GEN_21611; // @[sequencer-master.scala 154:24]
  wire  _GEN_21916 = _T_48 ? _GEN_21908 : _GEN_21612; // @[sequencer-master.scala 154:24]
  wire  _GEN_21917 = _T_48 ? _GEN_21909 : _GEN_21613; // @[sequencer-master.scala 154:24]
  wire  _GEN_21918 = _GEN_32729 | _GEN_21630; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21919 = _GEN_32730 | _GEN_21631; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21920 = _GEN_32731 | _GEN_21632; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21921 = _GEN_32732 | _GEN_21633; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21922 = _GEN_32733 | _GEN_21634; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21923 = _GEN_32734 | _GEN_21635; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21924 = _GEN_32735 | _GEN_21636; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21925 = _GEN_32736 | _GEN_21637; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21926 = _T_70 ? _GEN_21918 : _GEN_21630; // @[sequencer-master.scala 154:24]
  wire  _GEN_21927 = _T_70 ? _GEN_21919 : _GEN_21631; // @[sequencer-master.scala 154:24]
  wire  _GEN_21928 = _T_70 ? _GEN_21920 : _GEN_21632; // @[sequencer-master.scala 154:24]
  wire  _GEN_21929 = _T_70 ? _GEN_21921 : _GEN_21633; // @[sequencer-master.scala 154:24]
  wire  _GEN_21930 = _T_70 ? _GEN_21922 : _GEN_21634; // @[sequencer-master.scala 154:24]
  wire  _GEN_21931 = _T_70 ? _GEN_21923 : _GEN_21635; // @[sequencer-master.scala 154:24]
  wire  _GEN_21932 = _T_70 ? _GEN_21924 : _GEN_21636; // @[sequencer-master.scala 154:24]
  wire  _GEN_21933 = _T_70 ? _GEN_21925 : _GEN_21637; // @[sequencer-master.scala 154:24]
  wire  _GEN_21934 = _GEN_32729 | _GEN_21654; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21935 = _GEN_32730 | _GEN_21655; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21936 = _GEN_32731 | _GEN_21656; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21937 = _GEN_32732 | _GEN_21657; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21938 = _GEN_32733 | _GEN_21658; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21939 = _GEN_32734 | _GEN_21659; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21940 = _GEN_32735 | _GEN_21660; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21941 = _GEN_32736 | _GEN_21661; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21942 = _T_92 ? _GEN_21934 : _GEN_21654; // @[sequencer-master.scala 154:24]
  wire  _GEN_21943 = _T_92 ? _GEN_21935 : _GEN_21655; // @[sequencer-master.scala 154:24]
  wire  _GEN_21944 = _T_92 ? _GEN_21936 : _GEN_21656; // @[sequencer-master.scala 154:24]
  wire  _GEN_21945 = _T_92 ? _GEN_21937 : _GEN_21657; // @[sequencer-master.scala 154:24]
  wire  _GEN_21946 = _T_92 ? _GEN_21938 : _GEN_21658; // @[sequencer-master.scala 154:24]
  wire  _GEN_21947 = _T_92 ? _GEN_21939 : _GEN_21659; // @[sequencer-master.scala 154:24]
  wire  _GEN_21948 = _T_92 ? _GEN_21940 : _GEN_21660; // @[sequencer-master.scala 154:24]
  wire  _GEN_21949 = _T_92 ? _GEN_21941 : _GEN_21661; // @[sequencer-master.scala 154:24]
  wire  _GEN_21950 = _GEN_32729 | _GEN_21678; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21951 = _GEN_32730 | _GEN_21679; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21952 = _GEN_32731 | _GEN_21680; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21953 = _GEN_32732 | _GEN_21681; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21954 = _GEN_32733 | _GEN_21682; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21955 = _GEN_32734 | _GEN_21683; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21956 = _GEN_32735 | _GEN_21684; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21957 = _GEN_32736 | _GEN_21685; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21958 = _T_114 ? _GEN_21950 : _GEN_21678; // @[sequencer-master.scala 154:24]
  wire  _GEN_21959 = _T_114 ? _GEN_21951 : _GEN_21679; // @[sequencer-master.scala 154:24]
  wire  _GEN_21960 = _T_114 ? _GEN_21952 : _GEN_21680; // @[sequencer-master.scala 154:24]
  wire  _GEN_21961 = _T_114 ? _GEN_21953 : _GEN_21681; // @[sequencer-master.scala 154:24]
  wire  _GEN_21962 = _T_114 ? _GEN_21954 : _GEN_21682; // @[sequencer-master.scala 154:24]
  wire  _GEN_21963 = _T_114 ? _GEN_21955 : _GEN_21683; // @[sequencer-master.scala 154:24]
  wire  _GEN_21964 = _T_114 ? _GEN_21956 : _GEN_21684; // @[sequencer-master.scala 154:24]
  wire  _GEN_21965 = _T_114 ? _GEN_21957 : _GEN_21685; // @[sequencer-master.scala 154:24]
  wire  _GEN_21966 = _GEN_32729 | _GEN_21702; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21967 = _GEN_32730 | _GEN_21703; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21968 = _GEN_32731 | _GEN_21704; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21969 = _GEN_32732 | _GEN_21705; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21970 = _GEN_32733 | _GEN_21706; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21971 = _GEN_32734 | _GEN_21707; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21972 = _GEN_32735 | _GEN_21708; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21973 = _GEN_32736 | _GEN_21709; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21974 = _T_136 ? _GEN_21966 : _GEN_21702; // @[sequencer-master.scala 154:24]
  wire  _GEN_21975 = _T_136 ? _GEN_21967 : _GEN_21703; // @[sequencer-master.scala 154:24]
  wire  _GEN_21976 = _T_136 ? _GEN_21968 : _GEN_21704; // @[sequencer-master.scala 154:24]
  wire  _GEN_21977 = _T_136 ? _GEN_21969 : _GEN_21705; // @[sequencer-master.scala 154:24]
  wire  _GEN_21978 = _T_136 ? _GEN_21970 : _GEN_21706; // @[sequencer-master.scala 154:24]
  wire  _GEN_21979 = _T_136 ? _GEN_21971 : _GEN_21707; // @[sequencer-master.scala 154:24]
  wire  _GEN_21980 = _T_136 ? _GEN_21972 : _GEN_21708; // @[sequencer-master.scala 154:24]
  wire  _GEN_21981 = _T_136 ? _GEN_21973 : _GEN_21709; // @[sequencer-master.scala 154:24]
  wire  _GEN_21982 = _GEN_32729 | _GEN_21726; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21983 = _GEN_32730 | _GEN_21727; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21984 = _GEN_32731 | _GEN_21728; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21985 = _GEN_32732 | _GEN_21729; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21986 = _GEN_32733 | _GEN_21730; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21987 = _GEN_32734 | _GEN_21731; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21988 = _GEN_32735 | _GEN_21732; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21989 = _GEN_32736 | _GEN_21733; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21990 = _T_158 ? _GEN_21982 : _GEN_21726; // @[sequencer-master.scala 154:24]
  wire  _GEN_21991 = _T_158 ? _GEN_21983 : _GEN_21727; // @[sequencer-master.scala 154:24]
  wire  _GEN_21992 = _T_158 ? _GEN_21984 : _GEN_21728; // @[sequencer-master.scala 154:24]
  wire  _GEN_21993 = _T_158 ? _GEN_21985 : _GEN_21729; // @[sequencer-master.scala 154:24]
  wire  _GEN_21994 = _T_158 ? _GEN_21986 : _GEN_21730; // @[sequencer-master.scala 154:24]
  wire  _GEN_21995 = _T_158 ? _GEN_21987 : _GEN_21731; // @[sequencer-master.scala 154:24]
  wire  _GEN_21996 = _T_158 ? _GEN_21988 : _GEN_21732; // @[sequencer-master.scala 154:24]
  wire  _GEN_21997 = _T_158 ? _GEN_21989 : _GEN_21733; // @[sequencer-master.scala 154:24]
  wire  _GEN_21998 = _GEN_32729 | _GEN_21750; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_21999 = _GEN_32730 | _GEN_21751; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22000 = _GEN_32731 | _GEN_21752; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22001 = _GEN_32732 | _GEN_21753; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22002 = _GEN_32733 | _GEN_21754; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22003 = _GEN_32734 | _GEN_21755; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22004 = _GEN_32735 | _GEN_21756; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22005 = _GEN_32736 | _GEN_21757; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22006 = _T_180 ? _GEN_21998 : _GEN_21750; // @[sequencer-master.scala 154:24]
  wire  _GEN_22007 = _T_180 ? _GEN_21999 : _GEN_21751; // @[sequencer-master.scala 154:24]
  wire  _GEN_22008 = _T_180 ? _GEN_22000 : _GEN_21752; // @[sequencer-master.scala 154:24]
  wire  _GEN_22009 = _T_180 ? _GEN_22001 : _GEN_21753; // @[sequencer-master.scala 154:24]
  wire  _GEN_22010 = _T_180 ? _GEN_22002 : _GEN_21754; // @[sequencer-master.scala 154:24]
  wire  _GEN_22011 = _T_180 ? _GEN_22003 : _GEN_21755; // @[sequencer-master.scala 154:24]
  wire  _GEN_22012 = _T_180 ? _GEN_22004 : _GEN_21756; // @[sequencer-master.scala 154:24]
  wire  _GEN_22013 = _T_180 ? _GEN_22005 : _GEN_21757; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_22014 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_21380; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22015 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_21381; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22016 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_21382; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22017 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_21383; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22018 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_21384; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22019 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_21385; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22020 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_21386; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22021 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_21387; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22022 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_21542; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22023 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_21543; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22024 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_21544; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22025 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_21545; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22026 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_21546; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22027 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_21547; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22028 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_21548; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22029 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_21549; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22030 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_21388; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22031 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_21389; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22032 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_21390; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22033 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_21391; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22034 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_21392; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22035 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_21393; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22036 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_21394; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22037 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_21395; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22038 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_21396; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22039 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_21397; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22040 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_21398; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22041 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_21399; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22042 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_21400; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22043 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_21401; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22044 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_21402; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_22045 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_21403; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22046 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_21404; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22047 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_21405; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22048 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_21406; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22049 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_21407; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22050 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_21408; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22051 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_21409; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22052 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_21410; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_22053 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_21411; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_22054 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_21412; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22055 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_21413; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22056 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_21414; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22057 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_21415; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22058 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_21416; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22059 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_21417; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22060 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_21418; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_22061 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_21419; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_22062 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_21420; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22063 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_21421; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22064 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_21422; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22065 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_21423; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22066 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_21424; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22067 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_21425; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22068 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_21426; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22069 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_21427; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_22070 = _T_366 ? _GEN_22062 : _GEN_21420; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22071 = _T_366 ? _GEN_22063 : _GEN_21421; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22072 = _T_366 ? _GEN_22064 : _GEN_21422; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22073 = _T_366 ? _GEN_22065 : _GEN_21423; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22074 = _T_366 ? _GEN_22066 : _GEN_21424; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22075 = _T_366 ? _GEN_22067 : _GEN_21425; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22076 = _T_366 ? _GEN_22068 : _GEN_21426; // @[sequencer-master.scala 331:55]
  wire [63:0] _GEN_22077 = _T_366 ? _GEN_22069 : _GEN_21427; // @[sequencer-master.scala 331:55]
  wire [7:0] _GEN_22078 = io_op_bits_base_vs2_valid ? _GEN_22014 : _GEN_21380; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22079 = io_op_bits_base_vs2_valid ? _GEN_22015 : _GEN_21381; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22080 = io_op_bits_base_vs2_valid ? _GEN_22016 : _GEN_21382; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22081 = io_op_bits_base_vs2_valid ? _GEN_22017 : _GEN_21383; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22082 = io_op_bits_base_vs2_valid ? _GEN_22018 : _GEN_21384; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22083 = io_op_bits_base_vs2_valid ? _GEN_22019 : _GEN_21385; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22084 = io_op_bits_base_vs2_valid ? _GEN_22020 : _GEN_21386; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22085 = io_op_bits_base_vs2_valid ? _GEN_22021 : _GEN_21387; // @[sequencer-master.scala 328:47]
  wire  _GEN_22086 = io_op_bits_base_vs2_valid ? _GEN_22022 : _GEN_21542; // @[sequencer-master.scala 328:47]
  wire  _GEN_22087 = io_op_bits_base_vs2_valid ? _GEN_22023 : _GEN_21543; // @[sequencer-master.scala 328:47]
  wire  _GEN_22088 = io_op_bits_base_vs2_valid ? _GEN_22024 : _GEN_21544; // @[sequencer-master.scala 328:47]
  wire  _GEN_22089 = io_op_bits_base_vs2_valid ? _GEN_22025 : _GEN_21545; // @[sequencer-master.scala 328:47]
  wire  _GEN_22090 = io_op_bits_base_vs2_valid ? _GEN_22026 : _GEN_21546; // @[sequencer-master.scala 328:47]
  wire  _GEN_22091 = io_op_bits_base_vs2_valid ? _GEN_22027 : _GEN_21547; // @[sequencer-master.scala 328:47]
  wire  _GEN_22092 = io_op_bits_base_vs2_valid ? _GEN_22028 : _GEN_21548; // @[sequencer-master.scala 328:47]
  wire  _GEN_22093 = io_op_bits_base_vs2_valid ? _GEN_22029 : _GEN_21549; // @[sequencer-master.scala 328:47]
  wire  _GEN_22094 = io_op_bits_base_vs2_valid ? _GEN_22030 : _GEN_21388; // @[sequencer-master.scala 328:47]
  wire  _GEN_22095 = io_op_bits_base_vs2_valid ? _GEN_22031 : _GEN_21389; // @[sequencer-master.scala 328:47]
  wire  _GEN_22096 = io_op_bits_base_vs2_valid ? _GEN_22032 : _GEN_21390; // @[sequencer-master.scala 328:47]
  wire  _GEN_22097 = io_op_bits_base_vs2_valid ? _GEN_22033 : _GEN_21391; // @[sequencer-master.scala 328:47]
  wire  _GEN_22098 = io_op_bits_base_vs2_valid ? _GEN_22034 : _GEN_21392; // @[sequencer-master.scala 328:47]
  wire  _GEN_22099 = io_op_bits_base_vs2_valid ? _GEN_22035 : _GEN_21393; // @[sequencer-master.scala 328:47]
  wire  _GEN_22100 = io_op_bits_base_vs2_valid ? _GEN_22036 : _GEN_21394; // @[sequencer-master.scala 328:47]
  wire  _GEN_22101 = io_op_bits_base_vs2_valid ? _GEN_22037 : _GEN_21395; // @[sequencer-master.scala 328:47]
  wire  _GEN_22102 = io_op_bits_base_vs2_valid ? _GEN_22038 : _GEN_21396; // @[sequencer-master.scala 328:47]
  wire  _GEN_22103 = io_op_bits_base_vs2_valid ? _GEN_22039 : _GEN_21397; // @[sequencer-master.scala 328:47]
  wire  _GEN_22104 = io_op_bits_base_vs2_valid ? _GEN_22040 : _GEN_21398; // @[sequencer-master.scala 328:47]
  wire  _GEN_22105 = io_op_bits_base_vs2_valid ? _GEN_22041 : _GEN_21399; // @[sequencer-master.scala 328:47]
  wire  _GEN_22106 = io_op_bits_base_vs2_valid ? _GEN_22042 : _GEN_21400; // @[sequencer-master.scala 328:47]
  wire  _GEN_22107 = io_op_bits_base_vs2_valid ? _GEN_22043 : _GEN_21401; // @[sequencer-master.scala 328:47]
  wire  _GEN_22108 = io_op_bits_base_vs2_valid ? _GEN_22044 : _GEN_21402; // @[sequencer-master.scala 328:47]
  wire  _GEN_22109 = io_op_bits_base_vs2_valid ? _GEN_22045 : _GEN_21403; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22110 = io_op_bits_base_vs2_valid ? _GEN_22046 : _GEN_21404; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22111 = io_op_bits_base_vs2_valid ? _GEN_22047 : _GEN_21405; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22112 = io_op_bits_base_vs2_valid ? _GEN_22048 : _GEN_21406; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22113 = io_op_bits_base_vs2_valid ? _GEN_22049 : _GEN_21407; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22114 = io_op_bits_base_vs2_valid ? _GEN_22050 : _GEN_21408; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22115 = io_op_bits_base_vs2_valid ? _GEN_22051 : _GEN_21409; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22116 = io_op_bits_base_vs2_valid ? _GEN_22052 : _GEN_21410; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_22117 = io_op_bits_base_vs2_valid ? _GEN_22053 : _GEN_21411; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22118 = io_op_bits_base_vs2_valid ? _GEN_22054 : _GEN_21412; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22119 = io_op_bits_base_vs2_valid ? _GEN_22055 : _GEN_21413; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22120 = io_op_bits_base_vs2_valid ? _GEN_22056 : _GEN_21414; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22121 = io_op_bits_base_vs2_valid ? _GEN_22057 : _GEN_21415; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22122 = io_op_bits_base_vs2_valid ? _GEN_22058 : _GEN_21416; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22123 = io_op_bits_base_vs2_valid ? _GEN_22059 : _GEN_21417; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22124 = io_op_bits_base_vs2_valid ? _GEN_22060 : _GEN_21418; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_22125 = io_op_bits_base_vs2_valid ? _GEN_22061 : _GEN_21419; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22126 = io_op_bits_base_vs2_valid ? _GEN_22070 : _GEN_21420; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22127 = io_op_bits_base_vs2_valid ? _GEN_22071 : _GEN_21421; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22128 = io_op_bits_base_vs2_valid ? _GEN_22072 : _GEN_21422; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22129 = io_op_bits_base_vs2_valid ? _GEN_22073 : _GEN_21423; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22130 = io_op_bits_base_vs2_valid ? _GEN_22074 : _GEN_21424; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22131 = io_op_bits_base_vs2_valid ? _GEN_22075 : _GEN_21425; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22132 = io_op_bits_base_vs2_valid ? _GEN_22076 : _GEN_21426; // @[sequencer-master.scala 328:47]
  wire [63:0] _GEN_22133 = io_op_bits_base_vs2_valid ? _GEN_22077 : _GEN_21427; // @[sequencer-master.scala 328:47]
  wire  _GEN_22134 = _GEN_32729 | _GEN_21894; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22135 = _GEN_32730 | _GEN_21895; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22136 = _GEN_32731 | _GEN_21896; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22137 = _GEN_32732 | _GEN_21897; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22138 = _GEN_32733 | _GEN_21898; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22139 = _GEN_32734 | _GEN_21899; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22140 = _GEN_32735 | _GEN_21900; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22141 = _GEN_32736 | _GEN_21901; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22142 = _T_380 ? _GEN_22134 : _GEN_21894; // @[sequencer-master.scala 154:24]
  wire  _GEN_22143 = _T_380 ? _GEN_22135 : _GEN_21895; // @[sequencer-master.scala 154:24]
  wire  _GEN_22144 = _T_380 ? _GEN_22136 : _GEN_21896; // @[sequencer-master.scala 154:24]
  wire  _GEN_22145 = _T_380 ? _GEN_22137 : _GEN_21897; // @[sequencer-master.scala 154:24]
  wire  _GEN_22146 = _T_380 ? _GEN_22138 : _GEN_21898; // @[sequencer-master.scala 154:24]
  wire  _GEN_22147 = _T_380 ? _GEN_22139 : _GEN_21899; // @[sequencer-master.scala 154:24]
  wire  _GEN_22148 = _T_380 ? _GEN_22140 : _GEN_21900; // @[sequencer-master.scala 154:24]
  wire  _GEN_22149 = _T_380 ? _GEN_22141 : _GEN_21901; // @[sequencer-master.scala 154:24]
  wire  _GEN_22150 = _GEN_32729 | _GEN_21910; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22151 = _GEN_32730 | _GEN_21911; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22152 = _GEN_32731 | _GEN_21912; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22153 = _GEN_32732 | _GEN_21913; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22154 = _GEN_32733 | _GEN_21914; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22155 = _GEN_32734 | _GEN_21915; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22156 = _GEN_32735 | _GEN_21916; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22157 = _GEN_32736 | _GEN_21917; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22158 = _T_402 ? _GEN_22150 : _GEN_21910; // @[sequencer-master.scala 154:24]
  wire  _GEN_22159 = _T_402 ? _GEN_22151 : _GEN_21911; // @[sequencer-master.scala 154:24]
  wire  _GEN_22160 = _T_402 ? _GEN_22152 : _GEN_21912; // @[sequencer-master.scala 154:24]
  wire  _GEN_22161 = _T_402 ? _GEN_22153 : _GEN_21913; // @[sequencer-master.scala 154:24]
  wire  _GEN_22162 = _T_402 ? _GEN_22154 : _GEN_21914; // @[sequencer-master.scala 154:24]
  wire  _GEN_22163 = _T_402 ? _GEN_22155 : _GEN_21915; // @[sequencer-master.scala 154:24]
  wire  _GEN_22164 = _T_402 ? _GEN_22156 : _GEN_21916; // @[sequencer-master.scala 154:24]
  wire  _GEN_22165 = _T_402 ? _GEN_22157 : _GEN_21917; // @[sequencer-master.scala 154:24]
  wire  _GEN_22166 = _GEN_32729 | _GEN_21926; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22167 = _GEN_32730 | _GEN_21927; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22168 = _GEN_32731 | _GEN_21928; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22169 = _GEN_32732 | _GEN_21929; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22170 = _GEN_32733 | _GEN_21930; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22171 = _GEN_32734 | _GEN_21931; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22172 = _GEN_32735 | _GEN_21932; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22173 = _GEN_32736 | _GEN_21933; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22174 = _T_424 ? _GEN_22166 : _GEN_21926; // @[sequencer-master.scala 154:24]
  wire  _GEN_22175 = _T_424 ? _GEN_22167 : _GEN_21927; // @[sequencer-master.scala 154:24]
  wire  _GEN_22176 = _T_424 ? _GEN_22168 : _GEN_21928; // @[sequencer-master.scala 154:24]
  wire  _GEN_22177 = _T_424 ? _GEN_22169 : _GEN_21929; // @[sequencer-master.scala 154:24]
  wire  _GEN_22178 = _T_424 ? _GEN_22170 : _GEN_21930; // @[sequencer-master.scala 154:24]
  wire  _GEN_22179 = _T_424 ? _GEN_22171 : _GEN_21931; // @[sequencer-master.scala 154:24]
  wire  _GEN_22180 = _T_424 ? _GEN_22172 : _GEN_21932; // @[sequencer-master.scala 154:24]
  wire  _GEN_22181 = _T_424 ? _GEN_22173 : _GEN_21933; // @[sequencer-master.scala 154:24]
  wire  _GEN_22182 = _GEN_32729 | _GEN_21942; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22183 = _GEN_32730 | _GEN_21943; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22184 = _GEN_32731 | _GEN_21944; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22185 = _GEN_32732 | _GEN_21945; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22186 = _GEN_32733 | _GEN_21946; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22187 = _GEN_32734 | _GEN_21947; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22188 = _GEN_32735 | _GEN_21948; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22189 = _GEN_32736 | _GEN_21949; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22190 = _T_446 ? _GEN_22182 : _GEN_21942; // @[sequencer-master.scala 154:24]
  wire  _GEN_22191 = _T_446 ? _GEN_22183 : _GEN_21943; // @[sequencer-master.scala 154:24]
  wire  _GEN_22192 = _T_446 ? _GEN_22184 : _GEN_21944; // @[sequencer-master.scala 154:24]
  wire  _GEN_22193 = _T_446 ? _GEN_22185 : _GEN_21945; // @[sequencer-master.scala 154:24]
  wire  _GEN_22194 = _T_446 ? _GEN_22186 : _GEN_21946; // @[sequencer-master.scala 154:24]
  wire  _GEN_22195 = _T_446 ? _GEN_22187 : _GEN_21947; // @[sequencer-master.scala 154:24]
  wire  _GEN_22196 = _T_446 ? _GEN_22188 : _GEN_21948; // @[sequencer-master.scala 154:24]
  wire  _GEN_22197 = _T_446 ? _GEN_22189 : _GEN_21949; // @[sequencer-master.scala 154:24]
  wire  _GEN_22198 = _GEN_32729 | _GEN_21958; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22199 = _GEN_32730 | _GEN_21959; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22200 = _GEN_32731 | _GEN_21960; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22201 = _GEN_32732 | _GEN_21961; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22202 = _GEN_32733 | _GEN_21962; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22203 = _GEN_32734 | _GEN_21963; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22204 = _GEN_32735 | _GEN_21964; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22205 = _GEN_32736 | _GEN_21965; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22206 = _T_468 ? _GEN_22198 : _GEN_21958; // @[sequencer-master.scala 154:24]
  wire  _GEN_22207 = _T_468 ? _GEN_22199 : _GEN_21959; // @[sequencer-master.scala 154:24]
  wire  _GEN_22208 = _T_468 ? _GEN_22200 : _GEN_21960; // @[sequencer-master.scala 154:24]
  wire  _GEN_22209 = _T_468 ? _GEN_22201 : _GEN_21961; // @[sequencer-master.scala 154:24]
  wire  _GEN_22210 = _T_468 ? _GEN_22202 : _GEN_21962; // @[sequencer-master.scala 154:24]
  wire  _GEN_22211 = _T_468 ? _GEN_22203 : _GEN_21963; // @[sequencer-master.scala 154:24]
  wire  _GEN_22212 = _T_468 ? _GEN_22204 : _GEN_21964; // @[sequencer-master.scala 154:24]
  wire  _GEN_22213 = _T_468 ? _GEN_22205 : _GEN_21965; // @[sequencer-master.scala 154:24]
  wire  _GEN_22214 = _GEN_32729 | _GEN_21974; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22215 = _GEN_32730 | _GEN_21975; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22216 = _GEN_32731 | _GEN_21976; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22217 = _GEN_32732 | _GEN_21977; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22218 = _GEN_32733 | _GEN_21978; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22219 = _GEN_32734 | _GEN_21979; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22220 = _GEN_32735 | _GEN_21980; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22221 = _GEN_32736 | _GEN_21981; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22222 = _T_490 ? _GEN_22214 : _GEN_21974; // @[sequencer-master.scala 154:24]
  wire  _GEN_22223 = _T_490 ? _GEN_22215 : _GEN_21975; // @[sequencer-master.scala 154:24]
  wire  _GEN_22224 = _T_490 ? _GEN_22216 : _GEN_21976; // @[sequencer-master.scala 154:24]
  wire  _GEN_22225 = _T_490 ? _GEN_22217 : _GEN_21977; // @[sequencer-master.scala 154:24]
  wire  _GEN_22226 = _T_490 ? _GEN_22218 : _GEN_21978; // @[sequencer-master.scala 154:24]
  wire  _GEN_22227 = _T_490 ? _GEN_22219 : _GEN_21979; // @[sequencer-master.scala 154:24]
  wire  _GEN_22228 = _T_490 ? _GEN_22220 : _GEN_21980; // @[sequencer-master.scala 154:24]
  wire  _GEN_22229 = _T_490 ? _GEN_22221 : _GEN_21981; // @[sequencer-master.scala 154:24]
  wire  _GEN_22230 = _GEN_32729 | _GEN_21990; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22231 = _GEN_32730 | _GEN_21991; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22232 = _GEN_32731 | _GEN_21992; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22233 = _GEN_32732 | _GEN_21993; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22234 = _GEN_32733 | _GEN_21994; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22235 = _GEN_32734 | _GEN_21995; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22236 = _GEN_32735 | _GEN_21996; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22237 = _GEN_32736 | _GEN_21997; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22238 = _T_512 ? _GEN_22230 : _GEN_21990; // @[sequencer-master.scala 154:24]
  wire  _GEN_22239 = _T_512 ? _GEN_22231 : _GEN_21991; // @[sequencer-master.scala 154:24]
  wire  _GEN_22240 = _T_512 ? _GEN_22232 : _GEN_21992; // @[sequencer-master.scala 154:24]
  wire  _GEN_22241 = _T_512 ? _GEN_22233 : _GEN_21993; // @[sequencer-master.scala 154:24]
  wire  _GEN_22242 = _T_512 ? _GEN_22234 : _GEN_21994; // @[sequencer-master.scala 154:24]
  wire  _GEN_22243 = _T_512 ? _GEN_22235 : _GEN_21995; // @[sequencer-master.scala 154:24]
  wire  _GEN_22244 = _T_512 ? _GEN_22236 : _GEN_21996; // @[sequencer-master.scala 154:24]
  wire  _GEN_22245 = _T_512 ? _GEN_22237 : _GEN_21997; // @[sequencer-master.scala 154:24]
  wire  _GEN_22246 = _GEN_32729 | _GEN_22006; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22247 = _GEN_32730 | _GEN_22007; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22248 = _GEN_32731 | _GEN_22008; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22249 = _GEN_32732 | _GEN_22009; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22250 = _GEN_32733 | _GEN_22010; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22251 = _GEN_32734 | _GEN_22011; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22252 = _GEN_32735 | _GEN_22012; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22253 = _GEN_32736 | _GEN_22013; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_22254 = _T_534 ? _GEN_22246 : _GEN_22006; // @[sequencer-master.scala 154:24]
  wire  _GEN_22255 = _T_534 ? _GEN_22247 : _GEN_22007; // @[sequencer-master.scala 154:24]
  wire  _GEN_22256 = _T_534 ? _GEN_22248 : _GEN_22008; // @[sequencer-master.scala 154:24]
  wire  _GEN_22257 = _T_534 ? _GEN_22249 : _GEN_22009; // @[sequencer-master.scala 154:24]
  wire  _GEN_22258 = _T_534 ? _GEN_22250 : _GEN_22010; // @[sequencer-master.scala 154:24]
  wire  _GEN_22259 = _T_534 ? _GEN_22251 : _GEN_22011; // @[sequencer-master.scala 154:24]
  wire  _GEN_22260 = _T_534 ? _GEN_22252 : _GEN_22012; // @[sequencer-master.scala 154:24]
  wire  _GEN_22261 = _T_534 ? _GEN_22253 : _GEN_22013; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_22262 = 3'h0 == tail ? _e_T_1647_rports : _GEN_21428; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22263 = 3'h1 == tail ? _e_T_1647_rports : _GEN_21429; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22264 = 3'h2 == tail ? _e_T_1647_rports : _GEN_21430; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22265 = 3'h3 == tail ? _e_T_1647_rports : _GEN_21431; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22266 = 3'h4 == tail ? _e_T_1647_rports : _GEN_21432; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22267 = 3'h5 == tail ? _e_T_1647_rports : _GEN_21433; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22268 = 3'h6 == tail ? _e_T_1647_rports : _GEN_21434; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22269 = 3'h7 == tail ? _e_T_1647_rports : _GEN_21435; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_22270 = 3'h0 == tail ? 4'h0 : _GEN_21436; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22271 = 3'h1 == tail ? 4'h0 : _GEN_21437; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22272 = 3'h2 == tail ? 4'h0 : _GEN_21438; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22273 = 3'h3 == tail ? 4'h0 : _GEN_21439; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22274 = 3'h4 == tail ? 4'h0 : _GEN_21440; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22275 = 3'h5 == tail ? 4'h0 : _GEN_21441; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22276 = 3'h6 == tail ? 4'h0 : _GEN_21442; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22277 = 3'h7 == tail ? 4'h0 : _GEN_21443; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_22278 = 3'h0 == tail ? 3'h0 : _GEN_21444; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22279 = 3'h1 == tail ? 3'h0 : _GEN_21445; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22280 = 3'h2 == tail ? 3'h0 : _GEN_21446; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22281 = 3'h3 == tail ? 3'h0 : _GEN_21447; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22282 = 3'h4 == tail ? 3'h0 : _GEN_21448; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22283 = 3'h5 == tail ? 3'h0 : _GEN_21449; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22284 = 3'h6 == tail ? 3'h0 : _GEN_21450; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22285 = 3'h7 == tail ? 3'h0 : _GEN_21451; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_22302 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21854; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22303 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21855; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22304 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21856; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22305 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21857; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22306 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21858; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22307 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21859; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22308 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21860; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22309 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21861; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22310 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22086; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22311 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22087; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22312 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22088; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22313 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22089; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22314 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22090; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22315 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22091; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22316 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22092; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22317 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22093; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22318 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21550; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22319 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21551; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22320 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21552; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22321 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21553; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22322 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21554; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22323 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21555; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22324 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21556; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22325 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21557; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22326 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21558; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22327 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21559; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22328 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21560; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22329 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21561; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22330 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21562; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22331 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21563; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22332 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21564; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22333 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21565; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22334 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21566; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22335 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21567; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22336 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21568; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22337 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21569; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22338 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21570; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22339 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21571; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22340 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21572; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22341 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21573; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22350 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22142; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22351 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22143; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22352 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22144; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22353 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22145; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22354 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22146; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22355 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22147; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22356 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22148; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22357 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22149; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22358 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21590; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22359 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21591; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22360 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21592; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22361 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21593; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22362 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21594; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22363 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21595; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22364 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21596; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22365 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21597; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22366 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21598; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22367 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21599; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22368 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21600; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22369 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21601; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22370 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21602; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22371 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21603; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22372 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21604; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22373 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21605; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22374 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22158; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22375 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22159; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22376 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22160; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22377 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22161; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22378 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22162; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22379 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22163; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22380 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22164; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22381 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22165; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22382 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21614; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22383 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21615; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22384 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21616; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22385 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21617; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22386 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21618; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22387 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21619; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22388 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21620; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22389 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21621; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22390 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21622; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22391 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21623; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22392 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21624; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22393 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21625; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22394 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21626; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22395 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21627; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22396 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21628; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22397 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21629; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22398 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22174; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22399 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22175; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22400 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22176; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22401 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22177; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22402 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22178; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22403 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22179; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22404 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22180; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22405 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22181; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22406 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21638; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22407 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21639; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22408 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21640; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22409 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21641; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22410 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21642; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22411 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21643; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22412 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21644; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22413 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21645; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22414 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21646; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22415 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21647; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22416 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21648; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22417 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21649; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22418 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21650; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22419 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21651; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22420 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21652; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22421 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21653; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22422 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22190; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22423 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22191; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22424 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22192; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22425 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22193; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22426 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22194; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22427 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22195; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22428 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22196; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22429 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22197; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22430 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21662; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22431 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21663; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22432 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21664; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22433 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21665; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22434 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21666; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22435 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21667; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22436 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21668; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22437 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21669; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22438 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21670; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22439 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21671; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22440 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21672; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22441 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21673; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22442 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21674; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22443 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21675; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22444 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21676; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22445 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21677; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22446 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22206; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22447 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22207; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22448 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22208; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22449 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22209; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22450 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22210; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22451 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22211; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22452 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22212; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22453 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22213; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22454 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21686; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22455 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21687; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22456 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21688; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22457 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21689; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22458 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21690; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22459 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21691; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22460 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21692; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22461 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21693; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22462 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21694; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22463 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21695; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22464 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21696; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22465 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21697; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22466 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21698; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22467 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21699; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22468 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21700; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22469 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21701; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22470 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22222; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22471 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22223; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22472 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22224; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22473 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22225; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22474 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22226; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22475 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22227; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22476 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22228; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22477 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22229; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22478 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21710; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22479 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21711; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22480 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21712; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22481 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21713; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22482 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21714; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22483 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21715; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22484 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21716; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22485 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21717; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22486 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21718; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22487 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21719; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22488 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21720; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22489 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21721; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22490 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21722; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22491 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21723; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22492 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21724; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22493 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21725; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22494 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22238; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22495 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22239; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22496 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22240; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22497 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22241; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22498 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22242; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22499 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22243; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22500 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22244; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22501 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22245; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22502 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21734; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22503 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21735; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22504 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21736; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22505 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21737; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22506 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21738; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22507 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21739; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22508 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21740; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22509 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21741; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22510 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21742; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22511 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21743; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22512 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21744; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22513 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21745; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22514 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21746; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22515 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21747; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22516 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21748; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22517 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21749; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22518 = 3'h0 == _T_1645 ? 1'h0 : _GEN_22254; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22519 = 3'h1 == _T_1645 ? 1'h0 : _GEN_22255; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22520 = 3'h2 == _T_1645 ? 1'h0 : _GEN_22256; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22521 = 3'h3 == _T_1645 ? 1'h0 : _GEN_22257; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22522 = 3'h4 == _T_1645 ? 1'h0 : _GEN_22258; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22523 = 3'h5 == _T_1645 ? 1'h0 : _GEN_22259; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22524 = 3'h6 == _T_1645 ? 1'h0 : _GEN_22260; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22525 = 3'h7 == _T_1645 ? 1'h0 : _GEN_22261; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22526 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21758; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22527 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21759; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22528 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21760; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22529 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21761; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22530 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21762; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22531 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21763; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22532 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21764; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22533 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21765; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22534 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21766; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22535 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21767; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22536 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21768; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22537 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21769; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22538 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21770; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22539 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21771; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22540 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21772; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22541 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21773; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22542 = 3'h0 == _T_1645 ? 1'h0 : _GEN_21774; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22543 = 3'h1 == _T_1645 ? 1'h0 : _GEN_21775; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22544 = 3'h2 == _T_1645 ? 1'h0 : _GEN_21776; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22545 = 3'h3 == _T_1645 ? 1'h0 : _GEN_21777; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22546 = 3'h4 == _T_1645 ? 1'h0 : _GEN_21778; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22547 = 3'h5 == _T_1645 ? 1'h0 : _GEN_21779; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22548 = 3'h6 == _T_1645 ? 1'h0 : _GEN_21780; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22549 = 3'h7 == _T_1645 ? 1'h0 : _GEN_21781; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_22558 = _GEN_34121 | _GEN_21452; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22559 = _GEN_34122 | _GEN_21453; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22560 = _GEN_34123 | _GEN_21454; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22561 = _GEN_34124 | _GEN_21455; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22562 = _GEN_34125 | _GEN_21456; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22563 = _GEN_34126 | _GEN_21457; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22564 = _GEN_34127 | _GEN_21458; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_22565 = _GEN_34128 | _GEN_21459; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_22566 = 3'h0 == _T_1645 ? io_op_bits_fn_union : _GEN_21798; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22567 = 3'h1 == _T_1645 ? io_op_bits_fn_union : _GEN_21799; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22568 = 3'h2 == _T_1645 ? io_op_bits_fn_union : _GEN_21800; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22569 = 3'h3 == _T_1645 ? io_op_bits_fn_union : _GEN_21801; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22570 = 3'h4 == _T_1645 ? io_op_bits_fn_union : _GEN_21802; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22571 = 3'h5 == _T_1645 ? io_op_bits_fn_union : _GEN_21803; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22572 = 3'h6 == _T_1645 ? io_op_bits_fn_union : _GEN_21804; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_22573 = 3'h7 == _T_1645 ? io_op_bits_fn_union : _GEN_21805; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [1:0] _GEN_22574 = 3'h0 == _T_1645 ? 2'h0 : _GEN_22262; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22575 = 3'h1 == _T_1645 ? 2'h0 : _GEN_22263; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22576 = 3'h2 == _T_1645 ? 2'h0 : _GEN_22264; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22577 = 3'h3 == _T_1645 ? 2'h0 : _GEN_22265; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22578 = 3'h4 == _T_1645 ? 2'h0 : _GEN_22266; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22579 = 3'h5 == _T_1645 ? 2'h0 : _GEN_22267; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22580 = 3'h6 == _T_1645 ? 2'h0 : _GEN_22268; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_22581 = 3'h7 == _T_1645 ? 2'h0 : _GEN_22269; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_22582 = 3'h0 == _T_1645 ? 4'h0 : _GEN_22270; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22583 = 3'h1 == _T_1645 ? 4'h0 : _GEN_22271; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22584 = 3'h2 == _T_1645 ? 4'h0 : _GEN_22272; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22585 = 3'h3 == _T_1645 ? 4'h0 : _GEN_22273; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22586 = 3'h4 == _T_1645 ? 4'h0 : _GEN_22274; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22587 = 3'h5 == _T_1645 ? 4'h0 : _GEN_22275; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22588 = 3'h6 == _T_1645 ? 4'h0 : _GEN_22276; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_22589 = 3'h7 == _T_1645 ? 4'h0 : _GEN_22277; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_22590 = 3'h0 == _T_1645 ? 3'h0 : _GEN_22278; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22591 = 3'h1 == _T_1645 ? 3'h0 : _GEN_22279; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22592 = 3'h2 == _T_1645 ? 3'h0 : _GEN_22280; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22593 = 3'h3 == _T_1645 ? 3'h0 : _GEN_22281; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22594 = 3'h4 == _T_1645 ? 3'h0 : _GEN_22282; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22595 = 3'h5 == _T_1645 ? 3'h0 : _GEN_22283; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22596 = 3'h6 == _T_1645 ? 3'h0 : _GEN_22284; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_22597 = 3'h7 == _T_1645 ? 3'h0 : _GEN_22285; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_22598 = _GEN_34121 | _GEN_22358; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22599 = _GEN_34122 | _GEN_22359; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22600 = _GEN_34123 | _GEN_22360; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22601 = _GEN_34124 | _GEN_22361; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22602 = _GEN_34125 | _GEN_22362; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22603 = _GEN_34126 | _GEN_22363; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22604 = _GEN_34127 | _GEN_22364; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22605 = _GEN_34128 | _GEN_22365; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22606 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22598 : _GEN_22358; // @[sequencer-master.scala 161:86]
  wire  _GEN_22607 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22599 : _GEN_22359; // @[sequencer-master.scala 161:86]
  wire  _GEN_22608 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22600 : _GEN_22360; // @[sequencer-master.scala 161:86]
  wire  _GEN_22609 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22601 : _GEN_22361; // @[sequencer-master.scala 161:86]
  wire  _GEN_22610 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22602 : _GEN_22362; // @[sequencer-master.scala 161:86]
  wire  _GEN_22611 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22603 : _GEN_22363; // @[sequencer-master.scala 161:86]
  wire  _GEN_22612 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22604 : _GEN_22364; // @[sequencer-master.scala 161:86]
  wire  _GEN_22613 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_22605 : _GEN_22365; // @[sequencer-master.scala 161:86]
  wire  _GEN_22614 = _GEN_34121 | _GEN_22382; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22615 = _GEN_34122 | _GEN_22383; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22616 = _GEN_34123 | _GEN_22384; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22617 = _GEN_34124 | _GEN_22385; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22618 = _GEN_34125 | _GEN_22386; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22619 = _GEN_34126 | _GEN_22387; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22620 = _GEN_34127 | _GEN_22388; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22621 = _GEN_34128 | _GEN_22389; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22622 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22614 : _GEN_22382; // @[sequencer-master.scala 161:86]
  wire  _GEN_22623 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22615 : _GEN_22383; // @[sequencer-master.scala 161:86]
  wire  _GEN_22624 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22616 : _GEN_22384; // @[sequencer-master.scala 161:86]
  wire  _GEN_22625 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22617 : _GEN_22385; // @[sequencer-master.scala 161:86]
  wire  _GEN_22626 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22618 : _GEN_22386; // @[sequencer-master.scala 161:86]
  wire  _GEN_22627 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22619 : _GEN_22387; // @[sequencer-master.scala 161:86]
  wire  _GEN_22628 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22620 : _GEN_22388; // @[sequencer-master.scala 161:86]
  wire  _GEN_22629 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_22621 : _GEN_22389; // @[sequencer-master.scala 161:86]
  wire  _GEN_22630 = _GEN_34121 | _GEN_22406; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22631 = _GEN_34122 | _GEN_22407; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22632 = _GEN_34123 | _GEN_22408; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22633 = _GEN_34124 | _GEN_22409; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22634 = _GEN_34125 | _GEN_22410; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22635 = _GEN_34126 | _GEN_22411; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22636 = _GEN_34127 | _GEN_22412; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22637 = _GEN_34128 | _GEN_22413; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22638 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22630 : _GEN_22406; // @[sequencer-master.scala 161:86]
  wire  _GEN_22639 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22631 : _GEN_22407; // @[sequencer-master.scala 161:86]
  wire  _GEN_22640 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22632 : _GEN_22408; // @[sequencer-master.scala 161:86]
  wire  _GEN_22641 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22633 : _GEN_22409; // @[sequencer-master.scala 161:86]
  wire  _GEN_22642 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22634 : _GEN_22410; // @[sequencer-master.scala 161:86]
  wire  _GEN_22643 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22635 : _GEN_22411; // @[sequencer-master.scala 161:86]
  wire  _GEN_22644 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22636 : _GEN_22412; // @[sequencer-master.scala 161:86]
  wire  _GEN_22645 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_22637 : _GEN_22413; // @[sequencer-master.scala 161:86]
  wire  _GEN_22646 = _GEN_34121 | _GEN_22430; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22647 = _GEN_34122 | _GEN_22431; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22648 = _GEN_34123 | _GEN_22432; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22649 = _GEN_34124 | _GEN_22433; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22650 = _GEN_34125 | _GEN_22434; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22651 = _GEN_34126 | _GEN_22435; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22652 = _GEN_34127 | _GEN_22436; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22653 = _GEN_34128 | _GEN_22437; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22654 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22646 : _GEN_22430; // @[sequencer-master.scala 161:86]
  wire  _GEN_22655 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22647 : _GEN_22431; // @[sequencer-master.scala 161:86]
  wire  _GEN_22656 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22648 : _GEN_22432; // @[sequencer-master.scala 161:86]
  wire  _GEN_22657 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22649 : _GEN_22433; // @[sequencer-master.scala 161:86]
  wire  _GEN_22658 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22650 : _GEN_22434; // @[sequencer-master.scala 161:86]
  wire  _GEN_22659 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22651 : _GEN_22435; // @[sequencer-master.scala 161:86]
  wire  _GEN_22660 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22652 : _GEN_22436; // @[sequencer-master.scala 161:86]
  wire  _GEN_22661 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_22653 : _GEN_22437; // @[sequencer-master.scala 161:86]
  wire  _GEN_22662 = _GEN_34121 | _GEN_22454; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22663 = _GEN_34122 | _GEN_22455; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22664 = _GEN_34123 | _GEN_22456; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22665 = _GEN_34124 | _GEN_22457; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22666 = _GEN_34125 | _GEN_22458; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22667 = _GEN_34126 | _GEN_22459; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22668 = _GEN_34127 | _GEN_22460; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22669 = _GEN_34128 | _GEN_22461; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22670 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22662 : _GEN_22454; // @[sequencer-master.scala 161:86]
  wire  _GEN_22671 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22663 : _GEN_22455; // @[sequencer-master.scala 161:86]
  wire  _GEN_22672 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22664 : _GEN_22456; // @[sequencer-master.scala 161:86]
  wire  _GEN_22673 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22665 : _GEN_22457; // @[sequencer-master.scala 161:86]
  wire  _GEN_22674 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22666 : _GEN_22458; // @[sequencer-master.scala 161:86]
  wire  _GEN_22675 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22667 : _GEN_22459; // @[sequencer-master.scala 161:86]
  wire  _GEN_22676 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22668 : _GEN_22460; // @[sequencer-master.scala 161:86]
  wire  _GEN_22677 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_22669 : _GEN_22461; // @[sequencer-master.scala 161:86]
  wire  _GEN_22678 = _GEN_34121 | _GEN_22478; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22679 = _GEN_34122 | _GEN_22479; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22680 = _GEN_34123 | _GEN_22480; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22681 = _GEN_34124 | _GEN_22481; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22682 = _GEN_34125 | _GEN_22482; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22683 = _GEN_34126 | _GEN_22483; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22684 = _GEN_34127 | _GEN_22484; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22685 = _GEN_34128 | _GEN_22485; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22686 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22678 : _GEN_22478; // @[sequencer-master.scala 161:86]
  wire  _GEN_22687 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22679 : _GEN_22479; // @[sequencer-master.scala 161:86]
  wire  _GEN_22688 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22680 : _GEN_22480; // @[sequencer-master.scala 161:86]
  wire  _GEN_22689 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22681 : _GEN_22481; // @[sequencer-master.scala 161:86]
  wire  _GEN_22690 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22682 : _GEN_22482; // @[sequencer-master.scala 161:86]
  wire  _GEN_22691 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22683 : _GEN_22483; // @[sequencer-master.scala 161:86]
  wire  _GEN_22692 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22684 : _GEN_22484; // @[sequencer-master.scala 161:86]
  wire  _GEN_22693 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_22685 : _GEN_22485; // @[sequencer-master.scala 161:86]
  wire  _GEN_22694 = _GEN_34121 | _GEN_22502; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22695 = _GEN_34122 | _GEN_22503; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22696 = _GEN_34123 | _GEN_22504; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22697 = _GEN_34124 | _GEN_22505; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22698 = _GEN_34125 | _GEN_22506; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22699 = _GEN_34126 | _GEN_22507; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22700 = _GEN_34127 | _GEN_22508; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22701 = _GEN_34128 | _GEN_22509; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22702 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22694 : _GEN_22502; // @[sequencer-master.scala 161:86]
  wire  _GEN_22703 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22695 : _GEN_22503; // @[sequencer-master.scala 161:86]
  wire  _GEN_22704 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22696 : _GEN_22504; // @[sequencer-master.scala 161:86]
  wire  _GEN_22705 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22697 : _GEN_22505; // @[sequencer-master.scala 161:86]
  wire  _GEN_22706 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22698 : _GEN_22506; // @[sequencer-master.scala 161:86]
  wire  _GEN_22707 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22699 : _GEN_22507; // @[sequencer-master.scala 161:86]
  wire  _GEN_22708 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22700 : _GEN_22508; // @[sequencer-master.scala 161:86]
  wire  _GEN_22709 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_22701 : _GEN_22509; // @[sequencer-master.scala 161:86]
  wire  _GEN_22710 = _GEN_34121 | _GEN_22526; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22711 = _GEN_34122 | _GEN_22527; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22712 = _GEN_34123 | _GEN_22528; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22713 = _GEN_34124 | _GEN_22529; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22714 = _GEN_34125 | _GEN_22530; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22715 = _GEN_34126 | _GEN_22531; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22716 = _GEN_34127 | _GEN_22532; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22717 = _GEN_34128 | _GEN_22533; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_22718 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22710 : _GEN_22526; // @[sequencer-master.scala 161:86]
  wire  _GEN_22719 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22711 : _GEN_22527; // @[sequencer-master.scala 161:86]
  wire  _GEN_22720 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22712 : _GEN_22528; // @[sequencer-master.scala 161:86]
  wire  _GEN_22721 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22713 : _GEN_22529; // @[sequencer-master.scala 161:86]
  wire  _GEN_22722 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22714 : _GEN_22530; // @[sequencer-master.scala 161:86]
  wire  _GEN_22723 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22715 : _GEN_22531; // @[sequencer-master.scala 161:86]
  wire  _GEN_22724 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22716 : _GEN_22532; // @[sequencer-master.scala 161:86]
  wire  _GEN_22725 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_22717 : _GEN_22533; // @[sequencer-master.scala 161:86]
  wire  _GEN_22726 = _GEN_34121 | _GEN_22366; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22727 = _GEN_34122 | _GEN_22367; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22728 = _GEN_34123 | _GEN_22368; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22729 = _GEN_34124 | _GEN_22369; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22730 = _GEN_34125 | _GEN_22370; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22731 = _GEN_34126 | _GEN_22371; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22732 = _GEN_34127 | _GEN_22372; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22733 = _GEN_34128 | _GEN_22373; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22734 = _T_1442 ? _GEN_22726 : _GEN_22366; // @[sequencer-master.scala 168:32]
  wire  _GEN_22735 = _T_1442 ? _GEN_22727 : _GEN_22367; // @[sequencer-master.scala 168:32]
  wire  _GEN_22736 = _T_1442 ? _GEN_22728 : _GEN_22368; // @[sequencer-master.scala 168:32]
  wire  _GEN_22737 = _T_1442 ? _GEN_22729 : _GEN_22369; // @[sequencer-master.scala 168:32]
  wire  _GEN_22738 = _T_1442 ? _GEN_22730 : _GEN_22370; // @[sequencer-master.scala 168:32]
  wire  _GEN_22739 = _T_1442 ? _GEN_22731 : _GEN_22371; // @[sequencer-master.scala 168:32]
  wire  _GEN_22740 = _T_1442 ? _GEN_22732 : _GEN_22372; // @[sequencer-master.scala 168:32]
  wire  _GEN_22741 = _T_1442 ? _GEN_22733 : _GEN_22373; // @[sequencer-master.scala 168:32]
  wire  _GEN_22742 = _GEN_34121 | _GEN_22390; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22743 = _GEN_34122 | _GEN_22391; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22744 = _GEN_34123 | _GEN_22392; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22745 = _GEN_34124 | _GEN_22393; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22746 = _GEN_34125 | _GEN_22394; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22747 = _GEN_34126 | _GEN_22395; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22748 = _GEN_34127 | _GEN_22396; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22749 = _GEN_34128 | _GEN_22397; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22750 = _T_1464 ? _GEN_22742 : _GEN_22390; // @[sequencer-master.scala 168:32]
  wire  _GEN_22751 = _T_1464 ? _GEN_22743 : _GEN_22391; // @[sequencer-master.scala 168:32]
  wire  _GEN_22752 = _T_1464 ? _GEN_22744 : _GEN_22392; // @[sequencer-master.scala 168:32]
  wire  _GEN_22753 = _T_1464 ? _GEN_22745 : _GEN_22393; // @[sequencer-master.scala 168:32]
  wire  _GEN_22754 = _T_1464 ? _GEN_22746 : _GEN_22394; // @[sequencer-master.scala 168:32]
  wire  _GEN_22755 = _T_1464 ? _GEN_22747 : _GEN_22395; // @[sequencer-master.scala 168:32]
  wire  _GEN_22756 = _T_1464 ? _GEN_22748 : _GEN_22396; // @[sequencer-master.scala 168:32]
  wire  _GEN_22757 = _T_1464 ? _GEN_22749 : _GEN_22397; // @[sequencer-master.scala 168:32]
  wire  _GEN_22758 = _GEN_34121 | _GEN_22414; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22759 = _GEN_34122 | _GEN_22415; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22760 = _GEN_34123 | _GEN_22416; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22761 = _GEN_34124 | _GEN_22417; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22762 = _GEN_34125 | _GEN_22418; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22763 = _GEN_34126 | _GEN_22419; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22764 = _GEN_34127 | _GEN_22420; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22765 = _GEN_34128 | _GEN_22421; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22766 = _T_1486 ? _GEN_22758 : _GEN_22414; // @[sequencer-master.scala 168:32]
  wire  _GEN_22767 = _T_1486 ? _GEN_22759 : _GEN_22415; // @[sequencer-master.scala 168:32]
  wire  _GEN_22768 = _T_1486 ? _GEN_22760 : _GEN_22416; // @[sequencer-master.scala 168:32]
  wire  _GEN_22769 = _T_1486 ? _GEN_22761 : _GEN_22417; // @[sequencer-master.scala 168:32]
  wire  _GEN_22770 = _T_1486 ? _GEN_22762 : _GEN_22418; // @[sequencer-master.scala 168:32]
  wire  _GEN_22771 = _T_1486 ? _GEN_22763 : _GEN_22419; // @[sequencer-master.scala 168:32]
  wire  _GEN_22772 = _T_1486 ? _GEN_22764 : _GEN_22420; // @[sequencer-master.scala 168:32]
  wire  _GEN_22773 = _T_1486 ? _GEN_22765 : _GEN_22421; // @[sequencer-master.scala 168:32]
  wire  _GEN_22774 = _GEN_34121 | _GEN_22438; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22775 = _GEN_34122 | _GEN_22439; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22776 = _GEN_34123 | _GEN_22440; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22777 = _GEN_34124 | _GEN_22441; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22778 = _GEN_34125 | _GEN_22442; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22779 = _GEN_34126 | _GEN_22443; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22780 = _GEN_34127 | _GEN_22444; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22781 = _GEN_34128 | _GEN_22445; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22782 = _T_1508 ? _GEN_22774 : _GEN_22438; // @[sequencer-master.scala 168:32]
  wire  _GEN_22783 = _T_1508 ? _GEN_22775 : _GEN_22439; // @[sequencer-master.scala 168:32]
  wire  _GEN_22784 = _T_1508 ? _GEN_22776 : _GEN_22440; // @[sequencer-master.scala 168:32]
  wire  _GEN_22785 = _T_1508 ? _GEN_22777 : _GEN_22441; // @[sequencer-master.scala 168:32]
  wire  _GEN_22786 = _T_1508 ? _GEN_22778 : _GEN_22442; // @[sequencer-master.scala 168:32]
  wire  _GEN_22787 = _T_1508 ? _GEN_22779 : _GEN_22443; // @[sequencer-master.scala 168:32]
  wire  _GEN_22788 = _T_1508 ? _GEN_22780 : _GEN_22444; // @[sequencer-master.scala 168:32]
  wire  _GEN_22789 = _T_1508 ? _GEN_22781 : _GEN_22445; // @[sequencer-master.scala 168:32]
  wire  _GEN_22790 = _GEN_34121 | _GEN_22462; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22791 = _GEN_34122 | _GEN_22463; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22792 = _GEN_34123 | _GEN_22464; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22793 = _GEN_34124 | _GEN_22465; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22794 = _GEN_34125 | _GEN_22466; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22795 = _GEN_34126 | _GEN_22467; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22796 = _GEN_34127 | _GEN_22468; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22797 = _GEN_34128 | _GEN_22469; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22798 = _T_1530 ? _GEN_22790 : _GEN_22462; // @[sequencer-master.scala 168:32]
  wire  _GEN_22799 = _T_1530 ? _GEN_22791 : _GEN_22463; // @[sequencer-master.scala 168:32]
  wire  _GEN_22800 = _T_1530 ? _GEN_22792 : _GEN_22464; // @[sequencer-master.scala 168:32]
  wire  _GEN_22801 = _T_1530 ? _GEN_22793 : _GEN_22465; // @[sequencer-master.scala 168:32]
  wire  _GEN_22802 = _T_1530 ? _GEN_22794 : _GEN_22466; // @[sequencer-master.scala 168:32]
  wire  _GEN_22803 = _T_1530 ? _GEN_22795 : _GEN_22467; // @[sequencer-master.scala 168:32]
  wire  _GEN_22804 = _T_1530 ? _GEN_22796 : _GEN_22468; // @[sequencer-master.scala 168:32]
  wire  _GEN_22805 = _T_1530 ? _GEN_22797 : _GEN_22469; // @[sequencer-master.scala 168:32]
  wire  _GEN_22806 = _GEN_34121 | _GEN_22486; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22807 = _GEN_34122 | _GEN_22487; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22808 = _GEN_34123 | _GEN_22488; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22809 = _GEN_34124 | _GEN_22489; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22810 = _GEN_34125 | _GEN_22490; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22811 = _GEN_34126 | _GEN_22491; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22812 = _GEN_34127 | _GEN_22492; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22813 = _GEN_34128 | _GEN_22493; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22814 = _T_1552 ? _GEN_22806 : _GEN_22486; // @[sequencer-master.scala 168:32]
  wire  _GEN_22815 = _T_1552 ? _GEN_22807 : _GEN_22487; // @[sequencer-master.scala 168:32]
  wire  _GEN_22816 = _T_1552 ? _GEN_22808 : _GEN_22488; // @[sequencer-master.scala 168:32]
  wire  _GEN_22817 = _T_1552 ? _GEN_22809 : _GEN_22489; // @[sequencer-master.scala 168:32]
  wire  _GEN_22818 = _T_1552 ? _GEN_22810 : _GEN_22490; // @[sequencer-master.scala 168:32]
  wire  _GEN_22819 = _T_1552 ? _GEN_22811 : _GEN_22491; // @[sequencer-master.scala 168:32]
  wire  _GEN_22820 = _T_1552 ? _GEN_22812 : _GEN_22492; // @[sequencer-master.scala 168:32]
  wire  _GEN_22821 = _T_1552 ? _GEN_22813 : _GEN_22493; // @[sequencer-master.scala 168:32]
  wire  _GEN_22822 = _GEN_34121 | _GEN_22510; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22823 = _GEN_34122 | _GEN_22511; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22824 = _GEN_34123 | _GEN_22512; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22825 = _GEN_34124 | _GEN_22513; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22826 = _GEN_34125 | _GEN_22514; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22827 = _GEN_34126 | _GEN_22515; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22828 = _GEN_34127 | _GEN_22516; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22829 = _GEN_34128 | _GEN_22517; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22830 = _T_1574 ? _GEN_22822 : _GEN_22510; // @[sequencer-master.scala 168:32]
  wire  _GEN_22831 = _T_1574 ? _GEN_22823 : _GEN_22511; // @[sequencer-master.scala 168:32]
  wire  _GEN_22832 = _T_1574 ? _GEN_22824 : _GEN_22512; // @[sequencer-master.scala 168:32]
  wire  _GEN_22833 = _T_1574 ? _GEN_22825 : _GEN_22513; // @[sequencer-master.scala 168:32]
  wire  _GEN_22834 = _T_1574 ? _GEN_22826 : _GEN_22514; // @[sequencer-master.scala 168:32]
  wire  _GEN_22835 = _T_1574 ? _GEN_22827 : _GEN_22515; // @[sequencer-master.scala 168:32]
  wire  _GEN_22836 = _T_1574 ? _GEN_22828 : _GEN_22516; // @[sequencer-master.scala 168:32]
  wire  _GEN_22837 = _T_1574 ? _GEN_22829 : _GEN_22517; // @[sequencer-master.scala 168:32]
  wire  _GEN_22838 = _GEN_34121 | _GEN_22534; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22839 = _GEN_34122 | _GEN_22535; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22840 = _GEN_34123 | _GEN_22536; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22841 = _GEN_34124 | _GEN_22537; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22842 = _GEN_34125 | _GEN_22538; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22843 = _GEN_34126 | _GEN_22539; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22844 = _GEN_34127 | _GEN_22540; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22845 = _GEN_34128 | _GEN_22541; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_22846 = _T_1596 ? _GEN_22838 : _GEN_22534; // @[sequencer-master.scala 168:32]
  wire  _GEN_22847 = _T_1596 ? _GEN_22839 : _GEN_22535; // @[sequencer-master.scala 168:32]
  wire  _GEN_22848 = _T_1596 ? _GEN_22840 : _GEN_22536; // @[sequencer-master.scala 168:32]
  wire  _GEN_22849 = _T_1596 ? _GEN_22841 : _GEN_22537; // @[sequencer-master.scala 168:32]
  wire  _GEN_22850 = _T_1596 ? _GEN_22842 : _GEN_22538; // @[sequencer-master.scala 168:32]
  wire  _GEN_22851 = _T_1596 ? _GEN_22843 : _GEN_22539; // @[sequencer-master.scala 168:32]
  wire  _GEN_22852 = _T_1596 ? _GEN_22844 : _GEN_22540; // @[sequencer-master.scala 168:32]
  wire  _GEN_22853 = _T_1596 ? _GEN_22845 : _GEN_22541; // @[sequencer-master.scala 168:32]
  wire  _GEN_22854 = 3'h0 == _T_1647 | (3'h0 == _T_1645 | (_GEN_32729 | _GEN_21060)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22855 = 3'h1 == _T_1647 | (3'h1 == _T_1645 | (_GEN_32730 | _GEN_21061)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22856 = 3'h2 == _T_1647 | (3'h2 == _T_1645 | (_GEN_32731 | _GEN_21062)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22857 = 3'h3 == _T_1647 | (3'h3 == _T_1645 | (_GEN_32732 | _GEN_21063)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22858 = 3'h4 == _T_1647 | (3'h4 == _T_1645 | (_GEN_32733 | _GEN_21064)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22859 = 3'h5 == _T_1647 | (3'h5 == _T_1645 | (_GEN_32734 | _GEN_21065)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22860 = 3'h6 == _T_1647 | (3'h6 == _T_1645 | (_GEN_32735 | _GEN_21066)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22861 = 3'h7 == _T_1647 | (3'h7 == _T_1645 | (_GEN_32736 | _GEN_21067)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_22870 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22302; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22871 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22303; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22872 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22304; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22873 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22305; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22874 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22306; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22875 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22307; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22876 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22308; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22877 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22309; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_22878 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22310; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22879 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22311; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22880 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22312; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22881 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22313; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22882 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22314; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22883 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22315; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22884 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22316; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22885 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22317; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_22886 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22318; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22887 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22319; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22888 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22320; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22889 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22321; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22890 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22322; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22891 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22323; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22892 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22324; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22893 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22325; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_22894 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22326; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22895 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22327; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22896 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22328; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22897 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22329; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22898 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22330; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22899 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22331; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22900 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22332; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22901 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22333; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_22902 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22334; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22903 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22335; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22904 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22336; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22905 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22337; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22906 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22338; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22907 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22339; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22908 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22340; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22909 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22341; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_22910 = _GEN_36426 | (_GEN_34121 | (_GEN_32729 | _GEN_21116)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22911 = _GEN_36427 | (_GEN_34122 | (_GEN_32730 | _GEN_21117)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22912 = _GEN_36428 | (_GEN_34123 | (_GEN_32731 | _GEN_21118)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22913 = _GEN_36429 | (_GEN_34124 | (_GEN_32732 | _GEN_21119)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22914 = _GEN_36430 | (_GEN_34125 | (_GEN_32733 | _GEN_21120)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22915 = _GEN_36431 | (_GEN_34126 | (_GEN_32734 | _GEN_21121)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22916 = _GEN_36432 | (_GEN_34127 | (_GEN_32735 | _GEN_21122)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22917 = _GEN_36433 | (_GEN_34128 | (_GEN_32736 | _GEN_21123)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_22918 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22350; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22919 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22351; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22920 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22352; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22921 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22353; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22922 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22354; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22923 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22355; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22924 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22356; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22925 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22357; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22926 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22606; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22927 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22607; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22928 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22608; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22929 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22609; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22930 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22610; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22931 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22611; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22932 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22612; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22933 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22613; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22934 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22734; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22935 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22735; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22936 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22736; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22937 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22737; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22938 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22738; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22939 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22739; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22940 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22740; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22941 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22741; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22942 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22374; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22943 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22375; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22944 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22376; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22945 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22377; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22946 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22378; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22947 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22379; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22948 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22380; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22949 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22381; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22950 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22622; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22951 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22623; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22952 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22624; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22953 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22625; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22954 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22626; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22955 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22627; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22956 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22628; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22957 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22629; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22958 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22750; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22959 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22751; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22960 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22752; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22961 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22753; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22962 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22754; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22963 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22755; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22964 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22756; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22965 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22757; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22966 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22398; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22967 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22399; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22968 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22400; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22969 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22401; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22970 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22402; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22971 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22403; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22972 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22404; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22973 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22405; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22974 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22638; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22975 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22639; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22976 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22640; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22977 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22641; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22978 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22642; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22979 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22643; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22980 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22644; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22981 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22645; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22982 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22766; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22983 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22767; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22984 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22768; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22985 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22769; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22986 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22770; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22987 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22771; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22988 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22772; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22989 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22773; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_22990 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22422; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22991 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22423; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22992 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22424; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22993 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22425; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22994 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22426; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22995 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22427; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22996 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22428; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22997 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22429; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_22998 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22654; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_22999 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22655; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23000 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22656; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23001 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22657; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23002 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22658; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23003 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22659; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23004 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22660; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23005 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22661; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23006 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22782; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23007 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22783; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23008 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22784; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23009 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22785; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23010 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22786; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23011 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22787; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23012 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22788; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23013 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22789; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23014 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22446; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23015 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22447; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23016 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22448; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23017 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22449; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23018 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22450; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23019 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22451; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23020 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22452; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23021 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22453; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23022 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22670; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23023 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22671; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23024 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22672; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23025 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22673; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23026 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22674; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23027 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22675; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23028 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22676; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23029 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22677; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23030 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22798; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23031 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22799; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23032 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22800; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23033 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22801; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23034 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22802; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23035 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22803; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23036 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22804; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23037 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22805; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23038 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22470; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23039 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22471; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23040 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22472; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23041 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22473; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23042 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22474; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23043 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22475; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23044 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22476; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23045 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22477; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23046 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22686; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23047 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22687; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23048 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22688; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23049 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22689; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23050 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22690; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23051 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22691; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23052 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22692; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23053 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22693; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23054 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22814; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23055 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22815; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23056 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22816; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23057 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22817; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23058 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22818; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23059 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22819; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23060 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22820; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23061 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22821; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23062 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22494; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23063 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22495; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23064 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22496; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23065 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22497; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23066 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22498; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23067 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22499; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23068 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22500; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23069 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22501; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23070 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22702; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23071 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22703; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23072 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22704; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23073 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22705; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23074 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22706; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23075 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22707; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23076 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22708; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23077 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22709; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23078 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22830; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23079 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22831; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23080 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22832; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23081 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22833; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23082 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22834; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23083 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22835; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23084 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22836; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23085 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22837; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23086 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22518; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23087 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22519; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23088 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22520; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23089 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22521; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23090 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22522; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23091 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22523; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23092 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22524; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23093 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22525; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_23094 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22718; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23095 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22719; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23096 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22720; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23097 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22721; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23098 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22722; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23099 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22723; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23100 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22724; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23101 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22725; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_23102 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22846; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23103 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22847; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23104 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22848; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23105 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22849; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23106 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22850; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23107 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22851; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23108 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22852; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23109 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22853; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_23110 = 3'h0 == _T_1647 ? 1'h0 : _GEN_22542; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23111 = 3'h1 == _T_1647 ? 1'h0 : _GEN_22543; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23112 = 3'h2 == _T_1647 ? 1'h0 : _GEN_22544; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23113 = 3'h3 == _T_1647 ? 1'h0 : _GEN_22545; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23114 = 3'h4 == _T_1647 ? 1'h0 : _GEN_22546; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23115 = 3'h5 == _T_1647 ? 1'h0 : _GEN_22547; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23116 = 3'h6 == _T_1647 ? 1'h0 : _GEN_22548; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23117 = 3'h7 == _T_1647 ? 1'h0 : _GEN_22549; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_23126 = _GEN_36426 | _GEN_21468; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23127 = _GEN_36427 | _GEN_21469; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23128 = _GEN_36428 | _GEN_21470; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23129 = _GEN_36429 | _GEN_21471; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23130 = _GEN_36430 | _GEN_21472; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23131 = _GEN_36431 | _GEN_21473; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23132 = _GEN_36432 | _GEN_21474; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_23133 = _GEN_36433 | _GEN_21475; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_23134 = 3'h0 == _T_1647 ? io_op_bits_fn_union : _GEN_22566; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23135 = 3'h1 == _T_1647 ? io_op_bits_fn_union : _GEN_22567; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23136 = 3'h2 == _T_1647 ? io_op_bits_fn_union : _GEN_22568; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23137 = 3'h3 == _T_1647 ? io_op_bits_fn_union : _GEN_22569; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23138 = 3'h4 == _T_1647 ? io_op_bits_fn_union : _GEN_22570; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23139 = 3'h5 == _T_1647 ? io_op_bits_fn_union : _GEN_22571; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23140 = 3'h6 == _T_1647 ? io_op_bits_fn_union : _GEN_22572; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_23141 = 3'h7 == _T_1647 ? io_op_bits_fn_union : _GEN_22573; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [7:0] _GEN_23142 = 3'h0 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21476; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23143 = 3'h1 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21477; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23144 = 3'h2 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21478; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23145 = 3'h3 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21479; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23146 = 3'h4 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21480; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23147 = 3'h5 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21481; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23148 = 3'h6 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21482; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23149 = 3'h7 == _T_1647 ? io_op_bits_base_vd_id : _GEN_21483; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23150 = 3'h0 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22902; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23151 = 3'h1 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22903; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23152 = 3'h2 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22904; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23153 = 3'h3 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22905; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23154 = 3'h4 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22906; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23155 = 3'h5 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22907; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23156 = 3'h6 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22908; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23157 = 3'h7 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_22909; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23158 = 3'h0 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21484; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23159 = 3'h1 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21485; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23160 = 3'h2 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21486; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23161 = 3'h3 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21487; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23162 = 3'h4 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21488; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23163 = 3'h5 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21489; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23164 = 3'h6 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21490; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23165 = 3'h7 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_21491; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23166 = 3'h0 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21492; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23167 = 3'h1 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21493; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23168 = 3'h2 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21494; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23169 = 3'h3 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21495; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23170 = 3'h4 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21496; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23171 = 3'h5 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21497; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23172 = 3'h6 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21498; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_23173 = 3'h7 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_21499; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23174 = 3'h0 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21500; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23175 = 3'h1 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21501; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23176 = 3'h2 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21502; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23177 = 3'h3 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21503; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23178 = 3'h4 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21504; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23179 = 3'h5 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21505; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23180 = 3'h6 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21506; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [1:0] _GEN_23181 = 3'h7 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_21507; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_23182 = 3'h0 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21508; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23183 = 3'h1 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21509; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23184 = 3'h2 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21510; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23185 = 3'h3 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21511; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23186 = 3'h4 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21512; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23187 = 3'h5 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21513; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23188 = 3'h6 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21514; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23189 = 3'h7 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_21515; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_23190 = io_op_bits_base_vd_valid ? _GEN_23142 : _GEN_21476; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23191 = io_op_bits_base_vd_valid ? _GEN_23143 : _GEN_21477; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23192 = io_op_bits_base_vd_valid ? _GEN_23144 : _GEN_21478; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23193 = io_op_bits_base_vd_valid ? _GEN_23145 : _GEN_21479; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23194 = io_op_bits_base_vd_valid ? _GEN_23146 : _GEN_21480; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23195 = io_op_bits_base_vd_valid ? _GEN_23147 : _GEN_21481; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23196 = io_op_bits_base_vd_valid ? _GEN_23148 : _GEN_21482; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23197 = io_op_bits_base_vd_valid ? _GEN_23149 : _GEN_21483; // @[sequencer-master.scala 362:41]
  wire  _GEN_23198 = io_op_bits_base_vd_valid ? _GEN_23150 : _GEN_22902; // @[sequencer-master.scala 362:41]
  wire  _GEN_23199 = io_op_bits_base_vd_valid ? _GEN_23151 : _GEN_22903; // @[sequencer-master.scala 362:41]
  wire  _GEN_23200 = io_op_bits_base_vd_valid ? _GEN_23152 : _GEN_22904; // @[sequencer-master.scala 362:41]
  wire  _GEN_23201 = io_op_bits_base_vd_valid ? _GEN_23153 : _GEN_22905; // @[sequencer-master.scala 362:41]
  wire  _GEN_23202 = io_op_bits_base_vd_valid ? _GEN_23154 : _GEN_22906; // @[sequencer-master.scala 362:41]
  wire  _GEN_23203 = io_op_bits_base_vd_valid ? _GEN_23155 : _GEN_22907; // @[sequencer-master.scala 362:41]
  wire  _GEN_23204 = io_op_bits_base_vd_valid ? _GEN_23156 : _GEN_22908; // @[sequencer-master.scala 362:41]
  wire  _GEN_23205 = io_op_bits_base_vd_valid ? _GEN_23157 : _GEN_22909; // @[sequencer-master.scala 362:41]
  wire  _GEN_23206 = io_op_bits_base_vd_valid ? _GEN_23158 : _GEN_21484; // @[sequencer-master.scala 362:41]
  wire  _GEN_23207 = io_op_bits_base_vd_valid ? _GEN_23159 : _GEN_21485; // @[sequencer-master.scala 362:41]
  wire  _GEN_23208 = io_op_bits_base_vd_valid ? _GEN_23160 : _GEN_21486; // @[sequencer-master.scala 362:41]
  wire  _GEN_23209 = io_op_bits_base_vd_valid ? _GEN_23161 : _GEN_21487; // @[sequencer-master.scala 362:41]
  wire  _GEN_23210 = io_op_bits_base_vd_valid ? _GEN_23162 : _GEN_21488; // @[sequencer-master.scala 362:41]
  wire  _GEN_23211 = io_op_bits_base_vd_valid ? _GEN_23163 : _GEN_21489; // @[sequencer-master.scala 362:41]
  wire  _GEN_23212 = io_op_bits_base_vd_valid ? _GEN_23164 : _GEN_21490; // @[sequencer-master.scala 362:41]
  wire  _GEN_23213 = io_op_bits_base_vd_valid ? _GEN_23165 : _GEN_21491; // @[sequencer-master.scala 362:41]
  wire  _GEN_23214 = io_op_bits_base_vd_valid ? _GEN_23166 : _GEN_21492; // @[sequencer-master.scala 362:41]
  wire  _GEN_23215 = io_op_bits_base_vd_valid ? _GEN_23167 : _GEN_21493; // @[sequencer-master.scala 362:41]
  wire  _GEN_23216 = io_op_bits_base_vd_valid ? _GEN_23168 : _GEN_21494; // @[sequencer-master.scala 362:41]
  wire  _GEN_23217 = io_op_bits_base_vd_valid ? _GEN_23169 : _GEN_21495; // @[sequencer-master.scala 362:41]
  wire  _GEN_23218 = io_op_bits_base_vd_valid ? _GEN_23170 : _GEN_21496; // @[sequencer-master.scala 362:41]
  wire  _GEN_23219 = io_op_bits_base_vd_valid ? _GEN_23171 : _GEN_21497; // @[sequencer-master.scala 362:41]
  wire  _GEN_23220 = io_op_bits_base_vd_valid ? _GEN_23172 : _GEN_21498; // @[sequencer-master.scala 362:41]
  wire  _GEN_23221 = io_op_bits_base_vd_valid ? _GEN_23173 : _GEN_21499; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23222 = io_op_bits_base_vd_valid ? _GEN_23174 : _GEN_21500; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23223 = io_op_bits_base_vd_valid ? _GEN_23175 : _GEN_21501; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23224 = io_op_bits_base_vd_valid ? _GEN_23176 : _GEN_21502; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23225 = io_op_bits_base_vd_valid ? _GEN_23177 : _GEN_21503; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23226 = io_op_bits_base_vd_valid ? _GEN_23178 : _GEN_21504; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23227 = io_op_bits_base_vd_valid ? _GEN_23179 : _GEN_21505; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23228 = io_op_bits_base_vd_valid ? _GEN_23180 : _GEN_21506; // @[sequencer-master.scala 362:41]
  wire [1:0] _GEN_23229 = io_op_bits_base_vd_valid ? _GEN_23181 : _GEN_21507; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23230 = io_op_bits_base_vd_valid ? _GEN_23182 : _GEN_21508; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23231 = io_op_bits_base_vd_valid ? _GEN_23183 : _GEN_21509; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23232 = io_op_bits_base_vd_valid ? _GEN_23184 : _GEN_21510; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23233 = io_op_bits_base_vd_valid ? _GEN_23185 : _GEN_21511; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23234 = io_op_bits_base_vd_valid ? _GEN_23186 : _GEN_21512; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23235 = io_op_bits_base_vd_valid ? _GEN_23187 : _GEN_21513; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23236 = io_op_bits_base_vd_valid ? _GEN_23188 : _GEN_21514; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_23237 = io_op_bits_base_vd_valid ? _GEN_23189 : _GEN_21515; // @[sequencer-master.scala 362:41]
  wire  _GEN_23238 = _GEN_36426 | _GEN_22926; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23239 = _GEN_36427 | _GEN_22927; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23240 = _GEN_36428 | _GEN_22928; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23241 = _GEN_36429 | _GEN_22929; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23242 = _GEN_36430 | _GEN_22930; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23243 = _GEN_36431 | _GEN_22931; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23244 = _GEN_36432 | _GEN_22932; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23245 = _GEN_36433 | _GEN_22933; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23246 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23238 : _GEN_22926; // @[sequencer-master.scala 161:86]
  wire  _GEN_23247 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23239 : _GEN_22927; // @[sequencer-master.scala 161:86]
  wire  _GEN_23248 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23240 : _GEN_22928; // @[sequencer-master.scala 161:86]
  wire  _GEN_23249 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23241 : _GEN_22929; // @[sequencer-master.scala 161:86]
  wire  _GEN_23250 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23242 : _GEN_22930; // @[sequencer-master.scala 161:86]
  wire  _GEN_23251 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23243 : _GEN_22931; // @[sequencer-master.scala 161:86]
  wire  _GEN_23252 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23244 : _GEN_22932; // @[sequencer-master.scala 161:86]
  wire  _GEN_23253 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_23245 : _GEN_22933; // @[sequencer-master.scala 161:86]
  wire  _GEN_23254 = _GEN_36426 | _GEN_22950; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23255 = _GEN_36427 | _GEN_22951; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23256 = _GEN_36428 | _GEN_22952; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23257 = _GEN_36429 | _GEN_22953; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23258 = _GEN_36430 | _GEN_22954; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23259 = _GEN_36431 | _GEN_22955; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23260 = _GEN_36432 | _GEN_22956; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23261 = _GEN_36433 | _GEN_22957; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23262 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23254 : _GEN_22950; // @[sequencer-master.scala 161:86]
  wire  _GEN_23263 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23255 : _GEN_22951; // @[sequencer-master.scala 161:86]
  wire  _GEN_23264 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23256 : _GEN_22952; // @[sequencer-master.scala 161:86]
  wire  _GEN_23265 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23257 : _GEN_22953; // @[sequencer-master.scala 161:86]
  wire  _GEN_23266 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23258 : _GEN_22954; // @[sequencer-master.scala 161:86]
  wire  _GEN_23267 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23259 : _GEN_22955; // @[sequencer-master.scala 161:86]
  wire  _GEN_23268 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23260 : _GEN_22956; // @[sequencer-master.scala 161:86]
  wire  _GEN_23269 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_23261 : _GEN_22957; // @[sequencer-master.scala 161:86]
  wire  _GEN_23270 = _GEN_36426 | _GEN_22974; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23271 = _GEN_36427 | _GEN_22975; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23272 = _GEN_36428 | _GEN_22976; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23273 = _GEN_36429 | _GEN_22977; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23274 = _GEN_36430 | _GEN_22978; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23275 = _GEN_36431 | _GEN_22979; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23276 = _GEN_36432 | _GEN_22980; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23277 = _GEN_36433 | _GEN_22981; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23278 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23270 : _GEN_22974; // @[sequencer-master.scala 161:86]
  wire  _GEN_23279 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23271 : _GEN_22975; // @[sequencer-master.scala 161:86]
  wire  _GEN_23280 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23272 : _GEN_22976; // @[sequencer-master.scala 161:86]
  wire  _GEN_23281 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23273 : _GEN_22977; // @[sequencer-master.scala 161:86]
  wire  _GEN_23282 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23274 : _GEN_22978; // @[sequencer-master.scala 161:86]
  wire  _GEN_23283 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23275 : _GEN_22979; // @[sequencer-master.scala 161:86]
  wire  _GEN_23284 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23276 : _GEN_22980; // @[sequencer-master.scala 161:86]
  wire  _GEN_23285 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_23277 : _GEN_22981; // @[sequencer-master.scala 161:86]
  wire  _GEN_23286 = _GEN_36426 | _GEN_22998; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23287 = _GEN_36427 | _GEN_22999; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23288 = _GEN_36428 | _GEN_23000; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23289 = _GEN_36429 | _GEN_23001; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23290 = _GEN_36430 | _GEN_23002; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23291 = _GEN_36431 | _GEN_23003; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23292 = _GEN_36432 | _GEN_23004; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23293 = _GEN_36433 | _GEN_23005; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23294 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23286 : _GEN_22998; // @[sequencer-master.scala 161:86]
  wire  _GEN_23295 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23287 : _GEN_22999; // @[sequencer-master.scala 161:86]
  wire  _GEN_23296 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23288 : _GEN_23000; // @[sequencer-master.scala 161:86]
  wire  _GEN_23297 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23289 : _GEN_23001; // @[sequencer-master.scala 161:86]
  wire  _GEN_23298 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23290 : _GEN_23002; // @[sequencer-master.scala 161:86]
  wire  _GEN_23299 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23291 : _GEN_23003; // @[sequencer-master.scala 161:86]
  wire  _GEN_23300 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23292 : _GEN_23004; // @[sequencer-master.scala 161:86]
  wire  _GEN_23301 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_23293 : _GEN_23005; // @[sequencer-master.scala 161:86]
  wire  _GEN_23302 = _GEN_36426 | _GEN_23022; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23303 = _GEN_36427 | _GEN_23023; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23304 = _GEN_36428 | _GEN_23024; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23305 = _GEN_36429 | _GEN_23025; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23306 = _GEN_36430 | _GEN_23026; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23307 = _GEN_36431 | _GEN_23027; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23308 = _GEN_36432 | _GEN_23028; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23309 = _GEN_36433 | _GEN_23029; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23310 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23302 : _GEN_23022; // @[sequencer-master.scala 161:86]
  wire  _GEN_23311 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23303 : _GEN_23023; // @[sequencer-master.scala 161:86]
  wire  _GEN_23312 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23304 : _GEN_23024; // @[sequencer-master.scala 161:86]
  wire  _GEN_23313 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23305 : _GEN_23025; // @[sequencer-master.scala 161:86]
  wire  _GEN_23314 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23306 : _GEN_23026; // @[sequencer-master.scala 161:86]
  wire  _GEN_23315 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23307 : _GEN_23027; // @[sequencer-master.scala 161:86]
  wire  _GEN_23316 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23308 : _GEN_23028; // @[sequencer-master.scala 161:86]
  wire  _GEN_23317 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_23309 : _GEN_23029; // @[sequencer-master.scala 161:86]
  wire  _GEN_23318 = _GEN_36426 | _GEN_23046; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23319 = _GEN_36427 | _GEN_23047; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23320 = _GEN_36428 | _GEN_23048; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23321 = _GEN_36429 | _GEN_23049; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23322 = _GEN_36430 | _GEN_23050; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23323 = _GEN_36431 | _GEN_23051; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23324 = _GEN_36432 | _GEN_23052; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23325 = _GEN_36433 | _GEN_23053; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23326 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23318 : _GEN_23046; // @[sequencer-master.scala 161:86]
  wire  _GEN_23327 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23319 : _GEN_23047; // @[sequencer-master.scala 161:86]
  wire  _GEN_23328 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23320 : _GEN_23048; // @[sequencer-master.scala 161:86]
  wire  _GEN_23329 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23321 : _GEN_23049; // @[sequencer-master.scala 161:86]
  wire  _GEN_23330 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23322 : _GEN_23050; // @[sequencer-master.scala 161:86]
  wire  _GEN_23331 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23323 : _GEN_23051; // @[sequencer-master.scala 161:86]
  wire  _GEN_23332 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23324 : _GEN_23052; // @[sequencer-master.scala 161:86]
  wire  _GEN_23333 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_23325 : _GEN_23053; // @[sequencer-master.scala 161:86]
  wire  _GEN_23334 = _GEN_36426 | _GEN_23070; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23335 = _GEN_36427 | _GEN_23071; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23336 = _GEN_36428 | _GEN_23072; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23337 = _GEN_36429 | _GEN_23073; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23338 = _GEN_36430 | _GEN_23074; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23339 = _GEN_36431 | _GEN_23075; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23340 = _GEN_36432 | _GEN_23076; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23341 = _GEN_36433 | _GEN_23077; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23342 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23334 : _GEN_23070; // @[sequencer-master.scala 161:86]
  wire  _GEN_23343 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23335 : _GEN_23071; // @[sequencer-master.scala 161:86]
  wire  _GEN_23344 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23336 : _GEN_23072; // @[sequencer-master.scala 161:86]
  wire  _GEN_23345 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23337 : _GEN_23073; // @[sequencer-master.scala 161:86]
  wire  _GEN_23346 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23338 : _GEN_23074; // @[sequencer-master.scala 161:86]
  wire  _GEN_23347 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23339 : _GEN_23075; // @[sequencer-master.scala 161:86]
  wire  _GEN_23348 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23340 : _GEN_23076; // @[sequencer-master.scala 161:86]
  wire  _GEN_23349 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_23341 : _GEN_23077; // @[sequencer-master.scala 161:86]
  wire  _GEN_23350 = _GEN_36426 | _GEN_23094; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23351 = _GEN_36427 | _GEN_23095; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23352 = _GEN_36428 | _GEN_23096; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23353 = _GEN_36429 | _GEN_23097; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23354 = _GEN_36430 | _GEN_23098; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23355 = _GEN_36431 | _GEN_23099; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23356 = _GEN_36432 | _GEN_23100; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23357 = _GEN_36433 | _GEN_23101; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_23358 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23350 : _GEN_23094; // @[sequencer-master.scala 161:86]
  wire  _GEN_23359 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23351 : _GEN_23095; // @[sequencer-master.scala 161:86]
  wire  _GEN_23360 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23352 : _GEN_23096; // @[sequencer-master.scala 161:86]
  wire  _GEN_23361 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23353 : _GEN_23097; // @[sequencer-master.scala 161:86]
  wire  _GEN_23362 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23354 : _GEN_23098; // @[sequencer-master.scala 161:86]
  wire  _GEN_23363 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23355 : _GEN_23099; // @[sequencer-master.scala 161:86]
  wire  _GEN_23364 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23356 : _GEN_23100; // @[sequencer-master.scala 161:86]
  wire  _GEN_23365 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_23357 : _GEN_23101; // @[sequencer-master.scala 161:86]
  wire  _GEN_23366 = _GEN_36426 | _GEN_22934; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23367 = _GEN_36427 | _GEN_22935; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23368 = _GEN_36428 | _GEN_22936; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23369 = _GEN_36429 | _GEN_22937; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23370 = _GEN_36430 | _GEN_22938; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23371 = _GEN_36431 | _GEN_22939; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23372 = _GEN_36432 | _GEN_22940; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23373 = _GEN_36433 | _GEN_22941; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23374 = _T_1442 ? _GEN_23366 : _GEN_22934; // @[sequencer-master.scala 168:32]
  wire  _GEN_23375 = _T_1442 ? _GEN_23367 : _GEN_22935; // @[sequencer-master.scala 168:32]
  wire  _GEN_23376 = _T_1442 ? _GEN_23368 : _GEN_22936; // @[sequencer-master.scala 168:32]
  wire  _GEN_23377 = _T_1442 ? _GEN_23369 : _GEN_22937; // @[sequencer-master.scala 168:32]
  wire  _GEN_23378 = _T_1442 ? _GEN_23370 : _GEN_22938; // @[sequencer-master.scala 168:32]
  wire  _GEN_23379 = _T_1442 ? _GEN_23371 : _GEN_22939; // @[sequencer-master.scala 168:32]
  wire  _GEN_23380 = _T_1442 ? _GEN_23372 : _GEN_22940; // @[sequencer-master.scala 168:32]
  wire  _GEN_23381 = _T_1442 ? _GEN_23373 : _GEN_22941; // @[sequencer-master.scala 168:32]
  wire  _GEN_23382 = _GEN_36426 | _GEN_22958; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23383 = _GEN_36427 | _GEN_22959; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23384 = _GEN_36428 | _GEN_22960; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23385 = _GEN_36429 | _GEN_22961; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23386 = _GEN_36430 | _GEN_22962; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23387 = _GEN_36431 | _GEN_22963; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23388 = _GEN_36432 | _GEN_22964; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23389 = _GEN_36433 | _GEN_22965; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23390 = _T_1464 ? _GEN_23382 : _GEN_22958; // @[sequencer-master.scala 168:32]
  wire  _GEN_23391 = _T_1464 ? _GEN_23383 : _GEN_22959; // @[sequencer-master.scala 168:32]
  wire  _GEN_23392 = _T_1464 ? _GEN_23384 : _GEN_22960; // @[sequencer-master.scala 168:32]
  wire  _GEN_23393 = _T_1464 ? _GEN_23385 : _GEN_22961; // @[sequencer-master.scala 168:32]
  wire  _GEN_23394 = _T_1464 ? _GEN_23386 : _GEN_22962; // @[sequencer-master.scala 168:32]
  wire  _GEN_23395 = _T_1464 ? _GEN_23387 : _GEN_22963; // @[sequencer-master.scala 168:32]
  wire  _GEN_23396 = _T_1464 ? _GEN_23388 : _GEN_22964; // @[sequencer-master.scala 168:32]
  wire  _GEN_23397 = _T_1464 ? _GEN_23389 : _GEN_22965; // @[sequencer-master.scala 168:32]
  wire  _GEN_23398 = _GEN_36426 | _GEN_22982; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23399 = _GEN_36427 | _GEN_22983; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23400 = _GEN_36428 | _GEN_22984; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23401 = _GEN_36429 | _GEN_22985; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23402 = _GEN_36430 | _GEN_22986; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23403 = _GEN_36431 | _GEN_22987; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23404 = _GEN_36432 | _GEN_22988; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23405 = _GEN_36433 | _GEN_22989; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23406 = _T_1486 ? _GEN_23398 : _GEN_22982; // @[sequencer-master.scala 168:32]
  wire  _GEN_23407 = _T_1486 ? _GEN_23399 : _GEN_22983; // @[sequencer-master.scala 168:32]
  wire  _GEN_23408 = _T_1486 ? _GEN_23400 : _GEN_22984; // @[sequencer-master.scala 168:32]
  wire  _GEN_23409 = _T_1486 ? _GEN_23401 : _GEN_22985; // @[sequencer-master.scala 168:32]
  wire  _GEN_23410 = _T_1486 ? _GEN_23402 : _GEN_22986; // @[sequencer-master.scala 168:32]
  wire  _GEN_23411 = _T_1486 ? _GEN_23403 : _GEN_22987; // @[sequencer-master.scala 168:32]
  wire  _GEN_23412 = _T_1486 ? _GEN_23404 : _GEN_22988; // @[sequencer-master.scala 168:32]
  wire  _GEN_23413 = _T_1486 ? _GEN_23405 : _GEN_22989; // @[sequencer-master.scala 168:32]
  wire  _GEN_23414 = _GEN_36426 | _GEN_23006; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23415 = _GEN_36427 | _GEN_23007; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23416 = _GEN_36428 | _GEN_23008; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23417 = _GEN_36429 | _GEN_23009; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23418 = _GEN_36430 | _GEN_23010; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23419 = _GEN_36431 | _GEN_23011; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23420 = _GEN_36432 | _GEN_23012; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23421 = _GEN_36433 | _GEN_23013; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23422 = _T_1508 ? _GEN_23414 : _GEN_23006; // @[sequencer-master.scala 168:32]
  wire  _GEN_23423 = _T_1508 ? _GEN_23415 : _GEN_23007; // @[sequencer-master.scala 168:32]
  wire  _GEN_23424 = _T_1508 ? _GEN_23416 : _GEN_23008; // @[sequencer-master.scala 168:32]
  wire  _GEN_23425 = _T_1508 ? _GEN_23417 : _GEN_23009; // @[sequencer-master.scala 168:32]
  wire  _GEN_23426 = _T_1508 ? _GEN_23418 : _GEN_23010; // @[sequencer-master.scala 168:32]
  wire  _GEN_23427 = _T_1508 ? _GEN_23419 : _GEN_23011; // @[sequencer-master.scala 168:32]
  wire  _GEN_23428 = _T_1508 ? _GEN_23420 : _GEN_23012; // @[sequencer-master.scala 168:32]
  wire  _GEN_23429 = _T_1508 ? _GEN_23421 : _GEN_23013; // @[sequencer-master.scala 168:32]
  wire  _GEN_23430 = _GEN_36426 | _GEN_23030; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23431 = _GEN_36427 | _GEN_23031; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23432 = _GEN_36428 | _GEN_23032; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23433 = _GEN_36429 | _GEN_23033; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23434 = _GEN_36430 | _GEN_23034; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23435 = _GEN_36431 | _GEN_23035; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23436 = _GEN_36432 | _GEN_23036; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23437 = _GEN_36433 | _GEN_23037; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23438 = _T_1530 ? _GEN_23430 : _GEN_23030; // @[sequencer-master.scala 168:32]
  wire  _GEN_23439 = _T_1530 ? _GEN_23431 : _GEN_23031; // @[sequencer-master.scala 168:32]
  wire  _GEN_23440 = _T_1530 ? _GEN_23432 : _GEN_23032; // @[sequencer-master.scala 168:32]
  wire  _GEN_23441 = _T_1530 ? _GEN_23433 : _GEN_23033; // @[sequencer-master.scala 168:32]
  wire  _GEN_23442 = _T_1530 ? _GEN_23434 : _GEN_23034; // @[sequencer-master.scala 168:32]
  wire  _GEN_23443 = _T_1530 ? _GEN_23435 : _GEN_23035; // @[sequencer-master.scala 168:32]
  wire  _GEN_23444 = _T_1530 ? _GEN_23436 : _GEN_23036; // @[sequencer-master.scala 168:32]
  wire  _GEN_23445 = _T_1530 ? _GEN_23437 : _GEN_23037; // @[sequencer-master.scala 168:32]
  wire  _GEN_23446 = _GEN_36426 | _GEN_23054; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23447 = _GEN_36427 | _GEN_23055; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23448 = _GEN_36428 | _GEN_23056; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23449 = _GEN_36429 | _GEN_23057; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23450 = _GEN_36430 | _GEN_23058; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23451 = _GEN_36431 | _GEN_23059; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23452 = _GEN_36432 | _GEN_23060; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23453 = _GEN_36433 | _GEN_23061; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23454 = _T_1552 ? _GEN_23446 : _GEN_23054; // @[sequencer-master.scala 168:32]
  wire  _GEN_23455 = _T_1552 ? _GEN_23447 : _GEN_23055; // @[sequencer-master.scala 168:32]
  wire  _GEN_23456 = _T_1552 ? _GEN_23448 : _GEN_23056; // @[sequencer-master.scala 168:32]
  wire  _GEN_23457 = _T_1552 ? _GEN_23449 : _GEN_23057; // @[sequencer-master.scala 168:32]
  wire  _GEN_23458 = _T_1552 ? _GEN_23450 : _GEN_23058; // @[sequencer-master.scala 168:32]
  wire  _GEN_23459 = _T_1552 ? _GEN_23451 : _GEN_23059; // @[sequencer-master.scala 168:32]
  wire  _GEN_23460 = _T_1552 ? _GEN_23452 : _GEN_23060; // @[sequencer-master.scala 168:32]
  wire  _GEN_23461 = _T_1552 ? _GEN_23453 : _GEN_23061; // @[sequencer-master.scala 168:32]
  wire  _GEN_23462 = _GEN_36426 | _GEN_23078; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23463 = _GEN_36427 | _GEN_23079; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23464 = _GEN_36428 | _GEN_23080; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23465 = _GEN_36429 | _GEN_23081; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23466 = _GEN_36430 | _GEN_23082; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23467 = _GEN_36431 | _GEN_23083; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23468 = _GEN_36432 | _GEN_23084; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23469 = _GEN_36433 | _GEN_23085; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23470 = _T_1574 ? _GEN_23462 : _GEN_23078; // @[sequencer-master.scala 168:32]
  wire  _GEN_23471 = _T_1574 ? _GEN_23463 : _GEN_23079; // @[sequencer-master.scala 168:32]
  wire  _GEN_23472 = _T_1574 ? _GEN_23464 : _GEN_23080; // @[sequencer-master.scala 168:32]
  wire  _GEN_23473 = _T_1574 ? _GEN_23465 : _GEN_23081; // @[sequencer-master.scala 168:32]
  wire  _GEN_23474 = _T_1574 ? _GEN_23466 : _GEN_23082; // @[sequencer-master.scala 168:32]
  wire  _GEN_23475 = _T_1574 ? _GEN_23467 : _GEN_23083; // @[sequencer-master.scala 168:32]
  wire  _GEN_23476 = _T_1574 ? _GEN_23468 : _GEN_23084; // @[sequencer-master.scala 168:32]
  wire  _GEN_23477 = _T_1574 ? _GEN_23469 : _GEN_23085; // @[sequencer-master.scala 168:32]
  wire  _GEN_23478 = _GEN_36426 | _GEN_23102; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23479 = _GEN_36427 | _GEN_23103; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23480 = _GEN_36428 | _GEN_23104; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23481 = _GEN_36429 | _GEN_23105; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23482 = _GEN_36430 | _GEN_23106; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23483 = _GEN_36431 | _GEN_23107; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23484 = _GEN_36432 | _GEN_23108; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23485 = _GEN_36433 | _GEN_23109; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_23486 = _T_1596 ? _GEN_23478 : _GEN_23102; // @[sequencer-master.scala 168:32]
  wire  _GEN_23487 = _T_1596 ? _GEN_23479 : _GEN_23103; // @[sequencer-master.scala 168:32]
  wire  _GEN_23488 = _T_1596 ? _GEN_23480 : _GEN_23104; // @[sequencer-master.scala 168:32]
  wire  _GEN_23489 = _T_1596 ? _GEN_23481 : _GEN_23105; // @[sequencer-master.scala 168:32]
  wire  _GEN_23490 = _T_1596 ? _GEN_23482 : _GEN_23106; // @[sequencer-master.scala 168:32]
  wire  _GEN_23491 = _T_1596 ? _GEN_23483 : _GEN_23107; // @[sequencer-master.scala 168:32]
  wire  _GEN_23492 = _T_1596 ? _GEN_23484 : _GEN_23108; // @[sequencer-master.scala 168:32]
  wire  _GEN_23493 = _T_1596 ? _GEN_23485 : _GEN_23109; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_23494 = 3'h0 == _T_1647 ? 2'h0 : _GEN_22574; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23495 = 3'h1 == _T_1647 ? 2'h0 : _GEN_22575; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23496 = 3'h2 == _T_1647 ? 2'h0 : _GEN_22576; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23497 = 3'h3 == _T_1647 ? 2'h0 : _GEN_22577; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23498 = 3'h4 == _T_1647 ? 2'h0 : _GEN_22578; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23499 = 3'h5 == _T_1647 ? 2'h0 : _GEN_22579; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23500 = 3'h6 == _T_1647 ? 2'h0 : _GEN_22580; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_23501 = 3'h7 == _T_1647 ? 2'h0 : _GEN_22581; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_23502 = 3'h0 == _T_1647 ? 4'h0 : _GEN_22582; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23503 = 3'h1 == _T_1647 ? 4'h0 : _GEN_22583; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23504 = 3'h2 == _T_1647 ? 4'h0 : _GEN_22584; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23505 = 3'h3 == _T_1647 ? 4'h0 : _GEN_22585; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23506 = 3'h4 == _T_1647 ? 4'h0 : _GEN_22586; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23507 = 3'h5 == _T_1647 ? 4'h0 : _GEN_22587; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23508 = 3'h6 == _T_1647 ? 4'h0 : _GEN_22588; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_23509 = 3'h7 == _T_1647 ? 4'h0 : _GEN_22589; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_23510 = 3'h0 == _T_1647 ? 3'h0 : _GEN_22590; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23511 = 3'h1 == _T_1647 ? 3'h0 : _GEN_22591; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23512 = 3'h2 == _T_1647 ? 3'h0 : _GEN_22592; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23513 = 3'h3 == _T_1647 ? 3'h0 : _GEN_22593; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23514 = 3'h4 == _T_1647 ? 3'h0 : _GEN_22594; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23515 = 3'h5 == _T_1647 ? 3'h0 : _GEN_22595; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23516 = 3'h6 == _T_1647 ? 3'h0 : _GEN_22596; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_23517 = 3'h7 == _T_1647 ? 3'h0 : _GEN_22597; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_23518 = io_op_bits_active_vldx ? _GEN_22854 : _GEN_21060; // @[sequencer-master.scala 651:39]
  wire  _GEN_23519 = io_op_bits_active_vldx ? _GEN_22855 : _GEN_21061; // @[sequencer-master.scala 651:39]
  wire  _GEN_23520 = io_op_bits_active_vldx ? _GEN_22856 : _GEN_21062; // @[sequencer-master.scala 651:39]
  wire  _GEN_23521 = io_op_bits_active_vldx ? _GEN_22857 : _GEN_21063; // @[sequencer-master.scala 651:39]
  wire  _GEN_23522 = io_op_bits_active_vldx ? _GEN_22858 : _GEN_21064; // @[sequencer-master.scala 651:39]
  wire  _GEN_23523 = io_op_bits_active_vldx ? _GEN_22859 : _GEN_21065; // @[sequencer-master.scala 651:39]
  wire  _GEN_23524 = io_op_bits_active_vldx ? _GEN_22860 : _GEN_21066; // @[sequencer-master.scala 651:39]
  wire  _GEN_23525 = io_op_bits_active_vldx ? _GEN_22861 : _GEN_21067; // @[sequencer-master.scala 651:39]
  wire  _GEN_23534 = io_op_bits_active_vldx ? _GEN_22870 : _GEN_21076; // @[sequencer-master.scala 651:39]
  wire  _GEN_23535 = io_op_bits_active_vldx ? _GEN_22871 : _GEN_21077; // @[sequencer-master.scala 651:39]
  wire  _GEN_23536 = io_op_bits_active_vldx ? _GEN_22872 : _GEN_21078; // @[sequencer-master.scala 651:39]
  wire  _GEN_23537 = io_op_bits_active_vldx ? _GEN_22873 : _GEN_21079; // @[sequencer-master.scala 651:39]
  wire  _GEN_23538 = io_op_bits_active_vldx ? _GEN_22874 : _GEN_21080; // @[sequencer-master.scala 651:39]
  wire  _GEN_23539 = io_op_bits_active_vldx ? _GEN_22875 : _GEN_21081; // @[sequencer-master.scala 651:39]
  wire  _GEN_23540 = io_op_bits_active_vldx ? _GEN_22876 : _GEN_21082; // @[sequencer-master.scala 651:39]
  wire  _GEN_23541 = io_op_bits_active_vldx ? _GEN_22877 : _GEN_21083; // @[sequencer-master.scala 651:39]
  wire  _GEN_23542 = io_op_bits_active_vldx ? _GEN_22878 : _GEN_21084; // @[sequencer-master.scala 651:39]
  wire  _GEN_23543 = io_op_bits_active_vldx ? _GEN_22879 : _GEN_21085; // @[sequencer-master.scala 651:39]
  wire  _GEN_23544 = io_op_bits_active_vldx ? _GEN_22880 : _GEN_21086; // @[sequencer-master.scala 651:39]
  wire  _GEN_23545 = io_op_bits_active_vldx ? _GEN_22881 : _GEN_21087; // @[sequencer-master.scala 651:39]
  wire  _GEN_23546 = io_op_bits_active_vldx ? _GEN_22882 : _GEN_21088; // @[sequencer-master.scala 651:39]
  wire  _GEN_23547 = io_op_bits_active_vldx ? _GEN_22883 : _GEN_21089; // @[sequencer-master.scala 651:39]
  wire  _GEN_23548 = io_op_bits_active_vldx ? _GEN_22884 : _GEN_21090; // @[sequencer-master.scala 651:39]
  wire  _GEN_23549 = io_op_bits_active_vldx ? _GEN_22885 : _GEN_21091; // @[sequencer-master.scala 651:39]
  wire  _GEN_23550 = io_op_bits_active_vldx ? _GEN_22886 : _GEN_21092; // @[sequencer-master.scala 651:39]
  wire  _GEN_23551 = io_op_bits_active_vldx ? _GEN_22887 : _GEN_21093; // @[sequencer-master.scala 651:39]
  wire  _GEN_23552 = io_op_bits_active_vldx ? _GEN_22888 : _GEN_21094; // @[sequencer-master.scala 651:39]
  wire  _GEN_23553 = io_op_bits_active_vldx ? _GEN_22889 : _GEN_21095; // @[sequencer-master.scala 651:39]
  wire  _GEN_23554 = io_op_bits_active_vldx ? _GEN_22890 : _GEN_21096; // @[sequencer-master.scala 651:39]
  wire  _GEN_23555 = io_op_bits_active_vldx ? _GEN_22891 : _GEN_21097; // @[sequencer-master.scala 651:39]
  wire  _GEN_23556 = io_op_bits_active_vldx ? _GEN_22892 : _GEN_21098; // @[sequencer-master.scala 651:39]
  wire  _GEN_23557 = io_op_bits_active_vldx ? _GEN_22893 : _GEN_21099; // @[sequencer-master.scala 651:39]
  wire  _GEN_23558 = io_op_bits_active_vldx ? _GEN_22894 : _GEN_21100; // @[sequencer-master.scala 651:39]
  wire  _GEN_23559 = io_op_bits_active_vldx ? _GEN_22895 : _GEN_21101; // @[sequencer-master.scala 651:39]
  wire  _GEN_23560 = io_op_bits_active_vldx ? _GEN_22896 : _GEN_21102; // @[sequencer-master.scala 651:39]
  wire  _GEN_23561 = io_op_bits_active_vldx ? _GEN_22897 : _GEN_21103; // @[sequencer-master.scala 651:39]
  wire  _GEN_23562 = io_op_bits_active_vldx ? _GEN_22898 : _GEN_21104; // @[sequencer-master.scala 651:39]
  wire  _GEN_23563 = io_op_bits_active_vldx ? _GEN_22899 : _GEN_21105; // @[sequencer-master.scala 651:39]
  wire  _GEN_23564 = io_op_bits_active_vldx ? _GEN_22900 : _GEN_21106; // @[sequencer-master.scala 651:39]
  wire  _GEN_23565 = io_op_bits_active_vldx ? _GEN_22901 : _GEN_21107; // @[sequencer-master.scala 651:39]
  wire  _GEN_23566 = io_op_bits_active_vldx ? _GEN_23198 : _GEN_21108; // @[sequencer-master.scala 651:39]
  wire  _GEN_23567 = io_op_bits_active_vldx ? _GEN_23199 : _GEN_21109; // @[sequencer-master.scala 651:39]
  wire  _GEN_23568 = io_op_bits_active_vldx ? _GEN_23200 : _GEN_21110; // @[sequencer-master.scala 651:39]
  wire  _GEN_23569 = io_op_bits_active_vldx ? _GEN_23201 : _GEN_21111; // @[sequencer-master.scala 651:39]
  wire  _GEN_23570 = io_op_bits_active_vldx ? _GEN_23202 : _GEN_21112; // @[sequencer-master.scala 651:39]
  wire  _GEN_23571 = io_op_bits_active_vldx ? _GEN_23203 : _GEN_21113; // @[sequencer-master.scala 651:39]
  wire  _GEN_23572 = io_op_bits_active_vldx ? _GEN_23204 : _GEN_21114; // @[sequencer-master.scala 651:39]
  wire  _GEN_23573 = io_op_bits_active_vldx ? _GEN_23205 : _GEN_21115; // @[sequencer-master.scala 651:39]
  wire  _GEN_23574 = io_op_bits_active_vldx ? _GEN_22910 : _GEN_21116; // @[sequencer-master.scala 651:39]
  wire  _GEN_23575 = io_op_bits_active_vldx ? _GEN_22911 : _GEN_21117; // @[sequencer-master.scala 651:39]
  wire  _GEN_23576 = io_op_bits_active_vldx ? _GEN_22912 : _GEN_21118; // @[sequencer-master.scala 651:39]
  wire  _GEN_23577 = io_op_bits_active_vldx ? _GEN_22913 : _GEN_21119; // @[sequencer-master.scala 651:39]
  wire  _GEN_23578 = io_op_bits_active_vldx ? _GEN_22914 : _GEN_21120; // @[sequencer-master.scala 651:39]
  wire  _GEN_23579 = io_op_bits_active_vldx ? _GEN_22915 : _GEN_21121; // @[sequencer-master.scala 651:39]
  wire  _GEN_23580 = io_op_bits_active_vldx ? _GEN_22916 : _GEN_21122; // @[sequencer-master.scala 651:39]
  wire  _GEN_23581 = io_op_bits_active_vldx ? _GEN_22917 : _GEN_21123; // @[sequencer-master.scala 651:39]
  wire  _GEN_23582 = io_op_bits_active_vldx ? _GEN_22918 : _GEN_21124; // @[sequencer-master.scala 651:39]
  wire  _GEN_23583 = io_op_bits_active_vldx ? _GEN_22919 : _GEN_21125; // @[sequencer-master.scala 651:39]
  wire  _GEN_23584 = io_op_bits_active_vldx ? _GEN_22920 : _GEN_21126; // @[sequencer-master.scala 651:39]
  wire  _GEN_23585 = io_op_bits_active_vldx ? _GEN_22921 : _GEN_21127; // @[sequencer-master.scala 651:39]
  wire  _GEN_23586 = io_op_bits_active_vldx ? _GEN_22922 : _GEN_21128; // @[sequencer-master.scala 651:39]
  wire  _GEN_23587 = io_op_bits_active_vldx ? _GEN_22923 : _GEN_21129; // @[sequencer-master.scala 651:39]
  wire  _GEN_23588 = io_op_bits_active_vldx ? _GEN_22924 : _GEN_21130; // @[sequencer-master.scala 651:39]
  wire  _GEN_23589 = io_op_bits_active_vldx ? _GEN_22925 : _GEN_21131; // @[sequencer-master.scala 651:39]
  wire  _GEN_23590 = io_op_bits_active_vldx ? _GEN_23246 : _GEN_21132; // @[sequencer-master.scala 651:39]
  wire  _GEN_23591 = io_op_bits_active_vldx ? _GEN_23247 : _GEN_21133; // @[sequencer-master.scala 651:39]
  wire  _GEN_23592 = io_op_bits_active_vldx ? _GEN_23248 : _GEN_21134; // @[sequencer-master.scala 651:39]
  wire  _GEN_23593 = io_op_bits_active_vldx ? _GEN_23249 : _GEN_21135; // @[sequencer-master.scala 651:39]
  wire  _GEN_23594 = io_op_bits_active_vldx ? _GEN_23250 : _GEN_21136; // @[sequencer-master.scala 651:39]
  wire  _GEN_23595 = io_op_bits_active_vldx ? _GEN_23251 : _GEN_21137; // @[sequencer-master.scala 651:39]
  wire  _GEN_23596 = io_op_bits_active_vldx ? _GEN_23252 : _GEN_21138; // @[sequencer-master.scala 651:39]
  wire  _GEN_23597 = io_op_bits_active_vldx ? _GEN_23253 : _GEN_21139; // @[sequencer-master.scala 651:39]
  wire  _GEN_23598 = io_op_bits_active_vldx ? _GEN_23374 : _GEN_21140; // @[sequencer-master.scala 651:39]
  wire  _GEN_23599 = io_op_bits_active_vldx ? _GEN_23375 : _GEN_21141; // @[sequencer-master.scala 651:39]
  wire  _GEN_23600 = io_op_bits_active_vldx ? _GEN_23376 : _GEN_21142; // @[sequencer-master.scala 651:39]
  wire  _GEN_23601 = io_op_bits_active_vldx ? _GEN_23377 : _GEN_21143; // @[sequencer-master.scala 651:39]
  wire  _GEN_23602 = io_op_bits_active_vldx ? _GEN_23378 : _GEN_21144; // @[sequencer-master.scala 651:39]
  wire  _GEN_23603 = io_op_bits_active_vldx ? _GEN_23379 : _GEN_21145; // @[sequencer-master.scala 651:39]
  wire  _GEN_23604 = io_op_bits_active_vldx ? _GEN_23380 : _GEN_21146; // @[sequencer-master.scala 651:39]
  wire  _GEN_23605 = io_op_bits_active_vldx ? _GEN_23381 : _GEN_21147; // @[sequencer-master.scala 651:39]
  wire  _GEN_23606 = io_op_bits_active_vldx ? _GEN_22942 : _GEN_21148; // @[sequencer-master.scala 651:39]
  wire  _GEN_23607 = io_op_bits_active_vldx ? _GEN_22943 : _GEN_21149; // @[sequencer-master.scala 651:39]
  wire  _GEN_23608 = io_op_bits_active_vldx ? _GEN_22944 : _GEN_21150; // @[sequencer-master.scala 651:39]
  wire  _GEN_23609 = io_op_bits_active_vldx ? _GEN_22945 : _GEN_21151; // @[sequencer-master.scala 651:39]
  wire  _GEN_23610 = io_op_bits_active_vldx ? _GEN_22946 : _GEN_21152; // @[sequencer-master.scala 651:39]
  wire  _GEN_23611 = io_op_bits_active_vldx ? _GEN_22947 : _GEN_21153; // @[sequencer-master.scala 651:39]
  wire  _GEN_23612 = io_op_bits_active_vldx ? _GEN_22948 : _GEN_21154; // @[sequencer-master.scala 651:39]
  wire  _GEN_23613 = io_op_bits_active_vldx ? _GEN_22949 : _GEN_21155; // @[sequencer-master.scala 651:39]
  wire  _GEN_23614 = io_op_bits_active_vldx ? _GEN_23262 : _GEN_21156; // @[sequencer-master.scala 651:39]
  wire  _GEN_23615 = io_op_bits_active_vldx ? _GEN_23263 : _GEN_21157; // @[sequencer-master.scala 651:39]
  wire  _GEN_23616 = io_op_bits_active_vldx ? _GEN_23264 : _GEN_21158; // @[sequencer-master.scala 651:39]
  wire  _GEN_23617 = io_op_bits_active_vldx ? _GEN_23265 : _GEN_21159; // @[sequencer-master.scala 651:39]
  wire  _GEN_23618 = io_op_bits_active_vldx ? _GEN_23266 : _GEN_21160; // @[sequencer-master.scala 651:39]
  wire  _GEN_23619 = io_op_bits_active_vldx ? _GEN_23267 : _GEN_21161; // @[sequencer-master.scala 651:39]
  wire  _GEN_23620 = io_op_bits_active_vldx ? _GEN_23268 : _GEN_21162; // @[sequencer-master.scala 651:39]
  wire  _GEN_23621 = io_op_bits_active_vldx ? _GEN_23269 : _GEN_21163; // @[sequencer-master.scala 651:39]
  wire  _GEN_23622 = io_op_bits_active_vldx ? _GEN_23390 : _GEN_21164; // @[sequencer-master.scala 651:39]
  wire  _GEN_23623 = io_op_bits_active_vldx ? _GEN_23391 : _GEN_21165; // @[sequencer-master.scala 651:39]
  wire  _GEN_23624 = io_op_bits_active_vldx ? _GEN_23392 : _GEN_21166; // @[sequencer-master.scala 651:39]
  wire  _GEN_23625 = io_op_bits_active_vldx ? _GEN_23393 : _GEN_21167; // @[sequencer-master.scala 651:39]
  wire  _GEN_23626 = io_op_bits_active_vldx ? _GEN_23394 : _GEN_21168; // @[sequencer-master.scala 651:39]
  wire  _GEN_23627 = io_op_bits_active_vldx ? _GEN_23395 : _GEN_21169; // @[sequencer-master.scala 651:39]
  wire  _GEN_23628 = io_op_bits_active_vldx ? _GEN_23396 : _GEN_21170; // @[sequencer-master.scala 651:39]
  wire  _GEN_23629 = io_op_bits_active_vldx ? _GEN_23397 : _GEN_21171; // @[sequencer-master.scala 651:39]
  wire  _GEN_23630 = io_op_bits_active_vldx ? _GEN_22966 : _GEN_21172; // @[sequencer-master.scala 651:39]
  wire  _GEN_23631 = io_op_bits_active_vldx ? _GEN_22967 : _GEN_21173; // @[sequencer-master.scala 651:39]
  wire  _GEN_23632 = io_op_bits_active_vldx ? _GEN_22968 : _GEN_21174; // @[sequencer-master.scala 651:39]
  wire  _GEN_23633 = io_op_bits_active_vldx ? _GEN_22969 : _GEN_21175; // @[sequencer-master.scala 651:39]
  wire  _GEN_23634 = io_op_bits_active_vldx ? _GEN_22970 : _GEN_21176; // @[sequencer-master.scala 651:39]
  wire  _GEN_23635 = io_op_bits_active_vldx ? _GEN_22971 : _GEN_21177; // @[sequencer-master.scala 651:39]
  wire  _GEN_23636 = io_op_bits_active_vldx ? _GEN_22972 : _GEN_21178; // @[sequencer-master.scala 651:39]
  wire  _GEN_23637 = io_op_bits_active_vldx ? _GEN_22973 : _GEN_21179; // @[sequencer-master.scala 651:39]
  wire  _GEN_23638 = io_op_bits_active_vldx ? _GEN_23278 : _GEN_21180; // @[sequencer-master.scala 651:39]
  wire  _GEN_23639 = io_op_bits_active_vldx ? _GEN_23279 : _GEN_21181; // @[sequencer-master.scala 651:39]
  wire  _GEN_23640 = io_op_bits_active_vldx ? _GEN_23280 : _GEN_21182; // @[sequencer-master.scala 651:39]
  wire  _GEN_23641 = io_op_bits_active_vldx ? _GEN_23281 : _GEN_21183; // @[sequencer-master.scala 651:39]
  wire  _GEN_23642 = io_op_bits_active_vldx ? _GEN_23282 : _GEN_21184; // @[sequencer-master.scala 651:39]
  wire  _GEN_23643 = io_op_bits_active_vldx ? _GEN_23283 : _GEN_21185; // @[sequencer-master.scala 651:39]
  wire  _GEN_23644 = io_op_bits_active_vldx ? _GEN_23284 : _GEN_21186; // @[sequencer-master.scala 651:39]
  wire  _GEN_23645 = io_op_bits_active_vldx ? _GEN_23285 : _GEN_21187; // @[sequencer-master.scala 651:39]
  wire  _GEN_23646 = io_op_bits_active_vldx ? _GEN_23406 : _GEN_21188; // @[sequencer-master.scala 651:39]
  wire  _GEN_23647 = io_op_bits_active_vldx ? _GEN_23407 : _GEN_21189; // @[sequencer-master.scala 651:39]
  wire  _GEN_23648 = io_op_bits_active_vldx ? _GEN_23408 : _GEN_21190; // @[sequencer-master.scala 651:39]
  wire  _GEN_23649 = io_op_bits_active_vldx ? _GEN_23409 : _GEN_21191; // @[sequencer-master.scala 651:39]
  wire  _GEN_23650 = io_op_bits_active_vldx ? _GEN_23410 : _GEN_21192; // @[sequencer-master.scala 651:39]
  wire  _GEN_23651 = io_op_bits_active_vldx ? _GEN_23411 : _GEN_21193; // @[sequencer-master.scala 651:39]
  wire  _GEN_23652 = io_op_bits_active_vldx ? _GEN_23412 : _GEN_21194; // @[sequencer-master.scala 651:39]
  wire  _GEN_23653 = io_op_bits_active_vldx ? _GEN_23413 : _GEN_21195; // @[sequencer-master.scala 651:39]
  wire  _GEN_23654 = io_op_bits_active_vldx ? _GEN_22990 : _GEN_21196; // @[sequencer-master.scala 651:39]
  wire  _GEN_23655 = io_op_bits_active_vldx ? _GEN_22991 : _GEN_21197; // @[sequencer-master.scala 651:39]
  wire  _GEN_23656 = io_op_bits_active_vldx ? _GEN_22992 : _GEN_21198; // @[sequencer-master.scala 651:39]
  wire  _GEN_23657 = io_op_bits_active_vldx ? _GEN_22993 : _GEN_21199; // @[sequencer-master.scala 651:39]
  wire  _GEN_23658 = io_op_bits_active_vldx ? _GEN_22994 : _GEN_21200; // @[sequencer-master.scala 651:39]
  wire  _GEN_23659 = io_op_bits_active_vldx ? _GEN_22995 : _GEN_21201; // @[sequencer-master.scala 651:39]
  wire  _GEN_23660 = io_op_bits_active_vldx ? _GEN_22996 : _GEN_21202; // @[sequencer-master.scala 651:39]
  wire  _GEN_23661 = io_op_bits_active_vldx ? _GEN_22997 : _GEN_21203; // @[sequencer-master.scala 651:39]
  wire  _GEN_23662 = io_op_bits_active_vldx ? _GEN_23294 : _GEN_21204; // @[sequencer-master.scala 651:39]
  wire  _GEN_23663 = io_op_bits_active_vldx ? _GEN_23295 : _GEN_21205; // @[sequencer-master.scala 651:39]
  wire  _GEN_23664 = io_op_bits_active_vldx ? _GEN_23296 : _GEN_21206; // @[sequencer-master.scala 651:39]
  wire  _GEN_23665 = io_op_bits_active_vldx ? _GEN_23297 : _GEN_21207; // @[sequencer-master.scala 651:39]
  wire  _GEN_23666 = io_op_bits_active_vldx ? _GEN_23298 : _GEN_21208; // @[sequencer-master.scala 651:39]
  wire  _GEN_23667 = io_op_bits_active_vldx ? _GEN_23299 : _GEN_21209; // @[sequencer-master.scala 651:39]
  wire  _GEN_23668 = io_op_bits_active_vldx ? _GEN_23300 : _GEN_21210; // @[sequencer-master.scala 651:39]
  wire  _GEN_23669 = io_op_bits_active_vldx ? _GEN_23301 : _GEN_21211; // @[sequencer-master.scala 651:39]
  wire  _GEN_23670 = io_op_bits_active_vldx ? _GEN_23422 : _GEN_21212; // @[sequencer-master.scala 651:39]
  wire  _GEN_23671 = io_op_bits_active_vldx ? _GEN_23423 : _GEN_21213; // @[sequencer-master.scala 651:39]
  wire  _GEN_23672 = io_op_bits_active_vldx ? _GEN_23424 : _GEN_21214; // @[sequencer-master.scala 651:39]
  wire  _GEN_23673 = io_op_bits_active_vldx ? _GEN_23425 : _GEN_21215; // @[sequencer-master.scala 651:39]
  wire  _GEN_23674 = io_op_bits_active_vldx ? _GEN_23426 : _GEN_21216; // @[sequencer-master.scala 651:39]
  wire  _GEN_23675 = io_op_bits_active_vldx ? _GEN_23427 : _GEN_21217; // @[sequencer-master.scala 651:39]
  wire  _GEN_23676 = io_op_bits_active_vldx ? _GEN_23428 : _GEN_21218; // @[sequencer-master.scala 651:39]
  wire  _GEN_23677 = io_op_bits_active_vldx ? _GEN_23429 : _GEN_21219; // @[sequencer-master.scala 651:39]
  wire  _GEN_23678 = io_op_bits_active_vldx ? _GEN_23014 : _GEN_21220; // @[sequencer-master.scala 651:39]
  wire  _GEN_23679 = io_op_bits_active_vldx ? _GEN_23015 : _GEN_21221; // @[sequencer-master.scala 651:39]
  wire  _GEN_23680 = io_op_bits_active_vldx ? _GEN_23016 : _GEN_21222; // @[sequencer-master.scala 651:39]
  wire  _GEN_23681 = io_op_bits_active_vldx ? _GEN_23017 : _GEN_21223; // @[sequencer-master.scala 651:39]
  wire  _GEN_23682 = io_op_bits_active_vldx ? _GEN_23018 : _GEN_21224; // @[sequencer-master.scala 651:39]
  wire  _GEN_23683 = io_op_bits_active_vldx ? _GEN_23019 : _GEN_21225; // @[sequencer-master.scala 651:39]
  wire  _GEN_23684 = io_op_bits_active_vldx ? _GEN_23020 : _GEN_21226; // @[sequencer-master.scala 651:39]
  wire  _GEN_23685 = io_op_bits_active_vldx ? _GEN_23021 : _GEN_21227; // @[sequencer-master.scala 651:39]
  wire  _GEN_23686 = io_op_bits_active_vldx ? _GEN_23310 : _GEN_21228; // @[sequencer-master.scala 651:39]
  wire  _GEN_23687 = io_op_bits_active_vldx ? _GEN_23311 : _GEN_21229; // @[sequencer-master.scala 651:39]
  wire  _GEN_23688 = io_op_bits_active_vldx ? _GEN_23312 : _GEN_21230; // @[sequencer-master.scala 651:39]
  wire  _GEN_23689 = io_op_bits_active_vldx ? _GEN_23313 : _GEN_21231; // @[sequencer-master.scala 651:39]
  wire  _GEN_23690 = io_op_bits_active_vldx ? _GEN_23314 : _GEN_21232; // @[sequencer-master.scala 651:39]
  wire  _GEN_23691 = io_op_bits_active_vldx ? _GEN_23315 : _GEN_21233; // @[sequencer-master.scala 651:39]
  wire  _GEN_23692 = io_op_bits_active_vldx ? _GEN_23316 : _GEN_21234; // @[sequencer-master.scala 651:39]
  wire  _GEN_23693 = io_op_bits_active_vldx ? _GEN_23317 : _GEN_21235; // @[sequencer-master.scala 651:39]
  wire  _GEN_23694 = io_op_bits_active_vldx ? _GEN_23438 : _GEN_21236; // @[sequencer-master.scala 651:39]
  wire  _GEN_23695 = io_op_bits_active_vldx ? _GEN_23439 : _GEN_21237; // @[sequencer-master.scala 651:39]
  wire  _GEN_23696 = io_op_bits_active_vldx ? _GEN_23440 : _GEN_21238; // @[sequencer-master.scala 651:39]
  wire  _GEN_23697 = io_op_bits_active_vldx ? _GEN_23441 : _GEN_21239; // @[sequencer-master.scala 651:39]
  wire  _GEN_23698 = io_op_bits_active_vldx ? _GEN_23442 : _GEN_21240; // @[sequencer-master.scala 651:39]
  wire  _GEN_23699 = io_op_bits_active_vldx ? _GEN_23443 : _GEN_21241; // @[sequencer-master.scala 651:39]
  wire  _GEN_23700 = io_op_bits_active_vldx ? _GEN_23444 : _GEN_21242; // @[sequencer-master.scala 651:39]
  wire  _GEN_23701 = io_op_bits_active_vldx ? _GEN_23445 : _GEN_21243; // @[sequencer-master.scala 651:39]
  wire  _GEN_23702 = io_op_bits_active_vldx ? _GEN_23038 : _GEN_21244; // @[sequencer-master.scala 651:39]
  wire  _GEN_23703 = io_op_bits_active_vldx ? _GEN_23039 : _GEN_21245; // @[sequencer-master.scala 651:39]
  wire  _GEN_23704 = io_op_bits_active_vldx ? _GEN_23040 : _GEN_21246; // @[sequencer-master.scala 651:39]
  wire  _GEN_23705 = io_op_bits_active_vldx ? _GEN_23041 : _GEN_21247; // @[sequencer-master.scala 651:39]
  wire  _GEN_23706 = io_op_bits_active_vldx ? _GEN_23042 : _GEN_21248; // @[sequencer-master.scala 651:39]
  wire  _GEN_23707 = io_op_bits_active_vldx ? _GEN_23043 : _GEN_21249; // @[sequencer-master.scala 651:39]
  wire  _GEN_23708 = io_op_bits_active_vldx ? _GEN_23044 : _GEN_21250; // @[sequencer-master.scala 651:39]
  wire  _GEN_23709 = io_op_bits_active_vldx ? _GEN_23045 : _GEN_21251; // @[sequencer-master.scala 651:39]
  wire  _GEN_23710 = io_op_bits_active_vldx ? _GEN_23326 : _GEN_21252; // @[sequencer-master.scala 651:39]
  wire  _GEN_23711 = io_op_bits_active_vldx ? _GEN_23327 : _GEN_21253; // @[sequencer-master.scala 651:39]
  wire  _GEN_23712 = io_op_bits_active_vldx ? _GEN_23328 : _GEN_21254; // @[sequencer-master.scala 651:39]
  wire  _GEN_23713 = io_op_bits_active_vldx ? _GEN_23329 : _GEN_21255; // @[sequencer-master.scala 651:39]
  wire  _GEN_23714 = io_op_bits_active_vldx ? _GEN_23330 : _GEN_21256; // @[sequencer-master.scala 651:39]
  wire  _GEN_23715 = io_op_bits_active_vldx ? _GEN_23331 : _GEN_21257; // @[sequencer-master.scala 651:39]
  wire  _GEN_23716 = io_op_bits_active_vldx ? _GEN_23332 : _GEN_21258; // @[sequencer-master.scala 651:39]
  wire  _GEN_23717 = io_op_bits_active_vldx ? _GEN_23333 : _GEN_21259; // @[sequencer-master.scala 651:39]
  wire  _GEN_23718 = io_op_bits_active_vldx ? _GEN_23454 : _GEN_21260; // @[sequencer-master.scala 651:39]
  wire  _GEN_23719 = io_op_bits_active_vldx ? _GEN_23455 : _GEN_21261; // @[sequencer-master.scala 651:39]
  wire  _GEN_23720 = io_op_bits_active_vldx ? _GEN_23456 : _GEN_21262; // @[sequencer-master.scala 651:39]
  wire  _GEN_23721 = io_op_bits_active_vldx ? _GEN_23457 : _GEN_21263; // @[sequencer-master.scala 651:39]
  wire  _GEN_23722 = io_op_bits_active_vldx ? _GEN_23458 : _GEN_21264; // @[sequencer-master.scala 651:39]
  wire  _GEN_23723 = io_op_bits_active_vldx ? _GEN_23459 : _GEN_21265; // @[sequencer-master.scala 651:39]
  wire  _GEN_23724 = io_op_bits_active_vldx ? _GEN_23460 : _GEN_21266; // @[sequencer-master.scala 651:39]
  wire  _GEN_23725 = io_op_bits_active_vldx ? _GEN_23461 : _GEN_21267; // @[sequencer-master.scala 651:39]
  wire  _GEN_23726 = io_op_bits_active_vldx ? _GEN_23062 : _GEN_21268; // @[sequencer-master.scala 651:39]
  wire  _GEN_23727 = io_op_bits_active_vldx ? _GEN_23063 : _GEN_21269; // @[sequencer-master.scala 651:39]
  wire  _GEN_23728 = io_op_bits_active_vldx ? _GEN_23064 : _GEN_21270; // @[sequencer-master.scala 651:39]
  wire  _GEN_23729 = io_op_bits_active_vldx ? _GEN_23065 : _GEN_21271; // @[sequencer-master.scala 651:39]
  wire  _GEN_23730 = io_op_bits_active_vldx ? _GEN_23066 : _GEN_21272; // @[sequencer-master.scala 651:39]
  wire  _GEN_23731 = io_op_bits_active_vldx ? _GEN_23067 : _GEN_21273; // @[sequencer-master.scala 651:39]
  wire  _GEN_23732 = io_op_bits_active_vldx ? _GEN_23068 : _GEN_21274; // @[sequencer-master.scala 651:39]
  wire  _GEN_23733 = io_op_bits_active_vldx ? _GEN_23069 : _GEN_21275; // @[sequencer-master.scala 651:39]
  wire  _GEN_23734 = io_op_bits_active_vldx ? _GEN_23342 : _GEN_21276; // @[sequencer-master.scala 651:39]
  wire  _GEN_23735 = io_op_bits_active_vldx ? _GEN_23343 : _GEN_21277; // @[sequencer-master.scala 651:39]
  wire  _GEN_23736 = io_op_bits_active_vldx ? _GEN_23344 : _GEN_21278; // @[sequencer-master.scala 651:39]
  wire  _GEN_23737 = io_op_bits_active_vldx ? _GEN_23345 : _GEN_21279; // @[sequencer-master.scala 651:39]
  wire  _GEN_23738 = io_op_bits_active_vldx ? _GEN_23346 : _GEN_21280; // @[sequencer-master.scala 651:39]
  wire  _GEN_23739 = io_op_bits_active_vldx ? _GEN_23347 : _GEN_21281; // @[sequencer-master.scala 651:39]
  wire  _GEN_23740 = io_op_bits_active_vldx ? _GEN_23348 : _GEN_21282; // @[sequencer-master.scala 651:39]
  wire  _GEN_23741 = io_op_bits_active_vldx ? _GEN_23349 : _GEN_21283; // @[sequencer-master.scala 651:39]
  wire  _GEN_23742 = io_op_bits_active_vldx ? _GEN_23470 : _GEN_21284; // @[sequencer-master.scala 651:39]
  wire  _GEN_23743 = io_op_bits_active_vldx ? _GEN_23471 : _GEN_21285; // @[sequencer-master.scala 651:39]
  wire  _GEN_23744 = io_op_bits_active_vldx ? _GEN_23472 : _GEN_21286; // @[sequencer-master.scala 651:39]
  wire  _GEN_23745 = io_op_bits_active_vldx ? _GEN_23473 : _GEN_21287; // @[sequencer-master.scala 651:39]
  wire  _GEN_23746 = io_op_bits_active_vldx ? _GEN_23474 : _GEN_21288; // @[sequencer-master.scala 651:39]
  wire  _GEN_23747 = io_op_bits_active_vldx ? _GEN_23475 : _GEN_21289; // @[sequencer-master.scala 651:39]
  wire  _GEN_23748 = io_op_bits_active_vldx ? _GEN_23476 : _GEN_21290; // @[sequencer-master.scala 651:39]
  wire  _GEN_23749 = io_op_bits_active_vldx ? _GEN_23477 : _GEN_21291; // @[sequencer-master.scala 651:39]
  wire  _GEN_23750 = io_op_bits_active_vldx ? _GEN_23086 : _GEN_21292; // @[sequencer-master.scala 651:39]
  wire  _GEN_23751 = io_op_bits_active_vldx ? _GEN_23087 : _GEN_21293; // @[sequencer-master.scala 651:39]
  wire  _GEN_23752 = io_op_bits_active_vldx ? _GEN_23088 : _GEN_21294; // @[sequencer-master.scala 651:39]
  wire  _GEN_23753 = io_op_bits_active_vldx ? _GEN_23089 : _GEN_21295; // @[sequencer-master.scala 651:39]
  wire  _GEN_23754 = io_op_bits_active_vldx ? _GEN_23090 : _GEN_21296; // @[sequencer-master.scala 651:39]
  wire  _GEN_23755 = io_op_bits_active_vldx ? _GEN_23091 : _GEN_21297; // @[sequencer-master.scala 651:39]
  wire  _GEN_23756 = io_op_bits_active_vldx ? _GEN_23092 : _GEN_21298; // @[sequencer-master.scala 651:39]
  wire  _GEN_23757 = io_op_bits_active_vldx ? _GEN_23093 : _GEN_21299; // @[sequencer-master.scala 651:39]
  wire  _GEN_23758 = io_op_bits_active_vldx ? _GEN_23358 : _GEN_21300; // @[sequencer-master.scala 651:39]
  wire  _GEN_23759 = io_op_bits_active_vldx ? _GEN_23359 : _GEN_21301; // @[sequencer-master.scala 651:39]
  wire  _GEN_23760 = io_op_bits_active_vldx ? _GEN_23360 : _GEN_21302; // @[sequencer-master.scala 651:39]
  wire  _GEN_23761 = io_op_bits_active_vldx ? _GEN_23361 : _GEN_21303; // @[sequencer-master.scala 651:39]
  wire  _GEN_23762 = io_op_bits_active_vldx ? _GEN_23362 : _GEN_21304; // @[sequencer-master.scala 651:39]
  wire  _GEN_23763 = io_op_bits_active_vldx ? _GEN_23363 : _GEN_21305; // @[sequencer-master.scala 651:39]
  wire  _GEN_23764 = io_op_bits_active_vldx ? _GEN_23364 : _GEN_21306; // @[sequencer-master.scala 651:39]
  wire  _GEN_23765 = io_op_bits_active_vldx ? _GEN_23365 : _GEN_21307; // @[sequencer-master.scala 651:39]
  wire  _GEN_23766 = io_op_bits_active_vldx ? _GEN_23486 : _GEN_21308; // @[sequencer-master.scala 651:39]
  wire  _GEN_23767 = io_op_bits_active_vldx ? _GEN_23487 : _GEN_21309; // @[sequencer-master.scala 651:39]
  wire  _GEN_23768 = io_op_bits_active_vldx ? _GEN_23488 : _GEN_21310; // @[sequencer-master.scala 651:39]
  wire  _GEN_23769 = io_op_bits_active_vldx ? _GEN_23489 : _GEN_21311; // @[sequencer-master.scala 651:39]
  wire  _GEN_23770 = io_op_bits_active_vldx ? _GEN_23490 : _GEN_21312; // @[sequencer-master.scala 651:39]
  wire  _GEN_23771 = io_op_bits_active_vldx ? _GEN_23491 : _GEN_21313; // @[sequencer-master.scala 651:39]
  wire  _GEN_23772 = io_op_bits_active_vldx ? _GEN_23492 : _GEN_21314; // @[sequencer-master.scala 651:39]
  wire  _GEN_23773 = io_op_bits_active_vldx ? _GEN_23493 : _GEN_21315; // @[sequencer-master.scala 651:39]
  wire  _GEN_23774 = io_op_bits_active_vldx ? _GEN_23110 : _GEN_21316; // @[sequencer-master.scala 651:39]
  wire  _GEN_23775 = io_op_bits_active_vldx ? _GEN_23111 : _GEN_21317; // @[sequencer-master.scala 651:39]
  wire  _GEN_23776 = io_op_bits_active_vldx ? _GEN_23112 : _GEN_21318; // @[sequencer-master.scala 651:39]
  wire  _GEN_23777 = io_op_bits_active_vldx ? _GEN_23113 : _GEN_21319; // @[sequencer-master.scala 651:39]
  wire  _GEN_23778 = io_op_bits_active_vldx ? _GEN_23114 : _GEN_21320; // @[sequencer-master.scala 651:39]
  wire  _GEN_23779 = io_op_bits_active_vldx ? _GEN_23115 : _GEN_21321; // @[sequencer-master.scala 651:39]
  wire  _GEN_23780 = io_op_bits_active_vldx ? _GEN_23116 : _GEN_21322; // @[sequencer-master.scala 651:39]
  wire  _GEN_23781 = io_op_bits_active_vldx ? _GEN_23117 : _GEN_21323; // @[sequencer-master.scala 651:39]
  wire  _GEN_23790 = io_op_bits_active_vldx ? _GEN_21790 : _GEN_21332; // @[sequencer-master.scala 651:39]
  wire  _GEN_23791 = io_op_bits_active_vldx ? _GEN_21791 : _GEN_21333; // @[sequencer-master.scala 651:39]
  wire  _GEN_23792 = io_op_bits_active_vldx ? _GEN_21792 : _GEN_21334; // @[sequencer-master.scala 651:39]
  wire  _GEN_23793 = io_op_bits_active_vldx ? _GEN_21793 : _GEN_21335; // @[sequencer-master.scala 651:39]
  wire  _GEN_23794 = io_op_bits_active_vldx ? _GEN_21794 : _GEN_21336; // @[sequencer-master.scala 651:39]
  wire  _GEN_23795 = io_op_bits_active_vldx ? _GEN_21795 : _GEN_21337; // @[sequencer-master.scala 651:39]
  wire  _GEN_23796 = io_op_bits_active_vldx ? _GEN_21796 : _GEN_21338; // @[sequencer-master.scala 651:39]
  wire  _GEN_23797 = io_op_bits_active_vldx ? _GEN_21797 : _GEN_21339; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23798 = io_op_bits_active_vldx ? _GEN_23134 : _GEN_21340; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23799 = io_op_bits_active_vldx ? _GEN_23135 : _GEN_21341; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23800 = io_op_bits_active_vldx ? _GEN_23136 : _GEN_21342; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23801 = io_op_bits_active_vldx ? _GEN_23137 : _GEN_21343; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23802 = io_op_bits_active_vldx ? _GEN_23138 : _GEN_21344; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23803 = io_op_bits_active_vldx ? _GEN_23139 : _GEN_21345; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23804 = io_op_bits_active_vldx ? _GEN_23140 : _GEN_21346; // @[sequencer-master.scala 651:39]
  wire [9:0] _GEN_23805 = io_op_bits_active_vldx ? _GEN_23141 : _GEN_21347; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23806 = io_op_bits_active_vldx ? _GEN_21846 : _GEN_21348; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23807 = io_op_bits_active_vldx ? _GEN_21847 : _GEN_21349; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23808 = io_op_bits_active_vldx ? _GEN_21848 : _GEN_21350; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23809 = io_op_bits_active_vldx ? _GEN_21849 : _GEN_21351; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23810 = io_op_bits_active_vldx ? _GEN_21850 : _GEN_21352; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23811 = io_op_bits_active_vldx ? _GEN_21851 : _GEN_21353; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23812 = io_op_bits_active_vldx ? _GEN_21852 : _GEN_21354; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23813 = io_op_bits_active_vldx ? _GEN_21853 : _GEN_21355; // @[sequencer-master.scala 651:39]
  wire  _GEN_23814 = io_op_bits_active_vldx ? _GEN_21862 : _GEN_21356; // @[sequencer-master.scala 651:39]
  wire  _GEN_23815 = io_op_bits_active_vldx ? _GEN_21863 : _GEN_21357; // @[sequencer-master.scala 651:39]
  wire  _GEN_23816 = io_op_bits_active_vldx ? _GEN_21864 : _GEN_21358; // @[sequencer-master.scala 651:39]
  wire  _GEN_23817 = io_op_bits_active_vldx ? _GEN_21865 : _GEN_21359; // @[sequencer-master.scala 651:39]
  wire  _GEN_23818 = io_op_bits_active_vldx ? _GEN_21866 : _GEN_21360; // @[sequencer-master.scala 651:39]
  wire  _GEN_23819 = io_op_bits_active_vldx ? _GEN_21867 : _GEN_21361; // @[sequencer-master.scala 651:39]
  wire  _GEN_23820 = io_op_bits_active_vldx ? _GEN_21868 : _GEN_21362; // @[sequencer-master.scala 651:39]
  wire  _GEN_23821 = io_op_bits_active_vldx ? _GEN_21869 : _GEN_21363; // @[sequencer-master.scala 651:39]
  wire  _GEN_23822 = io_op_bits_active_vldx ? _GEN_21870 : _GEN_21364; // @[sequencer-master.scala 651:39]
  wire  _GEN_23823 = io_op_bits_active_vldx ? _GEN_21871 : _GEN_21365; // @[sequencer-master.scala 651:39]
  wire  _GEN_23824 = io_op_bits_active_vldx ? _GEN_21872 : _GEN_21366; // @[sequencer-master.scala 651:39]
  wire  _GEN_23825 = io_op_bits_active_vldx ? _GEN_21873 : _GEN_21367; // @[sequencer-master.scala 651:39]
  wire  _GEN_23826 = io_op_bits_active_vldx ? _GEN_21874 : _GEN_21368; // @[sequencer-master.scala 651:39]
  wire  _GEN_23827 = io_op_bits_active_vldx ? _GEN_21875 : _GEN_21369; // @[sequencer-master.scala 651:39]
  wire  _GEN_23828 = io_op_bits_active_vldx ? _GEN_21876 : _GEN_21370; // @[sequencer-master.scala 651:39]
  wire  _GEN_23829 = io_op_bits_active_vldx ? _GEN_21877 : _GEN_21371; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23830 = io_op_bits_active_vldx ? _GEN_21878 : _GEN_21372; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23831 = io_op_bits_active_vldx ? _GEN_21879 : _GEN_21373; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23832 = io_op_bits_active_vldx ? _GEN_21880 : _GEN_21374; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23833 = io_op_bits_active_vldx ? _GEN_21881 : _GEN_21375; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23834 = io_op_bits_active_vldx ? _GEN_21882 : _GEN_21376; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23835 = io_op_bits_active_vldx ? _GEN_21883 : _GEN_21377; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23836 = io_op_bits_active_vldx ? _GEN_21884 : _GEN_21378; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23837 = io_op_bits_active_vldx ? _GEN_21885 : _GEN_21379; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23838 = io_op_bits_active_vldx ? _GEN_22078 : _GEN_21380; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23839 = io_op_bits_active_vldx ? _GEN_22079 : _GEN_21381; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23840 = io_op_bits_active_vldx ? _GEN_22080 : _GEN_21382; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23841 = io_op_bits_active_vldx ? _GEN_22081 : _GEN_21383; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23842 = io_op_bits_active_vldx ? _GEN_22082 : _GEN_21384; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23843 = io_op_bits_active_vldx ? _GEN_22083 : _GEN_21385; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23844 = io_op_bits_active_vldx ? _GEN_22084 : _GEN_21386; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23845 = io_op_bits_active_vldx ? _GEN_22085 : _GEN_21387; // @[sequencer-master.scala 651:39]
  wire  _GEN_23846 = io_op_bits_active_vldx ? _GEN_22094 : _GEN_21388; // @[sequencer-master.scala 651:39]
  wire  _GEN_23847 = io_op_bits_active_vldx ? _GEN_22095 : _GEN_21389; // @[sequencer-master.scala 651:39]
  wire  _GEN_23848 = io_op_bits_active_vldx ? _GEN_22096 : _GEN_21390; // @[sequencer-master.scala 651:39]
  wire  _GEN_23849 = io_op_bits_active_vldx ? _GEN_22097 : _GEN_21391; // @[sequencer-master.scala 651:39]
  wire  _GEN_23850 = io_op_bits_active_vldx ? _GEN_22098 : _GEN_21392; // @[sequencer-master.scala 651:39]
  wire  _GEN_23851 = io_op_bits_active_vldx ? _GEN_22099 : _GEN_21393; // @[sequencer-master.scala 651:39]
  wire  _GEN_23852 = io_op_bits_active_vldx ? _GEN_22100 : _GEN_21394; // @[sequencer-master.scala 651:39]
  wire  _GEN_23853 = io_op_bits_active_vldx ? _GEN_22101 : _GEN_21395; // @[sequencer-master.scala 651:39]
  wire  _GEN_23854 = io_op_bits_active_vldx ? _GEN_22102 : _GEN_21396; // @[sequencer-master.scala 651:39]
  wire  _GEN_23855 = io_op_bits_active_vldx ? _GEN_22103 : _GEN_21397; // @[sequencer-master.scala 651:39]
  wire  _GEN_23856 = io_op_bits_active_vldx ? _GEN_22104 : _GEN_21398; // @[sequencer-master.scala 651:39]
  wire  _GEN_23857 = io_op_bits_active_vldx ? _GEN_22105 : _GEN_21399; // @[sequencer-master.scala 651:39]
  wire  _GEN_23858 = io_op_bits_active_vldx ? _GEN_22106 : _GEN_21400; // @[sequencer-master.scala 651:39]
  wire  _GEN_23859 = io_op_bits_active_vldx ? _GEN_22107 : _GEN_21401; // @[sequencer-master.scala 651:39]
  wire  _GEN_23860 = io_op_bits_active_vldx ? _GEN_22108 : _GEN_21402; // @[sequencer-master.scala 651:39]
  wire  _GEN_23861 = io_op_bits_active_vldx ? _GEN_22109 : _GEN_21403; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23862 = io_op_bits_active_vldx ? _GEN_22110 : _GEN_21404; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23863 = io_op_bits_active_vldx ? _GEN_22111 : _GEN_21405; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23864 = io_op_bits_active_vldx ? _GEN_22112 : _GEN_21406; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23865 = io_op_bits_active_vldx ? _GEN_22113 : _GEN_21407; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23866 = io_op_bits_active_vldx ? _GEN_22114 : _GEN_21408; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23867 = io_op_bits_active_vldx ? _GEN_22115 : _GEN_21409; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23868 = io_op_bits_active_vldx ? _GEN_22116 : _GEN_21410; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23869 = io_op_bits_active_vldx ? _GEN_22117 : _GEN_21411; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23870 = io_op_bits_active_vldx ? _GEN_22118 : _GEN_21412; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23871 = io_op_bits_active_vldx ? _GEN_22119 : _GEN_21413; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23872 = io_op_bits_active_vldx ? _GEN_22120 : _GEN_21414; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23873 = io_op_bits_active_vldx ? _GEN_22121 : _GEN_21415; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23874 = io_op_bits_active_vldx ? _GEN_22122 : _GEN_21416; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23875 = io_op_bits_active_vldx ? _GEN_22123 : _GEN_21417; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23876 = io_op_bits_active_vldx ? _GEN_22124 : _GEN_21418; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23877 = io_op_bits_active_vldx ? _GEN_22125 : _GEN_21419; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23878 = io_op_bits_active_vldx ? _GEN_22126 : _GEN_21420; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23879 = io_op_bits_active_vldx ? _GEN_22127 : _GEN_21421; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23880 = io_op_bits_active_vldx ? _GEN_22128 : _GEN_21422; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23881 = io_op_bits_active_vldx ? _GEN_22129 : _GEN_21423; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23882 = io_op_bits_active_vldx ? _GEN_22130 : _GEN_21424; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23883 = io_op_bits_active_vldx ? _GEN_22131 : _GEN_21425; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23884 = io_op_bits_active_vldx ? _GEN_22132 : _GEN_21426; // @[sequencer-master.scala 651:39]
  wire [63:0] _GEN_23885 = io_op_bits_active_vldx ? _GEN_22133 : _GEN_21427; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23886 = io_op_bits_active_vldx ? _GEN_23494 : _GEN_21428; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23887 = io_op_bits_active_vldx ? _GEN_23495 : _GEN_21429; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23888 = io_op_bits_active_vldx ? _GEN_23496 : _GEN_21430; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23889 = io_op_bits_active_vldx ? _GEN_23497 : _GEN_21431; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23890 = io_op_bits_active_vldx ? _GEN_23498 : _GEN_21432; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23891 = io_op_bits_active_vldx ? _GEN_23499 : _GEN_21433; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23892 = io_op_bits_active_vldx ? _GEN_23500 : _GEN_21434; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23893 = io_op_bits_active_vldx ? _GEN_23501 : _GEN_21435; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23894 = io_op_bits_active_vldx ? _GEN_23502 : _GEN_21436; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23895 = io_op_bits_active_vldx ? _GEN_23503 : _GEN_21437; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23896 = io_op_bits_active_vldx ? _GEN_23504 : _GEN_21438; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23897 = io_op_bits_active_vldx ? _GEN_23505 : _GEN_21439; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23898 = io_op_bits_active_vldx ? _GEN_23506 : _GEN_21440; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23899 = io_op_bits_active_vldx ? _GEN_23507 : _GEN_21441; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23900 = io_op_bits_active_vldx ? _GEN_23508 : _GEN_21442; // @[sequencer-master.scala 651:39]
  wire [3:0] _GEN_23901 = io_op_bits_active_vldx ? _GEN_23509 : _GEN_21443; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23902 = io_op_bits_active_vldx ? _GEN_23510 : _GEN_21444; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23903 = io_op_bits_active_vldx ? _GEN_23511 : _GEN_21445; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23904 = io_op_bits_active_vldx ? _GEN_23512 : _GEN_21446; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23905 = io_op_bits_active_vldx ? _GEN_23513 : _GEN_21447; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23906 = io_op_bits_active_vldx ? _GEN_23514 : _GEN_21448; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23907 = io_op_bits_active_vldx ? _GEN_23515 : _GEN_21449; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23908 = io_op_bits_active_vldx ? _GEN_23516 : _GEN_21450; // @[sequencer-master.scala 651:39]
  wire [2:0] _GEN_23909 = io_op_bits_active_vldx ? _GEN_23517 : _GEN_21451; // @[sequencer-master.scala 651:39]
  wire  _GEN_23910 = io_op_bits_active_vldx ? _GEN_22558 : _GEN_21452; // @[sequencer-master.scala 651:39]
  wire  _GEN_23911 = io_op_bits_active_vldx ? _GEN_22559 : _GEN_21453; // @[sequencer-master.scala 651:39]
  wire  _GEN_23912 = io_op_bits_active_vldx ? _GEN_22560 : _GEN_21454; // @[sequencer-master.scala 651:39]
  wire  _GEN_23913 = io_op_bits_active_vldx ? _GEN_22561 : _GEN_21455; // @[sequencer-master.scala 651:39]
  wire  _GEN_23914 = io_op_bits_active_vldx ? _GEN_22562 : _GEN_21456; // @[sequencer-master.scala 651:39]
  wire  _GEN_23915 = io_op_bits_active_vldx ? _GEN_22563 : _GEN_21457; // @[sequencer-master.scala 651:39]
  wire  _GEN_23916 = io_op_bits_active_vldx ? _GEN_22564 : _GEN_21458; // @[sequencer-master.scala 651:39]
  wire  _GEN_23917 = io_op_bits_active_vldx ? _GEN_22565 : _GEN_21459; // @[sequencer-master.scala 651:39]
  wire  _GEN_23918 = io_op_bits_active_vldx ? _GEN_23126 : _GEN_21468; // @[sequencer-master.scala 651:39]
  wire  _GEN_23919 = io_op_bits_active_vldx ? _GEN_23127 : _GEN_21469; // @[sequencer-master.scala 651:39]
  wire  _GEN_23920 = io_op_bits_active_vldx ? _GEN_23128 : _GEN_21470; // @[sequencer-master.scala 651:39]
  wire  _GEN_23921 = io_op_bits_active_vldx ? _GEN_23129 : _GEN_21471; // @[sequencer-master.scala 651:39]
  wire  _GEN_23922 = io_op_bits_active_vldx ? _GEN_23130 : _GEN_21472; // @[sequencer-master.scala 651:39]
  wire  _GEN_23923 = io_op_bits_active_vldx ? _GEN_23131 : _GEN_21473; // @[sequencer-master.scala 651:39]
  wire  _GEN_23924 = io_op_bits_active_vldx ? _GEN_23132 : _GEN_21474; // @[sequencer-master.scala 651:39]
  wire  _GEN_23925 = io_op_bits_active_vldx ? _GEN_23133 : _GEN_21475; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23926 = io_op_bits_active_vldx ? _GEN_23190 : _GEN_21476; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23927 = io_op_bits_active_vldx ? _GEN_23191 : _GEN_21477; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23928 = io_op_bits_active_vldx ? _GEN_23192 : _GEN_21478; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23929 = io_op_bits_active_vldx ? _GEN_23193 : _GEN_21479; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23930 = io_op_bits_active_vldx ? _GEN_23194 : _GEN_21480; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23931 = io_op_bits_active_vldx ? _GEN_23195 : _GEN_21481; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23932 = io_op_bits_active_vldx ? _GEN_23196 : _GEN_21482; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23933 = io_op_bits_active_vldx ? _GEN_23197 : _GEN_21483; // @[sequencer-master.scala 651:39]
  wire  _GEN_23934 = io_op_bits_active_vldx ? _GEN_23206 : _GEN_21484; // @[sequencer-master.scala 651:39]
  wire  _GEN_23935 = io_op_bits_active_vldx ? _GEN_23207 : _GEN_21485; // @[sequencer-master.scala 651:39]
  wire  _GEN_23936 = io_op_bits_active_vldx ? _GEN_23208 : _GEN_21486; // @[sequencer-master.scala 651:39]
  wire  _GEN_23937 = io_op_bits_active_vldx ? _GEN_23209 : _GEN_21487; // @[sequencer-master.scala 651:39]
  wire  _GEN_23938 = io_op_bits_active_vldx ? _GEN_23210 : _GEN_21488; // @[sequencer-master.scala 651:39]
  wire  _GEN_23939 = io_op_bits_active_vldx ? _GEN_23211 : _GEN_21489; // @[sequencer-master.scala 651:39]
  wire  _GEN_23940 = io_op_bits_active_vldx ? _GEN_23212 : _GEN_21490; // @[sequencer-master.scala 651:39]
  wire  _GEN_23941 = io_op_bits_active_vldx ? _GEN_23213 : _GEN_21491; // @[sequencer-master.scala 651:39]
  wire  _GEN_23942 = io_op_bits_active_vldx ? _GEN_23214 : _GEN_21492; // @[sequencer-master.scala 651:39]
  wire  _GEN_23943 = io_op_bits_active_vldx ? _GEN_23215 : _GEN_21493; // @[sequencer-master.scala 651:39]
  wire  _GEN_23944 = io_op_bits_active_vldx ? _GEN_23216 : _GEN_21494; // @[sequencer-master.scala 651:39]
  wire  _GEN_23945 = io_op_bits_active_vldx ? _GEN_23217 : _GEN_21495; // @[sequencer-master.scala 651:39]
  wire  _GEN_23946 = io_op_bits_active_vldx ? _GEN_23218 : _GEN_21496; // @[sequencer-master.scala 651:39]
  wire  _GEN_23947 = io_op_bits_active_vldx ? _GEN_23219 : _GEN_21497; // @[sequencer-master.scala 651:39]
  wire  _GEN_23948 = io_op_bits_active_vldx ? _GEN_23220 : _GEN_21498; // @[sequencer-master.scala 651:39]
  wire  _GEN_23949 = io_op_bits_active_vldx ? _GEN_23221 : _GEN_21499; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23950 = io_op_bits_active_vldx ? _GEN_23222 : _GEN_21500; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23951 = io_op_bits_active_vldx ? _GEN_23223 : _GEN_21501; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23952 = io_op_bits_active_vldx ? _GEN_23224 : _GEN_21502; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23953 = io_op_bits_active_vldx ? _GEN_23225 : _GEN_21503; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23954 = io_op_bits_active_vldx ? _GEN_23226 : _GEN_21504; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23955 = io_op_bits_active_vldx ? _GEN_23227 : _GEN_21505; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23956 = io_op_bits_active_vldx ? _GEN_23228 : _GEN_21506; // @[sequencer-master.scala 651:39]
  wire [1:0] _GEN_23957 = io_op_bits_active_vldx ? _GEN_23229 : _GEN_21507; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23958 = io_op_bits_active_vldx ? _GEN_23230 : _GEN_21508; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23959 = io_op_bits_active_vldx ? _GEN_23231 : _GEN_21509; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23960 = io_op_bits_active_vldx ? _GEN_23232 : _GEN_21510; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23961 = io_op_bits_active_vldx ? _GEN_23233 : _GEN_21511; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23962 = io_op_bits_active_vldx ? _GEN_23234 : _GEN_21512; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23963 = io_op_bits_active_vldx ? _GEN_23235 : _GEN_21513; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23964 = io_op_bits_active_vldx ? _GEN_23236 : _GEN_21514; // @[sequencer-master.scala 651:39]
  wire [7:0] _GEN_23965 = io_op_bits_active_vldx ? _GEN_23237 : _GEN_21515; // @[sequencer-master.scala 651:39]
  wire  _GEN_23966 = io_op_bits_active_vldx | _GEN_21516; // @[sequencer-master.scala 651:39 sequencer-master.scala 265:41]
  wire [2:0] _GEN_23967 = io_op_bits_active_vldx ? _T_1649 : _GEN_21517; // @[sequencer-master.scala 651:39 sequencer-master.scala 265:66]
  wire  _GEN_23984 = 3'h0 == tail ? 1'h0 : _GEN_23534; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23985 = 3'h1 == tail ? 1'h0 : _GEN_23535; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23986 = 3'h2 == tail ? 1'h0 : _GEN_23536; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23987 = 3'h3 == tail ? 1'h0 : _GEN_23537; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23988 = 3'h4 == tail ? 1'h0 : _GEN_23538; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23989 = 3'h5 == tail ? 1'h0 : _GEN_23539; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23990 = 3'h6 == tail ? 1'h0 : _GEN_23540; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23991 = 3'h7 == tail ? 1'h0 : _GEN_23541; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_23992 = 3'h0 == tail ? 1'h0 : _GEN_23542; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23993 = 3'h1 == tail ? 1'h0 : _GEN_23543; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23994 = 3'h2 == tail ? 1'h0 : _GEN_23544; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23995 = 3'h3 == tail ? 1'h0 : _GEN_23545; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23996 = 3'h4 == tail ? 1'h0 : _GEN_23546; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23997 = 3'h5 == tail ? 1'h0 : _GEN_23547; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23998 = 3'h6 == tail ? 1'h0 : _GEN_23548; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_23999 = 3'h7 == tail ? 1'h0 : _GEN_23549; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24000 = 3'h0 == tail ? 1'h0 : _GEN_23550; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24001 = 3'h1 == tail ? 1'h0 : _GEN_23551; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24002 = 3'h2 == tail ? 1'h0 : _GEN_23552; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24003 = 3'h3 == tail ? 1'h0 : _GEN_23553; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24004 = 3'h4 == tail ? 1'h0 : _GEN_23554; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24005 = 3'h5 == tail ? 1'h0 : _GEN_23555; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24006 = 3'h6 == tail ? 1'h0 : _GEN_23556; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24007 = 3'h7 == tail ? 1'h0 : _GEN_23557; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24008 = 3'h0 == tail ? 1'h0 : _GEN_23558; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24009 = 3'h1 == tail ? 1'h0 : _GEN_23559; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24010 = 3'h2 == tail ? 1'h0 : _GEN_23560; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24011 = 3'h3 == tail ? 1'h0 : _GEN_23561; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24012 = 3'h4 == tail ? 1'h0 : _GEN_23562; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24013 = 3'h5 == tail ? 1'h0 : _GEN_23563; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24014 = 3'h6 == tail ? 1'h0 : _GEN_23564; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24015 = 3'h7 == tail ? 1'h0 : _GEN_23565; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24016 = 3'h0 == tail ? 1'h0 : _GEN_23566; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24017 = 3'h1 == tail ? 1'h0 : _GEN_23567; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24018 = 3'h2 == tail ? 1'h0 : _GEN_23568; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24019 = 3'h3 == tail ? 1'h0 : _GEN_23569; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24020 = 3'h4 == tail ? 1'h0 : _GEN_23570; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24021 = 3'h5 == tail ? 1'h0 : _GEN_23571; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24022 = 3'h6 == tail ? 1'h0 : _GEN_23572; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24023 = 3'h7 == tail ? 1'h0 : _GEN_23573; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24032 = 3'h0 == tail ? 1'h0 : _GEN_23582; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24033 = 3'h1 == tail ? 1'h0 : _GEN_23583; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24034 = 3'h2 == tail ? 1'h0 : _GEN_23584; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24035 = 3'h3 == tail ? 1'h0 : _GEN_23585; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24036 = 3'h4 == tail ? 1'h0 : _GEN_23586; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24037 = 3'h5 == tail ? 1'h0 : _GEN_23587; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24038 = 3'h6 == tail ? 1'h0 : _GEN_23588; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24039 = 3'h7 == tail ? 1'h0 : _GEN_23589; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24040 = 3'h0 == tail ? 1'h0 : _GEN_23590; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24041 = 3'h1 == tail ? 1'h0 : _GEN_23591; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24042 = 3'h2 == tail ? 1'h0 : _GEN_23592; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24043 = 3'h3 == tail ? 1'h0 : _GEN_23593; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24044 = 3'h4 == tail ? 1'h0 : _GEN_23594; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24045 = 3'h5 == tail ? 1'h0 : _GEN_23595; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24046 = 3'h6 == tail ? 1'h0 : _GEN_23596; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24047 = 3'h7 == tail ? 1'h0 : _GEN_23597; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24048 = 3'h0 == tail ? 1'h0 : _GEN_23598; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24049 = 3'h1 == tail ? 1'h0 : _GEN_23599; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24050 = 3'h2 == tail ? 1'h0 : _GEN_23600; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24051 = 3'h3 == tail ? 1'h0 : _GEN_23601; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24052 = 3'h4 == tail ? 1'h0 : _GEN_23602; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24053 = 3'h5 == tail ? 1'h0 : _GEN_23603; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24054 = 3'h6 == tail ? 1'h0 : _GEN_23604; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24055 = 3'h7 == tail ? 1'h0 : _GEN_23605; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24056 = 3'h0 == tail ? 1'h0 : _GEN_23606; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24057 = 3'h1 == tail ? 1'h0 : _GEN_23607; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24058 = 3'h2 == tail ? 1'h0 : _GEN_23608; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24059 = 3'h3 == tail ? 1'h0 : _GEN_23609; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24060 = 3'h4 == tail ? 1'h0 : _GEN_23610; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24061 = 3'h5 == tail ? 1'h0 : _GEN_23611; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24062 = 3'h6 == tail ? 1'h0 : _GEN_23612; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24063 = 3'h7 == tail ? 1'h0 : _GEN_23613; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24064 = 3'h0 == tail ? 1'h0 : _GEN_23614; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24065 = 3'h1 == tail ? 1'h0 : _GEN_23615; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24066 = 3'h2 == tail ? 1'h0 : _GEN_23616; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24067 = 3'h3 == tail ? 1'h0 : _GEN_23617; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24068 = 3'h4 == tail ? 1'h0 : _GEN_23618; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24069 = 3'h5 == tail ? 1'h0 : _GEN_23619; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24070 = 3'h6 == tail ? 1'h0 : _GEN_23620; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24071 = 3'h7 == tail ? 1'h0 : _GEN_23621; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24072 = 3'h0 == tail ? 1'h0 : _GEN_23622; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24073 = 3'h1 == tail ? 1'h0 : _GEN_23623; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24074 = 3'h2 == tail ? 1'h0 : _GEN_23624; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24075 = 3'h3 == tail ? 1'h0 : _GEN_23625; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24076 = 3'h4 == tail ? 1'h0 : _GEN_23626; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24077 = 3'h5 == tail ? 1'h0 : _GEN_23627; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24078 = 3'h6 == tail ? 1'h0 : _GEN_23628; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24079 = 3'h7 == tail ? 1'h0 : _GEN_23629; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24080 = 3'h0 == tail ? 1'h0 : _GEN_23630; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24081 = 3'h1 == tail ? 1'h0 : _GEN_23631; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24082 = 3'h2 == tail ? 1'h0 : _GEN_23632; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24083 = 3'h3 == tail ? 1'h0 : _GEN_23633; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24084 = 3'h4 == tail ? 1'h0 : _GEN_23634; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24085 = 3'h5 == tail ? 1'h0 : _GEN_23635; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24086 = 3'h6 == tail ? 1'h0 : _GEN_23636; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24087 = 3'h7 == tail ? 1'h0 : _GEN_23637; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24088 = 3'h0 == tail ? 1'h0 : _GEN_23638; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24089 = 3'h1 == tail ? 1'h0 : _GEN_23639; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24090 = 3'h2 == tail ? 1'h0 : _GEN_23640; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24091 = 3'h3 == tail ? 1'h0 : _GEN_23641; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24092 = 3'h4 == tail ? 1'h0 : _GEN_23642; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24093 = 3'h5 == tail ? 1'h0 : _GEN_23643; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24094 = 3'h6 == tail ? 1'h0 : _GEN_23644; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24095 = 3'h7 == tail ? 1'h0 : _GEN_23645; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24096 = 3'h0 == tail ? 1'h0 : _GEN_23646; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24097 = 3'h1 == tail ? 1'h0 : _GEN_23647; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24098 = 3'h2 == tail ? 1'h0 : _GEN_23648; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24099 = 3'h3 == tail ? 1'h0 : _GEN_23649; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24100 = 3'h4 == tail ? 1'h0 : _GEN_23650; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24101 = 3'h5 == tail ? 1'h0 : _GEN_23651; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24102 = 3'h6 == tail ? 1'h0 : _GEN_23652; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24103 = 3'h7 == tail ? 1'h0 : _GEN_23653; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24104 = 3'h0 == tail ? 1'h0 : _GEN_23654; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24105 = 3'h1 == tail ? 1'h0 : _GEN_23655; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24106 = 3'h2 == tail ? 1'h0 : _GEN_23656; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24107 = 3'h3 == tail ? 1'h0 : _GEN_23657; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24108 = 3'h4 == tail ? 1'h0 : _GEN_23658; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24109 = 3'h5 == tail ? 1'h0 : _GEN_23659; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24110 = 3'h6 == tail ? 1'h0 : _GEN_23660; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24111 = 3'h7 == tail ? 1'h0 : _GEN_23661; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24112 = 3'h0 == tail ? 1'h0 : _GEN_23662; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24113 = 3'h1 == tail ? 1'h0 : _GEN_23663; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24114 = 3'h2 == tail ? 1'h0 : _GEN_23664; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24115 = 3'h3 == tail ? 1'h0 : _GEN_23665; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24116 = 3'h4 == tail ? 1'h0 : _GEN_23666; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24117 = 3'h5 == tail ? 1'h0 : _GEN_23667; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24118 = 3'h6 == tail ? 1'h0 : _GEN_23668; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24119 = 3'h7 == tail ? 1'h0 : _GEN_23669; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24120 = 3'h0 == tail ? 1'h0 : _GEN_23670; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24121 = 3'h1 == tail ? 1'h0 : _GEN_23671; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24122 = 3'h2 == tail ? 1'h0 : _GEN_23672; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24123 = 3'h3 == tail ? 1'h0 : _GEN_23673; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24124 = 3'h4 == tail ? 1'h0 : _GEN_23674; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24125 = 3'h5 == tail ? 1'h0 : _GEN_23675; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24126 = 3'h6 == tail ? 1'h0 : _GEN_23676; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24127 = 3'h7 == tail ? 1'h0 : _GEN_23677; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24128 = 3'h0 == tail ? 1'h0 : _GEN_23678; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24129 = 3'h1 == tail ? 1'h0 : _GEN_23679; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24130 = 3'h2 == tail ? 1'h0 : _GEN_23680; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24131 = 3'h3 == tail ? 1'h0 : _GEN_23681; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24132 = 3'h4 == tail ? 1'h0 : _GEN_23682; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24133 = 3'h5 == tail ? 1'h0 : _GEN_23683; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24134 = 3'h6 == tail ? 1'h0 : _GEN_23684; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24135 = 3'h7 == tail ? 1'h0 : _GEN_23685; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24136 = 3'h0 == tail ? 1'h0 : _GEN_23686; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24137 = 3'h1 == tail ? 1'h0 : _GEN_23687; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24138 = 3'h2 == tail ? 1'h0 : _GEN_23688; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24139 = 3'h3 == tail ? 1'h0 : _GEN_23689; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24140 = 3'h4 == tail ? 1'h0 : _GEN_23690; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24141 = 3'h5 == tail ? 1'h0 : _GEN_23691; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24142 = 3'h6 == tail ? 1'h0 : _GEN_23692; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24143 = 3'h7 == tail ? 1'h0 : _GEN_23693; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24144 = 3'h0 == tail ? 1'h0 : _GEN_23694; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24145 = 3'h1 == tail ? 1'h0 : _GEN_23695; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24146 = 3'h2 == tail ? 1'h0 : _GEN_23696; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24147 = 3'h3 == tail ? 1'h0 : _GEN_23697; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24148 = 3'h4 == tail ? 1'h0 : _GEN_23698; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24149 = 3'h5 == tail ? 1'h0 : _GEN_23699; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24150 = 3'h6 == tail ? 1'h0 : _GEN_23700; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24151 = 3'h7 == tail ? 1'h0 : _GEN_23701; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24152 = 3'h0 == tail ? 1'h0 : _GEN_23702; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24153 = 3'h1 == tail ? 1'h0 : _GEN_23703; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24154 = 3'h2 == tail ? 1'h0 : _GEN_23704; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24155 = 3'h3 == tail ? 1'h0 : _GEN_23705; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24156 = 3'h4 == tail ? 1'h0 : _GEN_23706; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24157 = 3'h5 == tail ? 1'h0 : _GEN_23707; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24158 = 3'h6 == tail ? 1'h0 : _GEN_23708; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24159 = 3'h7 == tail ? 1'h0 : _GEN_23709; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24160 = 3'h0 == tail ? 1'h0 : _GEN_23710; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24161 = 3'h1 == tail ? 1'h0 : _GEN_23711; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24162 = 3'h2 == tail ? 1'h0 : _GEN_23712; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24163 = 3'h3 == tail ? 1'h0 : _GEN_23713; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24164 = 3'h4 == tail ? 1'h0 : _GEN_23714; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24165 = 3'h5 == tail ? 1'h0 : _GEN_23715; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24166 = 3'h6 == tail ? 1'h0 : _GEN_23716; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24167 = 3'h7 == tail ? 1'h0 : _GEN_23717; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24168 = 3'h0 == tail ? 1'h0 : _GEN_23718; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24169 = 3'h1 == tail ? 1'h0 : _GEN_23719; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24170 = 3'h2 == tail ? 1'h0 : _GEN_23720; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24171 = 3'h3 == tail ? 1'h0 : _GEN_23721; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24172 = 3'h4 == tail ? 1'h0 : _GEN_23722; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24173 = 3'h5 == tail ? 1'h0 : _GEN_23723; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24174 = 3'h6 == tail ? 1'h0 : _GEN_23724; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24175 = 3'h7 == tail ? 1'h0 : _GEN_23725; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24176 = 3'h0 == tail ? 1'h0 : _GEN_23726; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24177 = 3'h1 == tail ? 1'h0 : _GEN_23727; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24178 = 3'h2 == tail ? 1'h0 : _GEN_23728; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24179 = 3'h3 == tail ? 1'h0 : _GEN_23729; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24180 = 3'h4 == tail ? 1'h0 : _GEN_23730; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24181 = 3'h5 == tail ? 1'h0 : _GEN_23731; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24182 = 3'h6 == tail ? 1'h0 : _GEN_23732; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24183 = 3'h7 == tail ? 1'h0 : _GEN_23733; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24184 = 3'h0 == tail ? 1'h0 : _GEN_23734; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24185 = 3'h1 == tail ? 1'h0 : _GEN_23735; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24186 = 3'h2 == tail ? 1'h0 : _GEN_23736; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24187 = 3'h3 == tail ? 1'h0 : _GEN_23737; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24188 = 3'h4 == tail ? 1'h0 : _GEN_23738; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24189 = 3'h5 == tail ? 1'h0 : _GEN_23739; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24190 = 3'h6 == tail ? 1'h0 : _GEN_23740; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24191 = 3'h7 == tail ? 1'h0 : _GEN_23741; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24192 = 3'h0 == tail ? 1'h0 : _GEN_23742; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24193 = 3'h1 == tail ? 1'h0 : _GEN_23743; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24194 = 3'h2 == tail ? 1'h0 : _GEN_23744; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24195 = 3'h3 == tail ? 1'h0 : _GEN_23745; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24196 = 3'h4 == tail ? 1'h0 : _GEN_23746; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24197 = 3'h5 == tail ? 1'h0 : _GEN_23747; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24198 = 3'h6 == tail ? 1'h0 : _GEN_23748; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24199 = 3'h7 == tail ? 1'h0 : _GEN_23749; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24200 = 3'h0 == tail ? 1'h0 : _GEN_23750; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24201 = 3'h1 == tail ? 1'h0 : _GEN_23751; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24202 = 3'h2 == tail ? 1'h0 : _GEN_23752; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24203 = 3'h3 == tail ? 1'h0 : _GEN_23753; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24204 = 3'h4 == tail ? 1'h0 : _GEN_23754; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24205 = 3'h5 == tail ? 1'h0 : _GEN_23755; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24206 = 3'h6 == tail ? 1'h0 : _GEN_23756; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24207 = 3'h7 == tail ? 1'h0 : _GEN_23757; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24208 = 3'h0 == tail ? 1'h0 : _GEN_23758; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24209 = 3'h1 == tail ? 1'h0 : _GEN_23759; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24210 = 3'h2 == tail ? 1'h0 : _GEN_23760; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24211 = 3'h3 == tail ? 1'h0 : _GEN_23761; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24212 = 3'h4 == tail ? 1'h0 : _GEN_23762; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24213 = 3'h5 == tail ? 1'h0 : _GEN_23763; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24214 = 3'h6 == tail ? 1'h0 : _GEN_23764; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24215 = 3'h7 == tail ? 1'h0 : _GEN_23765; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24216 = 3'h0 == tail ? 1'h0 : _GEN_23766; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24217 = 3'h1 == tail ? 1'h0 : _GEN_23767; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24218 = 3'h2 == tail ? 1'h0 : _GEN_23768; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24219 = 3'h3 == tail ? 1'h0 : _GEN_23769; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24220 = 3'h4 == tail ? 1'h0 : _GEN_23770; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24221 = 3'h5 == tail ? 1'h0 : _GEN_23771; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24222 = 3'h6 == tail ? 1'h0 : _GEN_23772; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24223 = 3'h7 == tail ? 1'h0 : _GEN_23773; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24224 = 3'h0 == tail ? 1'h0 : _GEN_23774; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24225 = 3'h1 == tail ? 1'h0 : _GEN_23775; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24226 = 3'h2 == tail ? 1'h0 : _GEN_23776; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24227 = 3'h3 == tail ? 1'h0 : _GEN_23777; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24228 = 3'h4 == tail ? 1'h0 : _GEN_23778; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24229 = 3'h5 == tail ? 1'h0 : _GEN_23779; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24230 = 3'h6 == tail ? 1'h0 : _GEN_23780; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24231 = 3'h7 == tail ? 1'h0 : _GEN_23781; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24240 = _GEN_32729 | _GEN_23790; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24241 = _GEN_32730 | _GEN_23791; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24242 = _GEN_32731 | _GEN_23792; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24243 = _GEN_32732 | _GEN_23793; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24244 = _GEN_32733 | _GEN_23794; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24245 = _GEN_32734 | _GEN_23795; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24246 = _GEN_32735 | _GEN_23796; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_24247 = _GEN_32736 | _GEN_23797; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_24248 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_23798; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24249 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_23799; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24250 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_23800; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24251 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_23801; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24252 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_23802; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24253 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_23803; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24254 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_23804; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_24255 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_23805; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_24256 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_23806; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24257 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_23807; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24258 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_23808; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24259 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_23809; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24260 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_23810; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24261 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_23811; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24262 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_23812; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_24263 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_23813; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24264 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_23984; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24265 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_23985; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24266 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_23986; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24267 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_23987; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24268 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_23988; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24269 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_23989; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24270 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_23990; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24271 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_23991; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24272 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_23814; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24273 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_23815; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24274 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_23816; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24275 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_23817; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24276 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_23818; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24277 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_23819; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24278 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_23820; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24279 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_23821; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24280 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_23822; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24281 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_23823; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24282 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_23824; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24283 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_23825; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24284 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_23826; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24285 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_23827; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24286 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_23828; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_24287 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_23829; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_24288 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_23830; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24289 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_23831; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24290 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_23832; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24291 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_23833; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24292 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_23834; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24293 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_23835; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24294 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_23836; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_24295 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_23837; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_24296 = io_op_bits_base_vp_valid ? _GEN_24256 : _GEN_23806; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24297 = io_op_bits_base_vp_valid ? _GEN_24257 : _GEN_23807; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24298 = io_op_bits_base_vp_valid ? _GEN_24258 : _GEN_23808; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24299 = io_op_bits_base_vp_valid ? _GEN_24259 : _GEN_23809; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24300 = io_op_bits_base_vp_valid ? _GEN_24260 : _GEN_23810; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24301 = io_op_bits_base_vp_valid ? _GEN_24261 : _GEN_23811; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24302 = io_op_bits_base_vp_valid ? _GEN_24262 : _GEN_23812; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_24303 = io_op_bits_base_vp_valid ? _GEN_24263 : _GEN_23813; // @[sequencer-master.scala 320:41]
  wire  _GEN_24304 = io_op_bits_base_vp_valid ? _GEN_24264 : _GEN_23984; // @[sequencer-master.scala 320:41]
  wire  _GEN_24305 = io_op_bits_base_vp_valid ? _GEN_24265 : _GEN_23985; // @[sequencer-master.scala 320:41]
  wire  _GEN_24306 = io_op_bits_base_vp_valid ? _GEN_24266 : _GEN_23986; // @[sequencer-master.scala 320:41]
  wire  _GEN_24307 = io_op_bits_base_vp_valid ? _GEN_24267 : _GEN_23987; // @[sequencer-master.scala 320:41]
  wire  _GEN_24308 = io_op_bits_base_vp_valid ? _GEN_24268 : _GEN_23988; // @[sequencer-master.scala 320:41]
  wire  _GEN_24309 = io_op_bits_base_vp_valid ? _GEN_24269 : _GEN_23989; // @[sequencer-master.scala 320:41]
  wire  _GEN_24310 = io_op_bits_base_vp_valid ? _GEN_24270 : _GEN_23990; // @[sequencer-master.scala 320:41]
  wire  _GEN_24311 = io_op_bits_base_vp_valid ? _GEN_24271 : _GEN_23991; // @[sequencer-master.scala 320:41]
  wire  _GEN_24312 = io_op_bits_base_vp_valid ? _GEN_24272 : _GEN_23814; // @[sequencer-master.scala 320:41]
  wire  _GEN_24313 = io_op_bits_base_vp_valid ? _GEN_24273 : _GEN_23815; // @[sequencer-master.scala 320:41]
  wire  _GEN_24314 = io_op_bits_base_vp_valid ? _GEN_24274 : _GEN_23816; // @[sequencer-master.scala 320:41]
  wire  _GEN_24315 = io_op_bits_base_vp_valid ? _GEN_24275 : _GEN_23817; // @[sequencer-master.scala 320:41]
  wire  _GEN_24316 = io_op_bits_base_vp_valid ? _GEN_24276 : _GEN_23818; // @[sequencer-master.scala 320:41]
  wire  _GEN_24317 = io_op_bits_base_vp_valid ? _GEN_24277 : _GEN_23819; // @[sequencer-master.scala 320:41]
  wire  _GEN_24318 = io_op_bits_base_vp_valid ? _GEN_24278 : _GEN_23820; // @[sequencer-master.scala 320:41]
  wire  _GEN_24319 = io_op_bits_base_vp_valid ? _GEN_24279 : _GEN_23821; // @[sequencer-master.scala 320:41]
  wire  _GEN_24320 = io_op_bits_base_vp_valid ? _GEN_24280 : _GEN_23822; // @[sequencer-master.scala 320:41]
  wire  _GEN_24321 = io_op_bits_base_vp_valid ? _GEN_24281 : _GEN_23823; // @[sequencer-master.scala 320:41]
  wire  _GEN_24322 = io_op_bits_base_vp_valid ? _GEN_24282 : _GEN_23824; // @[sequencer-master.scala 320:41]
  wire  _GEN_24323 = io_op_bits_base_vp_valid ? _GEN_24283 : _GEN_23825; // @[sequencer-master.scala 320:41]
  wire  _GEN_24324 = io_op_bits_base_vp_valid ? _GEN_24284 : _GEN_23826; // @[sequencer-master.scala 320:41]
  wire  _GEN_24325 = io_op_bits_base_vp_valid ? _GEN_24285 : _GEN_23827; // @[sequencer-master.scala 320:41]
  wire  _GEN_24326 = io_op_bits_base_vp_valid ? _GEN_24286 : _GEN_23828; // @[sequencer-master.scala 320:41]
  wire  _GEN_24327 = io_op_bits_base_vp_valid ? _GEN_24287 : _GEN_23829; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24328 = io_op_bits_base_vp_valid ? _GEN_24288 : _GEN_23830; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24329 = io_op_bits_base_vp_valid ? _GEN_24289 : _GEN_23831; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24330 = io_op_bits_base_vp_valid ? _GEN_24290 : _GEN_23832; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24331 = io_op_bits_base_vp_valid ? _GEN_24291 : _GEN_23833; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24332 = io_op_bits_base_vp_valid ? _GEN_24292 : _GEN_23834; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24333 = io_op_bits_base_vp_valid ? _GEN_24293 : _GEN_23835; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24334 = io_op_bits_base_vp_valid ? _GEN_24294 : _GEN_23836; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_24335 = io_op_bits_base_vp_valid ? _GEN_24295 : _GEN_23837; // @[sequencer-master.scala 320:41]
  wire  _GEN_24336 = _GEN_32729 | _GEN_24032; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24337 = _GEN_32730 | _GEN_24033; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24338 = _GEN_32731 | _GEN_24034; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24339 = _GEN_32732 | _GEN_24035; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24340 = _GEN_32733 | _GEN_24036; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24341 = _GEN_32734 | _GEN_24037; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24342 = _GEN_32735 | _GEN_24038; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24343 = _GEN_32736 | _GEN_24039; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24344 = _T_26 ? _GEN_24336 : _GEN_24032; // @[sequencer-master.scala 154:24]
  wire  _GEN_24345 = _T_26 ? _GEN_24337 : _GEN_24033; // @[sequencer-master.scala 154:24]
  wire  _GEN_24346 = _T_26 ? _GEN_24338 : _GEN_24034; // @[sequencer-master.scala 154:24]
  wire  _GEN_24347 = _T_26 ? _GEN_24339 : _GEN_24035; // @[sequencer-master.scala 154:24]
  wire  _GEN_24348 = _T_26 ? _GEN_24340 : _GEN_24036; // @[sequencer-master.scala 154:24]
  wire  _GEN_24349 = _T_26 ? _GEN_24341 : _GEN_24037; // @[sequencer-master.scala 154:24]
  wire  _GEN_24350 = _T_26 ? _GEN_24342 : _GEN_24038; // @[sequencer-master.scala 154:24]
  wire  _GEN_24351 = _T_26 ? _GEN_24343 : _GEN_24039; // @[sequencer-master.scala 154:24]
  wire  _GEN_24352 = _GEN_32729 | _GEN_24056; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24353 = _GEN_32730 | _GEN_24057; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24354 = _GEN_32731 | _GEN_24058; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24355 = _GEN_32732 | _GEN_24059; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24356 = _GEN_32733 | _GEN_24060; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24357 = _GEN_32734 | _GEN_24061; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24358 = _GEN_32735 | _GEN_24062; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24359 = _GEN_32736 | _GEN_24063; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24360 = _T_48 ? _GEN_24352 : _GEN_24056; // @[sequencer-master.scala 154:24]
  wire  _GEN_24361 = _T_48 ? _GEN_24353 : _GEN_24057; // @[sequencer-master.scala 154:24]
  wire  _GEN_24362 = _T_48 ? _GEN_24354 : _GEN_24058; // @[sequencer-master.scala 154:24]
  wire  _GEN_24363 = _T_48 ? _GEN_24355 : _GEN_24059; // @[sequencer-master.scala 154:24]
  wire  _GEN_24364 = _T_48 ? _GEN_24356 : _GEN_24060; // @[sequencer-master.scala 154:24]
  wire  _GEN_24365 = _T_48 ? _GEN_24357 : _GEN_24061; // @[sequencer-master.scala 154:24]
  wire  _GEN_24366 = _T_48 ? _GEN_24358 : _GEN_24062; // @[sequencer-master.scala 154:24]
  wire  _GEN_24367 = _T_48 ? _GEN_24359 : _GEN_24063; // @[sequencer-master.scala 154:24]
  wire  _GEN_24368 = _GEN_32729 | _GEN_24080; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24369 = _GEN_32730 | _GEN_24081; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24370 = _GEN_32731 | _GEN_24082; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24371 = _GEN_32732 | _GEN_24083; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24372 = _GEN_32733 | _GEN_24084; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24373 = _GEN_32734 | _GEN_24085; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24374 = _GEN_32735 | _GEN_24086; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24375 = _GEN_32736 | _GEN_24087; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24376 = _T_70 ? _GEN_24368 : _GEN_24080; // @[sequencer-master.scala 154:24]
  wire  _GEN_24377 = _T_70 ? _GEN_24369 : _GEN_24081; // @[sequencer-master.scala 154:24]
  wire  _GEN_24378 = _T_70 ? _GEN_24370 : _GEN_24082; // @[sequencer-master.scala 154:24]
  wire  _GEN_24379 = _T_70 ? _GEN_24371 : _GEN_24083; // @[sequencer-master.scala 154:24]
  wire  _GEN_24380 = _T_70 ? _GEN_24372 : _GEN_24084; // @[sequencer-master.scala 154:24]
  wire  _GEN_24381 = _T_70 ? _GEN_24373 : _GEN_24085; // @[sequencer-master.scala 154:24]
  wire  _GEN_24382 = _T_70 ? _GEN_24374 : _GEN_24086; // @[sequencer-master.scala 154:24]
  wire  _GEN_24383 = _T_70 ? _GEN_24375 : _GEN_24087; // @[sequencer-master.scala 154:24]
  wire  _GEN_24384 = _GEN_32729 | _GEN_24104; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24385 = _GEN_32730 | _GEN_24105; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24386 = _GEN_32731 | _GEN_24106; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24387 = _GEN_32732 | _GEN_24107; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24388 = _GEN_32733 | _GEN_24108; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24389 = _GEN_32734 | _GEN_24109; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24390 = _GEN_32735 | _GEN_24110; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24391 = _GEN_32736 | _GEN_24111; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24392 = _T_92 ? _GEN_24384 : _GEN_24104; // @[sequencer-master.scala 154:24]
  wire  _GEN_24393 = _T_92 ? _GEN_24385 : _GEN_24105; // @[sequencer-master.scala 154:24]
  wire  _GEN_24394 = _T_92 ? _GEN_24386 : _GEN_24106; // @[sequencer-master.scala 154:24]
  wire  _GEN_24395 = _T_92 ? _GEN_24387 : _GEN_24107; // @[sequencer-master.scala 154:24]
  wire  _GEN_24396 = _T_92 ? _GEN_24388 : _GEN_24108; // @[sequencer-master.scala 154:24]
  wire  _GEN_24397 = _T_92 ? _GEN_24389 : _GEN_24109; // @[sequencer-master.scala 154:24]
  wire  _GEN_24398 = _T_92 ? _GEN_24390 : _GEN_24110; // @[sequencer-master.scala 154:24]
  wire  _GEN_24399 = _T_92 ? _GEN_24391 : _GEN_24111; // @[sequencer-master.scala 154:24]
  wire  _GEN_24400 = _GEN_32729 | _GEN_24128; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24401 = _GEN_32730 | _GEN_24129; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24402 = _GEN_32731 | _GEN_24130; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24403 = _GEN_32732 | _GEN_24131; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24404 = _GEN_32733 | _GEN_24132; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24405 = _GEN_32734 | _GEN_24133; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24406 = _GEN_32735 | _GEN_24134; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24407 = _GEN_32736 | _GEN_24135; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24408 = _T_114 ? _GEN_24400 : _GEN_24128; // @[sequencer-master.scala 154:24]
  wire  _GEN_24409 = _T_114 ? _GEN_24401 : _GEN_24129; // @[sequencer-master.scala 154:24]
  wire  _GEN_24410 = _T_114 ? _GEN_24402 : _GEN_24130; // @[sequencer-master.scala 154:24]
  wire  _GEN_24411 = _T_114 ? _GEN_24403 : _GEN_24131; // @[sequencer-master.scala 154:24]
  wire  _GEN_24412 = _T_114 ? _GEN_24404 : _GEN_24132; // @[sequencer-master.scala 154:24]
  wire  _GEN_24413 = _T_114 ? _GEN_24405 : _GEN_24133; // @[sequencer-master.scala 154:24]
  wire  _GEN_24414 = _T_114 ? _GEN_24406 : _GEN_24134; // @[sequencer-master.scala 154:24]
  wire  _GEN_24415 = _T_114 ? _GEN_24407 : _GEN_24135; // @[sequencer-master.scala 154:24]
  wire  _GEN_24416 = _GEN_32729 | _GEN_24152; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24417 = _GEN_32730 | _GEN_24153; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24418 = _GEN_32731 | _GEN_24154; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24419 = _GEN_32732 | _GEN_24155; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24420 = _GEN_32733 | _GEN_24156; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24421 = _GEN_32734 | _GEN_24157; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24422 = _GEN_32735 | _GEN_24158; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24423 = _GEN_32736 | _GEN_24159; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24424 = _T_136 ? _GEN_24416 : _GEN_24152; // @[sequencer-master.scala 154:24]
  wire  _GEN_24425 = _T_136 ? _GEN_24417 : _GEN_24153; // @[sequencer-master.scala 154:24]
  wire  _GEN_24426 = _T_136 ? _GEN_24418 : _GEN_24154; // @[sequencer-master.scala 154:24]
  wire  _GEN_24427 = _T_136 ? _GEN_24419 : _GEN_24155; // @[sequencer-master.scala 154:24]
  wire  _GEN_24428 = _T_136 ? _GEN_24420 : _GEN_24156; // @[sequencer-master.scala 154:24]
  wire  _GEN_24429 = _T_136 ? _GEN_24421 : _GEN_24157; // @[sequencer-master.scala 154:24]
  wire  _GEN_24430 = _T_136 ? _GEN_24422 : _GEN_24158; // @[sequencer-master.scala 154:24]
  wire  _GEN_24431 = _T_136 ? _GEN_24423 : _GEN_24159; // @[sequencer-master.scala 154:24]
  wire  _GEN_24432 = _GEN_32729 | _GEN_24176; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24433 = _GEN_32730 | _GEN_24177; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24434 = _GEN_32731 | _GEN_24178; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24435 = _GEN_32732 | _GEN_24179; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24436 = _GEN_32733 | _GEN_24180; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24437 = _GEN_32734 | _GEN_24181; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24438 = _GEN_32735 | _GEN_24182; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24439 = _GEN_32736 | _GEN_24183; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24440 = _T_158 ? _GEN_24432 : _GEN_24176; // @[sequencer-master.scala 154:24]
  wire  _GEN_24441 = _T_158 ? _GEN_24433 : _GEN_24177; // @[sequencer-master.scala 154:24]
  wire  _GEN_24442 = _T_158 ? _GEN_24434 : _GEN_24178; // @[sequencer-master.scala 154:24]
  wire  _GEN_24443 = _T_158 ? _GEN_24435 : _GEN_24179; // @[sequencer-master.scala 154:24]
  wire  _GEN_24444 = _T_158 ? _GEN_24436 : _GEN_24180; // @[sequencer-master.scala 154:24]
  wire  _GEN_24445 = _T_158 ? _GEN_24437 : _GEN_24181; // @[sequencer-master.scala 154:24]
  wire  _GEN_24446 = _T_158 ? _GEN_24438 : _GEN_24182; // @[sequencer-master.scala 154:24]
  wire  _GEN_24447 = _T_158 ? _GEN_24439 : _GEN_24183; // @[sequencer-master.scala 154:24]
  wire  _GEN_24448 = _GEN_32729 | _GEN_24200; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24449 = _GEN_32730 | _GEN_24201; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24450 = _GEN_32731 | _GEN_24202; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24451 = _GEN_32732 | _GEN_24203; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24452 = _GEN_32733 | _GEN_24204; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24453 = _GEN_32734 | _GEN_24205; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24454 = _GEN_32735 | _GEN_24206; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24455 = _GEN_32736 | _GEN_24207; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24456 = _T_180 ? _GEN_24448 : _GEN_24200; // @[sequencer-master.scala 154:24]
  wire  _GEN_24457 = _T_180 ? _GEN_24449 : _GEN_24201; // @[sequencer-master.scala 154:24]
  wire  _GEN_24458 = _T_180 ? _GEN_24450 : _GEN_24202; // @[sequencer-master.scala 154:24]
  wire  _GEN_24459 = _T_180 ? _GEN_24451 : _GEN_24203; // @[sequencer-master.scala 154:24]
  wire  _GEN_24460 = _T_180 ? _GEN_24452 : _GEN_24204; // @[sequencer-master.scala 154:24]
  wire  _GEN_24461 = _T_180 ? _GEN_24453 : _GEN_24205; // @[sequencer-master.scala 154:24]
  wire  _GEN_24462 = _T_180 ? _GEN_24454 : _GEN_24206; // @[sequencer-master.scala 154:24]
  wire  _GEN_24463 = _T_180 ? _GEN_24455 : _GEN_24207; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_24464 = 3'h0 == tail ? io_op_bits_base_vs2_id : _GEN_23838; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24465 = 3'h1 == tail ? io_op_bits_base_vs2_id : _GEN_23839; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24466 = 3'h2 == tail ? io_op_bits_base_vs2_id : _GEN_23840; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24467 = 3'h3 == tail ? io_op_bits_base_vs2_id : _GEN_23841; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24468 = 3'h4 == tail ? io_op_bits_base_vs2_id : _GEN_23842; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24469 = 3'h5 == tail ? io_op_bits_base_vs2_id : _GEN_23843; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24470 = 3'h6 == tail ? io_op_bits_base_vs2_id : _GEN_23844; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24471 = 3'h7 == tail ? io_op_bits_base_vs2_id : _GEN_23845; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24472 = 3'h0 == tail ? io_op_bits_base_vs2_valid : _GEN_23992; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24473 = 3'h1 == tail ? io_op_bits_base_vs2_valid : _GEN_23993; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24474 = 3'h2 == tail ? io_op_bits_base_vs2_valid : _GEN_23994; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24475 = 3'h3 == tail ? io_op_bits_base_vs2_valid : _GEN_23995; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24476 = 3'h4 == tail ? io_op_bits_base_vs2_valid : _GEN_23996; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24477 = 3'h5 == tail ? io_op_bits_base_vs2_valid : _GEN_23997; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24478 = 3'h6 == tail ? io_op_bits_base_vs2_valid : _GEN_23998; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24479 = 3'h7 == tail ? io_op_bits_base_vs2_valid : _GEN_23999; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24480 = 3'h0 == tail ? io_op_bits_base_vs2_scalar : _GEN_23846; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24481 = 3'h1 == tail ? io_op_bits_base_vs2_scalar : _GEN_23847; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24482 = 3'h2 == tail ? io_op_bits_base_vs2_scalar : _GEN_23848; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24483 = 3'h3 == tail ? io_op_bits_base_vs2_scalar : _GEN_23849; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24484 = 3'h4 == tail ? io_op_bits_base_vs2_scalar : _GEN_23850; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24485 = 3'h5 == tail ? io_op_bits_base_vs2_scalar : _GEN_23851; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24486 = 3'h6 == tail ? io_op_bits_base_vs2_scalar : _GEN_23852; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24487 = 3'h7 == tail ? io_op_bits_base_vs2_scalar : _GEN_23853; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24488 = 3'h0 == tail ? io_op_bits_base_vs2_pred : _GEN_23854; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24489 = 3'h1 == tail ? io_op_bits_base_vs2_pred : _GEN_23855; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24490 = 3'h2 == tail ? io_op_bits_base_vs2_pred : _GEN_23856; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24491 = 3'h3 == tail ? io_op_bits_base_vs2_pred : _GEN_23857; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24492 = 3'h4 == tail ? io_op_bits_base_vs2_pred : _GEN_23858; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24493 = 3'h5 == tail ? io_op_bits_base_vs2_pred : _GEN_23859; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24494 = 3'h6 == tail ? io_op_bits_base_vs2_pred : _GEN_23860; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire  _GEN_24495 = 3'h7 == tail ? io_op_bits_base_vs2_pred : _GEN_23861; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24496 = 3'h0 == tail ? io_op_bits_base_vs2_prec : _GEN_23862; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24497 = 3'h1 == tail ? io_op_bits_base_vs2_prec : _GEN_23863; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24498 = 3'h2 == tail ? io_op_bits_base_vs2_prec : _GEN_23864; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24499 = 3'h3 == tail ? io_op_bits_base_vs2_prec : _GEN_23865; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24500 = 3'h4 == tail ? io_op_bits_base_vs2_prec : _GEN_23866; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24501 = 3'h5 == tail ? io_op_bits_base_vs2_prec : _GEN_23867; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24502 = 3'h6 == tail ? io_op_bits_base_vs2_prec : _GEN_23868; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [1:0] _GEN_24503 = 3'h7 == tail ? io_op_bits_base_vs2_prec : _GEN_23869; // @[sequencer-master.scala 329:29 sequencer-master.scala 329:29]
  wire [7:0] _GEN_24504 = 3'h0 == tail ? io_op_bits_reg_vs2_id : _GEN_23870; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24505 = 3'h1 == tail ? io_op_bits_reg_vs2_id : _GEN_23871; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24506 = 3'h2 == tail ? io_op_bits_reg_vs2_id : _GEN_23872; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24507 = 3'h3 == tail ? io_op_bits_reg_vs2_id : _GEN_23873; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24508 = 3'h4 == tail ? io_op_bits_reg_vs2_id : _GEN_23874; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24509 = 3'h5 == tail ? io_op_bits_reg_vs2_id : _GEN_23875; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24510 = 3'h6 == tail ? io_op_bits_reg_vs2_id : _GEN_23876; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [7:0] _GEN_24511 = 3'h7 == tail ? io_op_bits_reg_vs2_id : _GEN_23877; // @[sequencer-master.scala 330:47 sequencer-master.scala 330:47]
  wire [63:0] _GEN_24512 = 3'h0 == tail ? io_op_bits_sreg_ss2 : _GEN_23878; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24513 = 3'h1 == tail ? io_op_bits_sreg_ss2 : _GEN_23879; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24514 = 3'h2 == tail ? io_op_bits_sreg_ss2 : _GEN_23880; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24515 = 3'h3 == tail ? io_op_bits_sreg_ss2 : _GEN_23881; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24516 = 3'h4 == tail ? io_op_bits_sreg_ss2 : _GEN_23882; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24517 = 3'h5 == tail ? io_op_bits_sreg_ss2 : _GEN_23883; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24518 = 3'h6 == tail ? io_op_bits_sreg_ss2 : _GEN_23884; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [63:0] _GEN_24519 = 3'h7 == tail ? io_op_bits_sreg_ss2 : _GEN_23885; // @[sequencer-master.scala 332:31 sequencer-master.scala 332:31]
  wire [7:0] _GEN_24528 = io_op_bits_base_vs2_valid ? _GEN_24464 : _GEN_23838; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24529 = io_op_bits_base_vs2_valid ? _GEN_24465 : _GEN_23839; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24530 = io_op_bits_base_vs2_valid ? _GEN_24466 : _GEN_23840; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24531 = io_op_bits_base_vs2_valid ? _GEN_24467 : _GEN_23841; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24532 = io_op_bits_base_vs2_valid ? _GEN_24468 : _GEN_23842; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24533 = io_op_bits_base_vs2_valid ? _GEN_24469 : _GEN_23843; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24534 = io_op_bits_base_vs2_valid ? _GEN_24470 : _GEN_23844; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24535 = io_op_bits_base_vs2_valid ? _GEN_24471 : _GEN_23845; // @[sequencer-master.scala 328:47]
  wire  _GEN_24536 = io_op_bits_base_vs2_valid ? _GEN_24472 : _GEN_23992; // @[sequencer-master.scala 328:47]
  wire  _GEN_24537 = io_op_bits_base_vs2_valid ? _GEN_24473 : _GEN_23993; // @[sequencer-master.scala 328:47]
  wire  _GEN_24538 = io_op_bits_base_vs2_valid ? _GEN_24474 : _GEN_23994; // @[sequencer-master.scala 328:47]
  wire  _GEN_24539 = io_op_bits_base_vs2_valid ? _GEN_24475 : _GEN_23995; // @[sequencer-master.scala 328:47]
  wire  _GEN_24540 = io_op_bits_base_vs2_valid ? _GEN_24476 : _GEN_23996; // @[sequencer-master.scala 328:47]
  wire  _GEN_24541 = io_op_bits_base_vs2_valid ? _GEN_24477 : _GEN_23997; // @[sequencer-master.scala 328:47]
  wire  _GEN_24542 = io_op_bits_base_vs2_valid ? _GEN_24478 : _GEN_23998; // @[sequencer-master.scala 328:47]
  wire  _GEN_24543 = io_op_bits_base_vs2_valid ? _GEN_24479 : _GEN_23999; // @[sequencer-master.scala 328:47]
  wire  _GEN_24544 = io_op_bits_base_vs2_valid ? _GEN_24480 : _GEN_23846; // @[sequencer-master.scala 328:47]
  wire  _GEN_24545 = io_op_bits_base_vs2_valid ? _GEN_24481 : _GEN_23847; // @[sequencer-master.scala 328:47]
  wire  _GEN_24546 = io_op_bits_base_vs2_valid ? _GEN_24482 : _GEN_23848; // @[sequencer-master.scala 328:47]
  wire  _GEN_24547 = io_op_bits_base_vs2_valid ? _GEN_24483 : _GEN_23849; // @[sequencer-master.scala 328:47]
  wire  _GEN_24548 = io_op_bits_base_vs2_valid ? _GEN_24484 : _GEN_23850; // @[sequencer-master.scala 328:47]
  wire  _GEN_24549 = io_op_bits_base_vs2_valid ? _GEN_24485 : _GEN_23851; // @[sequencer-master.scala 328:47]
  wire  _GEN_24550 = io_op_bits_base_vs2_valid ? _GEN_24486 : _GEN_23852; // @[sequencer-master.scala 328:47]
  wire  _GEN_24551 = io_op_bits_base_vs2_valid ? _GEN_24487 : _GEN_23853; // @[sequencer-master.scala 328:47]
  wire  _GEN_24552 = io_op_bits_base_vs2_valid ? _GEN_24488 : _GEN_23854; // @[sequencer-master.scala 328:47]
  wire  _GEN_24553 = io_op_bits_base_vs2_valid ? _GEN_24489 : _GEN_23855; // @[sequencer-master.scala 328:47]
  wire  _GEN_24554 = io_op_bits_base_vs2_valid ? _GEN_24490 : _GEN_23856; // @[sequencer-master.scala 328:47]
  wire  _GEN_24555 = io_op_bits_base_vs2_valid ? _GEN_24491 : _GEN_23857; // @[sequencer-master.scala 328:47]
  wire  _GEN_24556 = io_op_bits_base_vs2_valid ? _GEN_24492 : _GEN_23858; // @[sequencer-master.scala 328:47]
  wire  _GEN_24557 = io_op_bits_base_vs2_valid ? _GEN_24493 : _GEN_23859; // @[sequencer-master.scala 328:47]
  wire  _GEN_24558 = io_op_bits_base_vs2_valid ? _GEN_24494 : _GEN_23860; // @[sequencer-master.scala 328:47]
  wire  _GEN_24559 = io_op_bits_base_vs2_valid ? _GEN_24495 : _GEN_23861; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24560 = io_op_bits_base_vs2_valid ? _GEN_24496 : _GEN_23862; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24561 = io_op_bits_base_vs2_valid ? _GEN_24497 : _GEN_23863; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24562 = io_op_bits_base_vs2_valid ? _GEN_24498 : _GEN_23864; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24563 = io_op_bits_base_vs2_valid ? _GEN_24499 : _GEN_23865; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24564 = io_op_bits_base_vs2_valid ? _GEN_24500 : _GEN_23866; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24565 = io_op_bits_base_vs2_valid ? _GEN_24501 : _GEN_23867; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24566 = io_op_bits_base_vs2_valid ? _GEN_24502 : _GEN_23868; // @[sequencer-master.scala 328:47]
  wire [1:0] _GEN_24567 = io_op_bits_base_vs2_valid ? _GEN_24503 : _GEN_23869; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24568 = io_op_bits_base_vs2_valid ? _GEN_24504 : _GEN_23870; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24569 = io_op_bits_base_vs2_valid ? _GEN_24505 : _GEN_23871; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24570 = io_op_bits_base_vs2_valid ? _GEN_24506 : _GEN_23872; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24571 = io_op_bits_base_vs2_valid ? _GEN_24507 : _GEN_23873; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24572 = io_op_bits_base_vs2_valid ? _GEN_24508 : _GEN_23874; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24573 = io_op_bits_base_vs2_valid ? _GEN_24509 : _GEN_23875; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24574 = io_op_bits_base_vs2_valid ? _GEN_24510 : _GEN_23876; // @[sequencer-master.scala 328:47]
  wire [7:0] _GEN_24575 = io_op_bits_base_vs2_valid ? _GEN_24511 : _GEN_23877; // @[sequencer-master.scala 328:47]
  wire  _GEN_24584 = _GEN_32729 | _GEN_24344; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24585 = _GEN_32730 | _GEN_24345; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24586 = _GEN_32731 | _GEN_24346; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24587 = _GEN_32732 | _GEN_24347; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24588 = _GEN_32733 | _GEN_24348; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24589 = _GEN_32734 | _GEN_24349; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24590 = _GEN_32735 | _GEN_24350; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24591 = _GEN_32736 | _GEN_24351; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24592 = _T_380 ? _GEN_24584 : _GEN_24344; // @[sequencer-master.scala 154:24]
  wire  _GEN_24593 = _T_380 ? _GEN_24585 : _GEN_24345; // @[sequencer-master.scala 154:24]
  wire  _GEN_24594 = _T_380 ? _GEN_24586 : _GEN_24346; // @[sequencer-master.scala 154:24]
  wire  _GEN_24595 = _T_380 ? _GEN_24587 : _GEN_24347; // @[sequencer-master.scala 154:24]
  wire  _GEN_24596 = _T_380 ? _GEN_24588 : _GEN_24348; // @[sequencer-master.scala 154:24]
  wire  _GEN_24597 = _T_380 ? _GEN_24589 : _GEN_24349; // @[sequencer-master.scala 154:24]
  wire  _GEN_24598 = _T_380 ? _GEN_24590 : _GEN_24350; // @[sequencer-master.scala 154:24]
  wire  _GEN_24599 = _T_380 ? _GEN_24591 : _GEN_24351; // @[sequencer-master.scala 154:24]
  wire  _GEN_24600 = _GEN_32729 | _GEN_24360; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24601 = _GEN_32730 | _GEN_24361; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24602 = _GEN_32731 | _GEN_24362; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24603 = _GEN_32732 | _GEN_24363; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24604 = _GEN_32733 | _GEN_24364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24605 = _GEN_32734 | _GEN_24365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24606 = _GEN_32735 | _GEN_24366; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24607 = _GEN_32736 | _GEN_24367; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24608 = _T_402 ? _GEN_24600 : _GEN_24360; // @[sequencer-master.scala 154:24]
  wire  _GEN_24609 = _T_402 ? _GEN_24601 : _GEN_24361; // @[sequencer-master.scala 154:24]
  wire  _GEN_24610 = _T_402 ? _GEN_24602 : _GEN_24362; // @[sequencer-master.scala 154:24]
  wire  _GEN_24611 = _T_402 ? _GEN_24603 : _GEN_24363; // @[sequencer-master.scala 154:24]
  wire  _GEN_24612 = _T_402 ? _GEN_24604 : _GEN_24364; // @[sequencer-master.scala 154:24]
  wire  _GEN_24613 = _T_402 ? _GEN_24605 : _GEN_24365; // @[sequencer-master.scala 154:24]
  wire  _GEN_24614 = _T_402 ? _GEN_24606 : _GEN_24366; // @[sequencer-master.scala 154:24]
  wire  _GEN_24615 = _T_402 ? _GEN_24607 : _GEN_24367; // @[sequencer-master.scala 154:24]
  wire  _GEN_24616 = _GEN_32729 | _GEN_24376; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24617 = _GEN_32730 | _GEN_24377; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24618 = _GEN_32731 | _GEN_24378; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24619 = _GEN_32732 | _GEN_24379; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24620 = _GEN_32733 | _GEN_24380; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24621 = _GEN_32734 | _GEN_24381; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24622 = _GEN_32735 | _GEN_24382; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24623 = _GEN_32736 | _GEN_24383; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24624 = _T_424 ? _GEN_24616 : _GEN_24376; // @[sequencer-master.scala 154:24]
  wire  _GEN_24625 = _T_424 ? _GEN_24617 : _GEN_24377; // @[sequencer-master.scala 154:24]
  wire  _GEN_24626 = _T_424 ? _GEN_24618 : _GEN_24378; // @[sequencer-master.scala 154:24]
  wire  _GEN_24627 = _T_424 ? _GEN_24619 : _GEN_24379; // @[sequencer-master.scala 154:24]
  wire  _GEN_24628 = _T_424 ? _GEN_24620 : _GEN_24380; // @[sequencer-master.scala 154:24]
  wire  _GEN_24629 = _T_424 ? _GEN_24621 : _GEN_24381; // @[sequencer-master.scala 154:24]
  wire  _GEN_24630 = _T_424 ? _GEN_24622 : _GEN_24382; // @[sequencer-master.scala 154:24]
  wire  _GEN_24631 = _T_424 ? _GEN_24623 : _GEN_24383; // @[sequencer-master.scala 154:24]
  wire  _GEN_24632 = _GEN_32729 | _GEN_24392; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24633 = _GEN_32730 | _GEN_24393; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24634 = _GEN_32731 | _GEN_24394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24635 = _GEN_32732 | _GEN_24395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24636 = _GEN_32733 | _GEN_24396; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24637 = _GEN_32734 | _GEN_24397; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24638 = _GEN_32735 | _GEN_24398; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24639 = _GEN_32736 | _GEN_24399; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24640 = _T_446 ? _GEN_24632 : _GEN_24392; // @[sequencer-master.scala 154:24]
  wire  _GEN_24641 = _T_446 ? _GEN_24633 : _GEN_24393; // @[sequencer-master.scala 154:24]
  wire  _GEN_24642 = _T_446 ? _GEN_24634 : _GEN_24394; // @[sequencer-master.scala 154:24]
  wire  _GEN_24643 = _T_446 ? _GEN_24635 : _GEN_24395; // @[sequencer-master.scala 154:24]
  wire  _GEN_24644 = _T_446 ? _GEN_24636 : _GEN_24396; // @[sequencer-master.scala 154:24]
  wire  _GEN_24645 = _T_446 ? _GEN_24637 : _GEN_24397; // @[sequencer-master.scala 154:24]
  wire  _GEN_24646 = _T_446 ? _GEN_24638 : _GEN_24398; // @[sequencer-master.scala 154:24]
  wire  _GEN_24647 = _T_446 ? _GEN_24639 : _GEN_24399; // @[sequencer-master.scala 154:24]
  wire  _GEN_24648 = _GEN_32729 | _GEN_24408; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24649 = _GEN_32730 | _GEN_24409; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24650 = _GEN_32731 | _GEN_24410; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24651 = _GEN_32732 | _GEN_24411; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24652 = _GEN_32733 | _GEN_24412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24653 = _GEN_32734 | _GEN_24413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24654 = _GEN_32735 | _GEN_24414; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24655 = _GEN_32736 | _GEN_24415; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24656 = _T_468 ? _GEN_24648 : _GEN_24408; // @[sequencer-master.scala 154:24]
  wire  _GEN_24657 = _T_468 ? _GEN_24649 : _GEN_24409; // @[sequencer-master.scala 154:24]
  wire  _GEN_24658 = _T_468 ? _GEN_24650 : _GEN_24410; // @[sequencer-master.scala 154:24]
  wire  _GEN_24659 = _T_468 ? _GEN_24651 : _GEN_24411; // @[sequencer-master.scala 154:24]
  wire  _GEN_24660 = _T_468 ? _GEN_24652 : _GEN_24412; // @[sequencer-master.scala 154:24]
  wire  _GEN_24661 = _T_468 ? _GEN_24653 : _GEN_24413; // @[sequencer-master.scala 154:24]
  wire  _GEN_24662 = _T_468 ? _GEN_24654 : _GEN_24414; // @[sequencer-master.scala 154:24]
  wire  _GEN_24663 = _T_468 ? _GEN_24655 : _GEN_24415; // @[sequencer-master.scala 154:24]
  wire  _GEN_24664 = _GEN_32729 | _GEN_24424; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24665 = _GEN_32730 | _GEN_24425; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24666 = _GEN_32731 | _GEN_24426; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24667 = _GEN_32732 | _GEN_24427; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24668 = _GEN_32733 | _GEN_24428; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24669 = _GEN_32734 | _GEN_24429; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24670 = _GEN_32735 | _GEN_24430; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24671 = _GEN_32736 | _GEN_24431; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24672 = _T_490 ? _GEN_24664 : _GEN_24424; // @[sequencer-master.scala 154:24]
  wire  _GEN_24673 = _T_490 ? _GEN_24665 : _GEN_24425; // @[sequencer-master.scala 154:24]
  wire  _GEN_24674 = _T_490 ? _GEN_24666 : _GEN_24426; // @[sequencer-master.scala 154:24]
  wire  _GEN_24675 = _T_490 ? _GEN_24667 : _GEN_24427; // @[sequencer-master.scala 154:24]
  wire  _GEN_24676 = _T_490 ? _GEN_24668 : _GEN_24428; // @[sequencer-master.scala 154:24]
  wire  _GEN_24677 = _T_490 ? _GEN_24669 : _GEN_24429; // @[sequencer-master.scala 154:24]
  wire  _GEN_24678 = _T_490 ? _GEN_24670 : _GEN_24430; // @[sequencer-master.scala 154:24]
  wire  _GEN_24679 = _T_490 ? _GEN_24671 : _GEN_24431; // @[sequencer-master.scala 154:24]
  wire  _GEN_24680 = _GEN_32729 | _GEN_24440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24681 = _GEN_32730 | _GEN_24441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24682 = _GEN_32731 | _GEN_24442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24683 = _GEN_32732 | _GEN_24443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24684 = _GEN_32733 | _GEN_24444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24685 = _GEN_32734 | _GEN_24445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24686 = _GEN_32735 | _GEN_24446; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24687 = _GEN_32736 | _GEN_24447; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24688 = _T_512 ? _GEN_24680 : _GEN_24440; // @[sequencer-master.scala 154:24]
  wire  _GEN_24689 = _T_512 ? _GEN_24681 : _GEN_24441; // @[sequencer-master.scala 154:24]
  wire  _GEN_24690 = _T_512 ? _GEN_24682 : _GEN_24442; // @[sequencer-master.scala 154:24]
  wire  _GEN_24691 = _T_512 ? _GEN_24683 : _GEN_24443; // @[sequencer-master.scala 154:24]
  wire  _GEN_24692 = _T_512 ? _GEN_24684 : _GEN_24444; // @[sequencer-master.scala 154:24]
  wire  _GEN_24693 = _T_512 ? _GEN_24685 : _GEN_24445; // @[sequencer-master.scala 154:24]
  wire  _GEN_24694 = _T_512 ? _GEN_24686 : _GEN_24446; // @[sequencer-master.scala 154:24]
  wire  _GEN_24695 = _T_512 ? _GEN_24687 : _GEN_24447; // @[sequencer-master.scala 154:24]
  wire  _GEN_24696 = _GEN_32729 | _GEN_24456; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24697 = _GEN_32730 | _GEN_24457; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24698 = _GEN_32731 | _GEN_24458; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24699 = _GEN_32732 | _GEN_24459; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24700 = _GEN_32733 | _GEN_24460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24701 = _GEN_32734 | _GEN_24461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24702 = _GEN_32735 | _GEN_24462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24703 = _GEN_32736 | _GEN_24463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_24704 = _T_534 ? _GEN_24696 : _GEN_24456; // @[sequencer-master.scala 154:24]
  wire  _GEN_24705 = _T_534 ? _GEN_24697 : _GEN_24457; // @[sequencer-master.scala 154:24]
  wire  _GEN_24706 = _T_534 ? _GEN_24698 : _GEN_24458; // @[sequencer-master.scala 154:24]
  wire  _GEN_24707 = _T_534 ? _GEN_24699 : _GEN_24459; // @[sequencer-master.scala 154:24]
  wire  _GEN_24708 = _T_534 ? _GEN_24700 : _GEN_24460; // @[sequencer-master.scala 154:24]
  wire  _GEN_24709 = _T_534 ? _GEN_24701 : _GEN_24461; // @[sequencer-master.scala 154:24]
  wire  _GEN_24710 = _T_534 ? _GEN_24702 : _GEN_24462; // @[sequencer-master.scala 154:24]
  wire  _GEN_24711 = _T_534 ? _GEN_24703 : _GEN_24463; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_24712 = 3'h0 == tail ? _e_T_1647_rports : _GEN_23886; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24713 = 3'h1 == tail ? _e_T_1647_rports : _GEN_23887; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24714 = 3'h2 == tail ? _e_T_1647_rports : _GEN_23888; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24715 = 3'h3 == tail ? _e_T_1647_rports : _GEN_23889; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24716 = 3'h4 == tail ? _e_T_1647_rports : _GEN_23890; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24717 = 3'h5 == tail ? _e_T_1647_rports : _GEN_23891; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24718 = 3'h6 == tail ? _e_T_1647_rports : _GEN_23892; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_24719 = 3'h7 == tail ? _e_T_1647_rports : _GEN_23893; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_24720 = 3'h0 == tail ? 4'h0 : _GEN_23894; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24721 = 3'h1 == tail ? 4'h0 : _GEN_23895; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24722 = 3'h2 == tail ? 4'h0 : _GEN_23896; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24723 = 3'h3 == tail ? 4'h0 : _GEN_23897; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24724 = 3'h4 == tail ? 4'h0 : _GEN_23898; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24725 = 3'h5 == tail ? 4'h0 : _GEN_23899; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24726 = 3'h6 == tail ? 4'h0 : _GEN_23900; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_24727 = 3'h7 == tail ? 4'h0 : _GEN_23901; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_24728 = 3'h0 == tail ? 3'h0 : _GEN_23902; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24729 = 3'h1 == tail ? 3'h0 : _GEN_23903; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24730 = 3'h2 == tail ? 3'h0 : _GEN_23904; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24731 = 3'h3 == tail ? 3'h0 : _GEN_23905; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24732 = 3'h4 == tail ? 3'h0 : _GEN_23906; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24733 = 3'h5 == tail ? 3'h0 : _GEN_23907; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24734 = 3'h6 == tail ? 3'h0 : _GEN_23908; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_24735 = 3'h7 == tail ? 3'h0 : _GEN_23909; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_24752 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24304; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24753 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24305; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24754 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24306; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24755 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24307; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24756 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24308; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24757 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24309; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24758 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24310; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24759 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24311; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_24760 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24536; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24761 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24537; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24762 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24538; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24763 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24539; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24764 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24540; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24765 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24541; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24766 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24542; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24767 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24543; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_24768 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24000; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24769 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24001; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24770 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24002; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24771 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24003; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24772 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24004; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24773 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24005; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24774 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24006; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24775 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24007; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_24776 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24008; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24777 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24009; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24778 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24010; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24779 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24011; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24780 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24012; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24781 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24013; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24782 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24014; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24783 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24015; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_24784 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24016; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24785 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24017; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24786 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24018; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24787 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24019; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24788 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24020; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24789 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24021; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24790 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24022; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24791 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24023; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_24800 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24592; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24801 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24593; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24802 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24594; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24803 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24595; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24804 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24596; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24805 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24597; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24806 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24598; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24807 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24599; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24808 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24040; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24809 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24041; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24810 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24042; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24811 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24043; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24812 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24044; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24813 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24045; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24814 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24046; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24815 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24047; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24816 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24048; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24817 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24049; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24818 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24050; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24819 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24051; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24820 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24052; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24821 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24053; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24822 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24054; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24823 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24055; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24824 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24608; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24825 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24609; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24826 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24610; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24827 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24611; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24828 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24612; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24829 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24613; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24830 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24614; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24831 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24615; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24832 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24064; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24833 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24065; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24834 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24066; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24835 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24067; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24836 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24068; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24837 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24069; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24838 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24070; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24839 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24071; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24840 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24072; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24841 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24073; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24842 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24074; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24843 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24075; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24844 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24076; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24845 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24077; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24846 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24078; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24847 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24079; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24848 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24624; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24849 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24625; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24850 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24626; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24851 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24627; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24852 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24628; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24853 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24629; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24854 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24630; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24855 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24631; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24856 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24088; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24857 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24089; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24858 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24090; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24859 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24091; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24860 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24092; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24861 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24093; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24862 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24094; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24863 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24095; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24864 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24096; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24865 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24097; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24866 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24098; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24867 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24099; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24868 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24100; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24869 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24101; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24870 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24102; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24871 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24103; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24872 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24640; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24873 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24641; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24874 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24642; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24875 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24643; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24876 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24644; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24877 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24645; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24878 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24646; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24879 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24647; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24880 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24112; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24881 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24113; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24882 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24114; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24883 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24115; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24884 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24116; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24885 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24117; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24886 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24118; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24887 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24119; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24888 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24120; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24889 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24121; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24890 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24122; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24891 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24123; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24892 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24124; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24893 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24125; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24894 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24126; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24895 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24127; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24896 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24656; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24897 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24657; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24898 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24658; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24899 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24659; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24900 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24660; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24901 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24661; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24902 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24662; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24903 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24663; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24904 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24136; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24905 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24137; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24906 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24138; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24907 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24139; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24908 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24140; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24909 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24141; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24910 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24142; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24911 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24143; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24912 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24144; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24913 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24145; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24914 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24146; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24915 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24147; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24916 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24148; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24917 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24149; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24918 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24150; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24919 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24151; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24920 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24672; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24921 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24673; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24922 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24674; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24923 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24675; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24924 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24676; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24925 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24677; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24926 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24678; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24927 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24679; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24928 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24160; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24929 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24161; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24930 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24162; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24931 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24163; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24932 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24164; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24933 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24165; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24934 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24166; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24935 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24167; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24936 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24168; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24937 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24169; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24938 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24170; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24939 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24171; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24940 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24172; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24941 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24173; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24942 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24174; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24943 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24175; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24944 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24688; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24945 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24689; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24946 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24690; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24947 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24691; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24948 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24692; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24949 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24693; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24950 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24694; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24951 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24695; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24952 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24184; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24953 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24185; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24954 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24186; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24955 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24187; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24956 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24188; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24957 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24189; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24958 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24190; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24959 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24191; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24960 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24192; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24961 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24193; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24962 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24194; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24963 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24195; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24964 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24196; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24965 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24197; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24966 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24198; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24967 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24199; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24968 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24704; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24969 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24705; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24970 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24706; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24971 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24707; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24972 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24708; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24973 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24709; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24974 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24710; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24975 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24711; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_24976 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24208; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24977 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24209; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24978 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24210; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24979 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24211; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24980 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24212; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24981 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24213; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24982 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24214; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24983 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24215; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_24984 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24216; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24985 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24217; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24986 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24218; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24987 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24219; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24988 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24220; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24989 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24221; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24990 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24222; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24991 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24223; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_24992 = 3'h0 == _T_1645 ? 1'h0 : _GEN_24224; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24993 = 3'h1 == _T_1645 ? 1'h0 : _GEN_24225; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24994 = 3'h2 == _T_1645 ? 1'h0 : _GEN_24226; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24995 = 3'h3 == _T_1645 ? 1'h0 : _GEN_24227; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24996 = 3'h4 == _T_1645 ? 1'h0 : _GEN_24228; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24997 = 3'h5 == _T_1645 ? 1'h0 : _GEN_24229; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24998 = 3'h6 == _T_1645 ? 1'h0 : _GEN_24230; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_24999 = 3'h7 == _T_1645 ? 1'h0 : _GEN_24231; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25008 = _GEN_34121 | _GEN_23910; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25009 = _GEN_34122 | _GEN_23911; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25010 = _GEN_34123 | _GEN_23912; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25011 = _GEN_34124 | _GEN_23913; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25012 = _GEN_34125 | _GEN_23914; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25013 = _GEN_34126 | _GEN_23915; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25014 = _GEN_34127 | _GEN_23916; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25015 = _GEN_34128 | _GEN_23917; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_25016 = 3'h0 == _T_1645 ? io_op_bits_fn_union : _GEN_24248; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25017 = 3'h1 == _T_1645 ? io_op_bits_fn_union : _GEN_24249; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25018 = 3'h2 == _T_1645 ? io_op_bits_fn_union : _GEN_24250; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25019 = 3'h3 == _T_1645 ? io_op_bits_fn_union : _GEN_24251; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25020 = 3'h4 == _T_1645 ? io_op_bits_fn_union : _GEN_24252; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25021 = 3'h5 == _T_1645 ? io_op_bits_fn_union : _GEN_24253; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25022 = 3'h6 == _T_1645 ? io_op_bits_fn_union : _GEN_24254; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25023 = 3'h7 == _T_1645 ? io_op_bits_fn_union : _GEN_24255; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [1:0] _GEN_25024 = 3'h0 == _T_1645 ? 2'h0 : _GEN_24712; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25025 = 3'h1 == _T_1645 ? 2'h0 : _GEN_24713; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25026 = 3'h2 == _T_1645 ? 2'h0 : _GEN_24714; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25027 = 3'h3 == _T_1645 ? 2'h0 : _GEN_24715; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25028 = 3'h4 == _T_1645 ? 2'h0 : _GEN_24716; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25029 = 3'h5 == _T_1645 ? 2'h0 : _GEN_24717; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25030 = 3'h6 == _T_1645 ? 2'h0 : _GEN_24718; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25031 = 3'h7 == _T_1645 ? 2'h0 : _GEN_24719; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_25032 = 3'h0 == _T_1645 ? 4'h0 : _GEN_24720; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25033 = 3'h1 == _T_1645 ? 4'h0 : _GEN_24721; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25034 = 3'h2 == _T_1645 ? 4'h0 : _GEN_24722; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25035 = 3'h3 == _T_1645 ? 4'h0 : _GEN_24723; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25036 = 3'h4 == _T_1645 ? 4'h0 : _GEN_24724; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25037 = 3'h5 == _T_1645 ? 4'h0 : _GEN_24725; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25038 = 3'h6 == _T_1645 ? 4'h0 : _GEN_24726; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25039 = 3'h7 == _T_1645 ? 4'h0 : _GEN_24727; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_25040 = 3'h0 == _T_1645 ? 3'h0 : _GEN_24728; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25041 = 3'h1 == _T_1645 ? 3'h0 : _GEN_24729; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25042 = 3'h2 == _T_1645 ? 3'h0 : _GEN_24730; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25043 = 3'h3 == _T_1645 ? 3'h0 : _GEN_24731; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25044 = 3'h4 == _T_1645 ? 3'h0 : _GEN_24732; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25045 = 3'h5 == _T_1645 ? 3'h0 : _GEN_24733; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25046 = 3'h6 == _T_1645 ? 3'h0 : _GEN_24734; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25047 = 3'h7 == _T_1645 ? 3'h0 : _GEN_24735; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_25048 = 3'h0 == _T_1647 | (3'h0 == _T_1645 | (_GEN_32729 | _GEN_23518)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25049 = 3'h1 == _T_1647 | (3'h1 == _T_1645 | (_GEN_32730 | _GEN_23519)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25050 = 3'h2 == _T_1647 | (3'h2 == _T_1645 | (_GEN_32731 | _GEN_23520)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25051 = 3'h3 == _T_1647 | (3'h3 == _T_1645 | (_GEN_32732 | _GEN_23521)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25052 = 3'h4 == _T_1647 | (3'h4 == _T_1645 | (_GEN_32733 | _GEN_23522)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25053 = 3'h5 == _T_1647 | (3'h5 == _T_1645 | (_GEN_32734 | _GEN_23523)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25054 = 3'h6 == _T_1647 | (3'h6 == _T_1645 | (_GEN_32735 | _GEN_23524)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25055 = 3'h7 == _T_1647 | (3'h7 == _T_1645 | (_GEN_32736 | _GEN_23525)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_25064 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24752; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25065 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24753; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25066 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24754; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25067 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24755; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25068 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24756; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25069 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24757; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25070 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24758; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25071 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24759; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_25072 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24760; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25073 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24761; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25074 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24762; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25075 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24763; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25076 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24764; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25077 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24765; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25078 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24766; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25079 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24767; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_25080 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24768; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25081 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24769; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25082 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24770; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25083 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24771; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25084 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24772; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25085 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24773; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25086 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24774; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25087 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24775; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_25088 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24776; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25089 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24777; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25090 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24778; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25091 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24779; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25092 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24780; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25093 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24781; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25094 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24782; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25095 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24783; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_25096 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24784; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25097 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24785; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25098 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24786; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25099 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24787; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25100 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24788; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25101 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24789; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25102 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24790; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25103 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24791; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_25104 = _GEN_36426 | (_GEN_34121 | (_GEN_32729 | _GEN_23574)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25105 = _GEN_36427 | (_GEN_34122 | (_GEN_32730 | _GEN_23575)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25106 = _GEN_36428 | (_GEN_34123 | (_GEN_32731 | _GEN_23576)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25107 = _GEN_36429 | (_GEN_34124 | (_GEN_32732 | _GEN_23577)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25108 = _GEN_36430 | (_GEN_34125 | (_GEN_32733 | _GEN_23578)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25109 = _GEN_36431 | (_GEN_34126 | (_GEN_32734 | _GEN_23579)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25110 = _GEN_36432 | (_GEN_34127 | (_GEN_32735 | _GEN_23580)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25111 = _GEN_36433 | (_GEN_34128 | (_GEN_32736 | _GEN_23581)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_25112 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24800; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25113 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24801; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25114 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24802; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25115 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24803; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25116 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24804; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25117 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24805; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25118 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24806; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25119 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24807; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25120 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24808; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25121 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24809; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25122 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24810; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25123 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24811; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25124 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24812; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25125 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24813; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25126 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24814; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25127 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24815; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25128 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24816; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25129 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24817; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25130 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24818; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25131 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24819; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25132 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24820; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25133 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24821; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25134 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24822; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25135 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24823; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25136 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24824; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25137 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24825; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25138 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24826; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25139 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24827; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25140 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24828; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25141 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24829; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25142 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24830; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25143 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24831; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25144 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24832; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25145 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24833; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25146 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24834; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25147 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24835; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25148 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24836; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25149 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24837; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25150 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24838; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25151 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24839; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25152 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24840; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25153 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24841; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25154 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24842; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25155 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24843; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25156 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24844; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25157 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24845; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25158 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24846; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25159 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24847; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25160 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24848; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25161 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24849; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25162 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24850; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25163 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24851; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25164 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24852; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25165 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24853; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25166 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24854; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25167 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24855; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25168 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24856; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25169 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24857; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25170 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24858; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25171 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24859; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25172 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24860; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25173 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24861; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25174 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24862; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25175 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24863; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25176 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24864; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25177 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24865; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25178 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24866; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25179 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24867; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25180 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24868; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25181 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24869; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25182 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24870; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25183 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24871; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25184 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24872; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25185 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24873; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25186 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24874; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25187 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24875; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25188 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24876; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25189 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24877; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25190 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24878; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25191 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24879; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25192 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24880; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25193 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24881; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25194 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24882; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25195 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24883; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25196 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24884; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25197 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24885; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25198 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24886; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25199 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24887; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25200 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24888; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25201 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24889; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25202 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24890; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25203 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24891; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25204 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24892; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25205 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24893; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25206 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24894; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25207 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24895; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25208 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24896; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25209 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24897; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25210 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24898; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25211 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24899; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25212 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24900; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25213 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24901; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25214 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24902; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25215 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24903; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25216 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24904; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25217 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24905; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25218 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24906; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25219 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24907; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25220 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24908; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25221 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24909; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25222 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24910; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25223 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24911; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25224 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24912; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25225 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24913; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25226 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24914; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25227 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24915; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25228 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24916; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25229 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24917; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25230 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24918; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25231 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24919; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25232 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24920; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25233 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24921; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25234 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24922; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25235 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24923; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25236 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24924; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25237 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24925; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25238 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24926; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25239 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24927; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25240 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24928; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25241 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24929; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25242 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24930; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25243 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24931; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25244 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24932; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25245 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24933; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25246 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24934; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25247 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24935; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25248 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24936; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25249 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24937; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25250 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24938; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25251 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24939; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25252 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24940; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25253 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24941; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25254 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24942; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25255 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24943; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25256 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24944; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25257 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24945; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25258 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24946; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25259 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24947; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25260 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24948; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25261 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24949; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25262 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24950; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25263 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24951; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25264 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24952; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25265 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24953; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25266 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24954; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25267 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24955; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25268 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24956; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25269 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24957; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25270 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24958; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25271 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24959; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25272 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24960; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25273 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24961; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25274 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24962; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25275 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24963; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25276 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24964; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25277 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24965; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25278 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24966; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25279 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24967; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25280 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24968; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25281 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24969; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25282 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24970; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25283 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24971; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25284 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24972; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25285 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24973; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25286 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24974; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25287 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24975; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_25288 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24976; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25289 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24977; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25290 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24978; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25291 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24979; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25292 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24980; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25293 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24981; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25294 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24982; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25295 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24983; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_25296 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24984; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25297 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24985; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25298 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24986; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25299 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24987; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25300 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24988; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25301 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24989; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25302 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24990; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25303 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24991; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_25304 = 3'h0 == _T_1647 ? 1'h0 : _GEN_24992; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25305 = 3'h1 == _T_1647 ? 1'h0 : _GEN_24993; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25306 = 3'h2 == _T_1647 ? 1'h0 : _GEN_24994; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25307 = 3'h3 == _T_1647 ? 1'h0 : _GEN_24995; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25308 = 3'h4 == _T_1647 ? 1'h0 : _GEN_24996; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25309 = 3'h5 == _T_1647 ? 1'h0 : _GEN_24997; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25310 = 3'h6 == _T_1647 ? 1'h0 : _GEN_24998; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25311 = 3'h7 == _T_1647 ? 1'h0 : _GEN_24999; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_25320 = _GEN_36426 | _GEN_21460; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25321 = _GEN_36427 | _GEN_21461; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25322 = _GEN_36428 | _GEN_21462; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25323 = _GEN_36429 | _GEN_21463; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25324 = _GEN_36430 | _GEN_21464; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25325 = _GEN_36431 | _GEN_21465; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25326 = _GEN_36432 | _GEN_21466; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_25327 = _GEN_36433 | _GEN_21467; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_25328 = 3'h0 == _T_1647 ? io_op_bits_fn_union : _GEN_25016; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25329 = 3'h1 == _T_1647 ? io_op_bits_fn_union : _GEN_25017; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25330 = 3'h2 == _T_1647 ? io_op_bits_fn_union : _GEN_25018; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25331 = 3'h3 == _T_1647 ? io_op_bits_fn_union : _GEN_25019; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25332 = 3'h4 == _T_1647 ? io_op_bits_fn_union : _GEN_25020; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25333 = 3'h5 == _T_1647 ? io_op_bits_fn_union : _GEN_25021; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25334 = 3'h6 == _T_1647 ? io_op_bits_fn_union : _GEN_25022; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_25335 = 3'h7 == _T_1647 ? io_op_bits_fn_union : _GEN_25023; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_25336 = 3'h0 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24296; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25337 = 3'h1 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24297; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25338 = 3'h2 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24298; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25339 = 3'h3 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24299; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25340 = 3'h4 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24300; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25341 = 3'h5 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24301; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25342 = 3'h6 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24302; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_25343 = 3'h7 == _T_1647 ? io_op_bits_base_vp_id : _GEN_24303; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25344 = 3'h0 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25064; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25345 = 3'h1 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25065; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25346 = 3'h2 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25066; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25347 = 3'h3 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25067; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25348 = 3'h4 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25068; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25349 = 3'h5 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25069; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25350 = 3'h6 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25070; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25351 = 3'h7 == _T_1647 ? io_op_bits_base_vp_valid : _GEN_25071; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25352 = 3'h0 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24312; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25353 = 3'h1 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24313; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25354 = 3'h2 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24314; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25355 = 3'h3 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24315; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25356 = 3'h4 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24316; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25357 = 3'h5 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24317; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25358 = 3'h6 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24318; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25359 = 3'h7 == _T_1647 ? io_op_bits_base_vp_scalar : _GEN_24319; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25360 = 3'h0 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24320; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25361 = 3'h1 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24321; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25362 = 3'h2 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24322; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25363 = 3'h3 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24323; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25364 = 3'h4 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24324; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25365 = 3'h5 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24325; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25366 = 3'h6 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24326; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_25367 = 3'h7 == _T_1647 ? io_op_bits_base_vp_pred : _GEN_24327; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_25368 = 3'h0 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24328; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25369 = 3'h1 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24329; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25370 = 3'h2 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24330; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25371 = 3'h3 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24331; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25372 = 3'h4 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24332; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25373 = 3'h5 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24333; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25374 = 3'h6 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24334; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_25375 = 3'h7 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_24335; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_25376 = io_op_bits_base_vp_valid ? _GEN_25336 : _GEN_24296; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25377 = io_op_bits_base_vp_valid ? _GEN_25337 : _GEN_24297; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25378 = io_op_bits_base_vp_valid ? _GEN_25338 : _GEN_24298; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25379 = io_op_bits_base_vp_valid ? _GEN_25339 : _GEN_24299; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25380 = io_op_bits_base_vp_valid ? _GEN_25340 : _GEN_24300; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25381 = io_op_bits_base_vp_valid ? _GEN_25341 : _GEN_24301; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25382 = io_op_bits_base_vp_valid ? _GEN_25342 : _GEN_24302; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_25383 = io_op_bits_base_vp_valid ? _GEN_25343 : _GEN_24303; // @[sequencer-master.scala 320:41]
  wire  _GEN_25384 = io_op_bits_base_vp_valid ? _GEN_25344 : _GEN_25064; // @[sequencer-master.scala 320:41]
  wire  _GEN_25385 = io_op_bits_base_vp_valid ? _GEN_25345 : _GEN_25065; // @[sequencer-master.scala 320:41]
  wire  _GEN_25386 = io_op_bits_base_vp_valid ? _GEN_25346 : _GEN_25066; // @[sequencer-master.scala 320:41]
  wire  _GEN_25387 = io_op_bits_base_vp_valid ? _GEN_25347 : _GEN_25067; // @[sequencer-master.scala 320:41]
  wire  _GEN_25388 = io_op_bits_base_vp_valid ? _GEN_25348 : _GEN_25068; // @[sequencer-master.scala 320:41]
  wire  _GEN_25389 = io_op_bits_base_vp_valid ? _GEN_25349 : _GEN_25069; // @[sequencer-master.scala 320:41]
  wire  _GEN_25390 = io_op_bits_base_vp_valid ? _GEN_25350 : _GEN_25070; // @[sequencer-master.scala 320:41]
  wire  _GEN_25391 = io_op_bits_base_vp_valid ? _GEN_25351 : _GEN_25071; // @[sequencer-master.scala 320:41]
  wire  _GEN_25392 = io_op_bits_base_vp_valid ? _GEN_25352 : _GEN_24312; // @[sequencer-master.scala 320:41]
  wire  _GEN_25393 = io_op_bits_base_vp_valid ? _GEN_25353 : _GEN_24313; // @[sequencer-master.scala 320:41]
  wire  _GEN_25394 = io_op_bits_base_vp_valid ? _GEN_25354 : _GEN_24314; // @[sequencer-master.scala 320:41]
  wire  _GEN_25395 = io_op_bits_base_vp_valid ? _GEN_25355 : _GEN_24315; // @[sequencer-master.scala 320:41]
  wire  _GEN_25396 = io_op_bits_base_vp_valid ? _GEN_25356 : _GEN_24316; // @[sequencer-master.scala 320:41]
  wire  _GEN_25397 = io_op_bits_base_vp_valid ? _GEN_25357 : _GEN_24317; // @[sequencer-master.scala 320:41]
  wire  _GEN_25398 = io_op_bits_base_vp_valid ? _GEN_25358 : _GEN_24318; // @[sequencer-master.scala 320:41]
  wire  _GEN_25399 = io_op_bits_base_vp_valid ? _GEN_25359 : _GEN_24319; // @[sequencer-master.scala 320:41]
  wire  _GEN_25400 = io_op_bits_base_vp_valid ? _GEN_25360 : _GEN_24320; // @[sequencer-master.scala 320:41]
  wire  _GEN_25401 = io_op_bits_base_vp_valid ? _GEN_25361 : _GEN_24321; // @[sequencer-master.scala 320:41]
  wire  _GEN_25402 = io_op_bits_base_vp_valid ? _GEN_25362 : _GEN_24322; // @[sequencer-master.scala 320:41]
  wire  _GEN_25403 = io_op_bits_base_vp_valid ? _GEN_25363 : _GEN_24323; // @[sequencer-master.scala 320:41]
  wire  _GEN_25404 = io_op_bits_base_vp_valid ? _GEN_25364 : _GEN_24324; // @[sequencer-master.scala 320:41]
  wire  _GEN_25405 = io_op_bits_base_vp_valid ? _GEN_25365 : _GEN_24325; // @[sequencer-master.scala 320:41]
  wire  _GEN_25406 = io_op_bits_base_vp_valid ? _GEN_25366 : _GEN_24326; // @[sequencer-master.scala 320:41]
  wire  _GEN_25407 = io_op_bits_base_vp_valid ? _GEN_25367 : _GEN_24327; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25408 = io_op_bits_base_vp_valid ? _GEN_25368 : _GEN_24328; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25409 = io_op_bits_base_vp_valid ? _GEN_25369 : _GEN_24329; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25410 = io_op_bits_base_vp_valid ? _GEN_25370 : _GEN_24330; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25411 = io_op_bits_base_vp_valid ? _GEN_25371 : _GEN_24331; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25412 = io_op_bits_base_vp_valid ? _GEN_25372 : _GEN_24332; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25413 = io_op_bits_base_vp_valid ? _GEN_25373 : _GEN_24333; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25414 = io_op_bits_base_vp_valid ? _GEN_25374 : _GEN_24334; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_25415 = io_op_bits_base_vp_valid ? _GEN_25375 : _GEN_24335; // @[sequencer-master.scala 320:41]
  wire  _GEN_25416 = _GEN_36426 | _GEN_25112; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25417 = _GEN_36427 | _GEN_25113; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25418 = _GEN_36428 | _GEN_25114; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25419 = _GEN_36429 | _GEN_25115; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25420 = _GEN_36430 | _GEN_25116; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25421 = _GEN_36431 | _GEN_25117; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25422 = _GEN_36432 | _GEN_25118; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25423 = _GEN_36433 | _GEN_25119; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25424 = _T_26 ? _GEN_25416 : _GEN_25112; // @[sequencer-master.scala 154:24]
  wire  _GEN_25425 = _T_26 ? _GEN_25417 : _GEN_25113; // @[sequencer-master.scala 154:24]
  wire  _GEN_25426 = _T_26 ? _GEN_25418 : _GEN_25114; // @[sequencer-master.scala 154:24]
  wire  _GEN_25427 = _T_26 ? _GEN_25419 : _GEN_25115; // @[sequencer-master.scala 154:24]
  wire  _GEN_25428 = _T_26 ? _GEN_25420 : _GEN_25116; // @[sequencer-master.scala 154:24]
  wire  _GEN_25429 = _T_26 ? _GEN_25421 : _GEN_25117; // @[sequencer-master.scala 154:24]
  wire  _GEN_25430 = _T_26 ? _GEN_25422 : _GEN_25118; // @[sequencer-master.scala 154:24]
  wire  _GEN_25431 = _T_26 ? _GEN_25423 : _GEN_25119; // @[sequencer-master.scala 154:24]
  wire  _GEN_25432 = _GEN_36426 | _GEN_25136; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25433 = _GEN_36427 | _GEN_25137; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25434 = _GEN_36428 | _GEN_25138; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25435 = _GEN_36429 | _GEN_25139; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25436 = _GEN_36430 | _GEN_25140; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25437 = _GEN_36431 | _GEN_25141; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25438 = _GEN_36432 | _GEN_25142; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25439 = _GEN_36433 | _GEN_25143; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25440 = _T_48 ? _GEN_25432 : _GEN_25136; // @[sequencer-master.scala 154:24]
  wire  _GEN_25441 = _T_48 ? _GEN_25433 : _GEN_25137; // @[sequencer-master.scala 154:24]
  wire  _GEN_25442 = _T_48 ? _GEN_25434 : _GEN_25138; // @[sequencer-master.scala 154:24]
  wire  _GEN_25443 = _T_48 ? _GEN_25435 : _GEN_25139; // @[sequencer-master.scala 154:24]
  wire  _GEN_25444 = _T_48 ? _GEN_25436 : _GEN_25140; // @[sequencer-master.scala 154:24]
  wire  _GEN_25445 = _T_48 ? _GEN_25437 : _GEN_25141; // @[sequencer-master.scala 154:24]
  wire  _GEN_25446 = _T_48 ? _GEN_25438 : _GEN_25142; // @[sequencer-master.scala 154:24]
  wire  _GEN_25447 = _T_48 ? _GEN_25439 : _GEN_25143; // @[sequencer-master.scala 154:24]
  wire  _GEN_25448 = _GEN_36426 | _GEN_25160; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25449 = _GEN_36427 | _GEN_25161; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25450 = _GEN_36428 | _GEN_25162; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25451 = _GEN_36429 | _GEN_25163; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25452 = _GEN_36430 | _GEN_25164; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25453 = _GEN_36431 | _GEN_25165; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25454 = _GEN_36432 | _GEN_25166; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25455 = _GEN_36433 | _GEN_25167; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25456 = _T_70 ? _GEN_25448 : _GEN_25160; // @[sequencer-master.scala 154:24]
  wire  _GEN_25457 = _T_70 ? _GEN_25449 : _GEN_25161; // @[sequencer-master.scala 154:24]
  wire  _GEN_25458 = _T_70 ? _GEN_25450 : _GEN_25162; // @[sequencer-master.scala 154:24]
  wire  _GEN_25459 = _T_70 ? _GEN_25451 : _GEN_25163; // @[sequencer-master.scala 154:24]
  wire  _GEN_25460 = _T_70 ? _GEN_25452 : _GEN_25164; // @[sequencer-master.scala 154:24]
  wire  _GEN_25461 = _T_70 ? _GEN_25453 : _GEN_25165; // @[sequencer-master.scala 154:24]
  wire  _GEN_25462 = _T_70 ? _GEN_25454 : _GEN_25166; // @[sequencer-master.scala 154:24]
  wire  _GEN_25463 = _T_70 ? _GEN_25455 : _GEN_25167; // @[sequencer-master.scala 154:24]
  wire  _GEN_25464 = _GEN_36426 | _GEN_25184; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25465 = _GEN_36427 | _GEN_25185; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25466 = _GEN_36428 | _GEN_25186; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25467 = _GEN_36429 | _GEN_25187; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25468 = _GEN_36430 | _GEN_25188; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25469 = _GEN_36431 | _GEN_25189; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25470 = _GEN_36432 | _GEN_25190; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25471 = _GEN_36433 | _GEN_25191; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25472 = _T_92 ? _GEN_25464 : _GEN_25184; // @[sequencer-master.scala 154:24]
  wire  _GEN_25473 = _T_92 ? _GEN_25465 : _GEN_25185; // @[sequencer-master.scala 154:24]
  wire  _GEN_25474 = _T_92 ? _GEN_25466 : _GEN_25186; // @[sequencer-master.scala 154:24]
  wire  _GEN_25475 = _T_92 ? _GEN_25467 : _GEN_25187; // @[sequencer-master.scala 154:24]
  wire  _GEN_25476 = _T_92 ? _GEN_25468 : _GEN_25188; // @[sequencer-master.scala 154:24]
  wire  _GEN_25477 = _T_92 ? _GEN_25469 : _GEN_25189; // @[sequencer-master.scala 154:24]
  wire  _GEN_25478 = _T_92 ? _GEN_25470 : _GEN_25190; // @[sequencer-master.scala 154:24]
  wire  _GEN_25479 = _T_92 ? _GEN_25471 : _GEN_25191; // @[sequencer-master.scala 154:24]
  wire  _GEN_25480 = _GEN_36426 | _GEN_25208; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25481 = _GEN_36427 | _GEN_25209; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25482 = _GEN_36428 | _GEN_25210; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25483 = _GEN_36429 | _GEN_25211; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25484 = _GEN_36430 | _GEN_25212; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25485 = _GEN_36431 | _GEN_25213; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25486 = _GEN_36432 | _GEN_25214; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25487 = _GEN_36433 | _GEN_25215; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25488 = _T_114 ? _GEN_25480 : _GEN_25208; // @[sequencer-master.scala 154:24]
  wire  _GEN_25489 = _T_114 ? _GEN_25481 : _GEN_25209; // @[sequencer-master.scala 154:24]
  wire  _GEN_25490 = _T_114 ? _GEN_25482 : _GEN_25210; // @[sequencer-master.scala 154:24]
  wire  _GEN_25491 = _T_114 ? _GEN_25483 : _GEN_25211; // @[sequencer-master.scala 154:24]
  wire  _GEN_25492 = _T_114 ? _GEN_25484 : _GEN_25212; // @[sequencer-master.scala 154:24]
  wire  _GEN_25493 = _T_114 ? _GEN_25485 : _GEN_25213; // @[sequencer-master.scala 154:24]
  wire  _GEN_25494 = _T_114 ? _GEN_25486 : _GEN_25214; // @[sequencer-master.scala 154:24]
  wire  _GEN_25495 = _T_114 ? _GEN_25487 : _GEN_25215; // @[sequencer-master.scala 154:24]
  wire  _GEN_25496 = _GEN_36426 | _GEN_25232; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25497 = _GEN_36427 | _GEN_25233; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25498 = _GEN_36428 | _GEN_25234; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25499 = _GEN_36429 | _GEN_25235; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25500 = _GEN_36430 | _GEN_25236; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25501 = _GEN_36431 | _GEN_25237; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25502 = _GEN_36432 | _GEN_25238; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25503 = _GEN_36433 | _GEN_25239; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25504 = _T_136 ? _GEN_25496 : _GEN_25232; // @[sequencer-master.scala 154:24]
  wire  _GEN_25505 = _T_136 ? _GEN_25497 : _GEN_25233; // @[sequencer-master.scala 154:24]
  wire  _GEN_25506 = _T_136 ? _GEN_25498 : _GEN_25234; // @[sequencer-master.scala 154:24]
  wire  _GEN_25507 = _T_136 ? _GEN_25499 : _GEN_25235; // @[sequencer-master.scala 154:24]
  wire  _GEN_25508 = _T_136 ? _GEN_25500 : _GEN_25236; // @[sequencer-master.scala 154:24]
  wire  _GEN_25509 = _T_136 ? _GEN_25501 : _GEN_25237; // @[sequencer-master.scala 154:24]
  wire  _GEN_25510 = _T_136 ? _GEN_25502 : _GEN_25238; // @[sequencer-master.scala 154:24]
  wire  _GEN_25511 = _T_136 ? _GEN_25503 : _GEN_25239; // @[sequencer-master.scala 154:24]
  wire  _GEN_25512 = _GEN_36426 | _GEN_25256; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25513 = _GEN_36427 | _GEN_25257; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25514 = _GEN_36428 | _GEN_25258; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25515 = _GEN_36429 | _GEN_25259; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25516 = _GEN_36430 | _GEN_25260; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25517 = _GEN_36431 | _GEN_25261; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25518 = _GEN_36432 | _GEN_25262; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25519 = _GEN_36433 | _GEN_25263; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25520 = _T_158 ? _GEN_25512 : _GEN_25256; // @[sequencer-master.scala 154:24]
  wire  _GEN_25521 = _T_158 ? _GEN_25513 : _GEN_25257; // @[sequencer-master.scala 154:24]
  wire  _GEN_25522 = _T_158 ? _GEN_25514 : _GEN_25258; // @[sequencer-master.scala 154:24]
  wire  _GEN_25523 = _T_158 ? _GEN_25515 : _GEN_25259; // @[sequencer-master.scala 154:24]
  wire  _GEN_25524 = _T_158 ? _GEN_25516 : _GEN_25260; // @[sequencer-master.scala 154:24]
  wire  _GEN_25525 = _T_158 ? _GEN_25517 : _GEN_25261; // @[sequencer-master.scala 154:24]
  wire  _GEN_25526 = _T_158 ? _GEN_25518 : _GEN_25262; // @[sequencer-master.scala 154:24]
  wire  _GEN_25527 = _T_158 ? _GEN_25519 : _GEN_25263; // @[sequencer-master.scala 154:24]
  wire  _GEN_25528 = _GEN_36426 | _GEN_25280; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25529 = _GEN_36427 | _GEN_25281; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25530 = _GEN_36428 | _GEN_25282; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25531 = _GEN_36429 | _GEN_25283; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25532 = _GEN_36430 | _GEN_25284; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25533 = _GEN_36431 | _GEN_25285; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25534 = _GEN_36432 | _GEN_25286; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25535 = _GEN_36433 | _GEN_25287; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25536 = _T_180 ? _GEN_25528 : _GEN_25280; // @[sequencer-master.scala 154:24]
  wire  _GEN_25537 = _T_180 ? _GEN_25529 : _GEN_25281; // @[sequencer-master.scala 154:24]
  wire  _GEN_25538 = _T_180 ? _GEN_25530 : _GEN_25282; // @[sequencer-master.scala 154:24]
  wire  _GEN_25539 = _T_180 ? _GEN_25531 : _GEN_25283; // @[sequencer-master.scala 154:24]
  wire  _GEN_25540 = _T_180 ? _GEN_25532 : _GEN_25284; // @[sequencer-master.scala 154:24]
  wire  _GEN_25541 = _T_180 ? _GEN_25533 : _GEN_25285; // @[sequencer-master.scala 154:24]
  wire  _GEN_25542 = _T_180 ? _GEN_25534 : _GEN_25286; // @[sequencer-master.scala 154:24]
  wire  _GEN_25543 = _T_180 ? _GEN_25535 : _GEN_25287; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_25544 = 3'h0 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24528; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25545 = 3'h1 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24529; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25546 = 3'h2 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24530; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25547 = 3'h3 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24531; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25548 = 3'h4 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24532; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25549 = 3'h5 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24533; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25550 = 3'h6 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24534; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25551 = 3'h7 == _T_1647 ? io_op_bits_base_vd_id : _GEN_24535; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25552 = 3'h0 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25072; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25553 = 3'h1 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25073; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25554 = 3'h2 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25074; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25555 = 3'h3 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25075; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25556 = 3'h4 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25076; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25557 = 3'h5 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25077; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25558 = 3'h6 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25078; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25559 = 3'h7 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_25079; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25560 = 3'h0 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24544; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25561 = 3'h1 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24545; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25562 = 3'h2 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24546; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25563 = 3'h3 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24547; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25564 = 3'h4 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24548; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25565 = 3'h5 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24549; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25566 = 3'h6 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24550; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25567 = 3'h7 == _T_1647 ? io_op_bits_base_vd_scalar : _GEN_24551; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25568 = 3'h0 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24552; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25569 = 3'h1 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24553; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25570 = 3'h2 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24554; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25571 = 3'h3 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24555; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25572 = 3'h4 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24556; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25573 = 3'h5 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24557; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25574 = 3'h6 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24558; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire  _GEN_25575 = 3'h7 == _T_1647 ? io_op_bits_base_vd_pred : _GEN_24559; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25576 = 3'h0 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24560; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25577 = 3'h1 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24561; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25578 = 3'h2 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24562; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25579 = 3'h3 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24563; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25580 = 3'h4 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24564; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25581 = 3'h5 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24565; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25582 = 3'h6 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24566; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [1:0] _GEN_25583 = 3'h7 == _T_1647 ? io_op_bits_base_vd_prec : _GEN_24567; // @[sequencer-master.scala 355:25 sequencer-master.scala 355:25]
  wire [7:0] _GEN_25584 = 3'h0 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24568; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25585 = 3'h1 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24569; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25586 = 3'h2 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24570; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25587 = 3'h3 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24571; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25588 = 3'h4 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24572; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25589 = 3'h5 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24573; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25590 = 3'h6 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24574; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25591 = 3'h7 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_24575; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_25592 = io_op_bits_base_vd_valid ? _GEN_25544 : _GEN_24528; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25593 = io_op_bits_base_vd_valid ? _GEN_25545 : _GEN_24529; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25594 = io_op_bits_base_vd_valid ? _GEN_25546 : _GEN_24530; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25595 = io_op_bits_base_vd_valid ? _GEN_25547 : _GEN_24531; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25596 = io_op_bits_base_vd_valid ? _GEN_25548 : _GEN_24532; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25597 = io_op_bits_base_vd_valid ? _GEN_25549 : _GEN_24533; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25598 = io_op_bits_base_vd_valid ? _GEN_25550 : _GEN_24534; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25599 = io_op_bits_base_vd_valid ? _GEN_25551 : _GEN_24535; // @[sequencer-master.scala 354:41]
  wire  _GEN_25600 = io_op_bits_base_vd_valid ? _GEN_25552 : _GEN_25072; // @[sequencer-master.scala 354:41]
  wire  _GEN_25601 = io_op_bits_base_vd_valid ? _GEN_25553 : _GEN_25073; // @[sequencer-master.scala 354:41]
  wire  _GEN_25602 = io_op_bits_base_vd_valid ? _GEN_25554 : _GEN_25074; // @[sequencer-master.scala 354:41]
  wire  _GEN_25603 = io_op_bits_base_vd_valid ? _GEN_25555 : _GEN_25075; // @[sequencer-master.scala 354:41]
  wire  _GEN_25604 = io_op_bits_base_vd_valid ? _GEN_25556 : _GEN_25076; // @[sequencer-master.scala 354:41]
  wire  _GEN_25605 = io_op_bits_base_vd_valid ? _GEN_25557 : _GEN_25077; // @[sequencer-master.scala 354:41]
  wire  _GEN_25606 = io_op_bits_base_vd_valid ? _GEN_25558 : _GEN_25078; // @[sequencer-master.scala 354:41]
  wire  _GEN_25607 = io_op_bits_base_vd_valid ? _GEN_25559 : _GEN_25079; // @[sequencer-master.scala 354:41]
  wire  _GEN_25608 = io_op_bits_base_vd_valid ? _GEN_25560 : _GEN_24544; // @[sequencer-master.scala 354:41]
  wire  _GEN_25609 = io_op_bits_base_vd_valid ? _GEN_25561 : _GEN_24545; // @[sequencer-master.scala 354:41]
  wire  _GEN_25610 = io_op_bits_base_vd_valid ? _GEN_25562 : _GEN_24546; // @[sequencer-master.scala 354:41]
  wire  _GEN_25611 = io_op_bits_base_vd_valid ? _GEN_25563 : _GEN_24547; // @[sequencer-master.scala 354:41]
  wire  _GEN_25612 = io_op_bits_base_vd_valid ? _GEN_25564 : _GEN_24548; // @[sequencer-master.scala 354:41]
  wire  _GEN_25613 = io_op_bits_base_vd_valid ? _GEN_25565 : _GEN_24549; // @[sequencer-master.scala 354:41]
  wire  _GEN_25614 = io_op_bits_base_vd_valid ? _GEN_25566 : _GEN_24550; // @[sequencer-master.scala 354:41]
  wire  _GEN_25615 = io_op_bits_base_vd_valid ? _GEN_25567 : _GEN_24551; // @[sequencer-master.scala 354:41]
  wire  _GEN_25616 = io_op_bits_base_vd_valid ? _GEN_25568 : _GEN_24552; // @[sequencer-master.scala 354:41]
  wire  _GEN_25617 = io_op_bits_base_vd_valid ? _GEN_25569 : _GEN_24553; // @[sequencer-master.scala 354:41]
  wire  _GEN_25618 = io_op_bits_base_vd_valid ? _GEN_25570 : _GEN_24554; // @[sequencer-master.scala 354:41]
  wire  _GEN_25619 = io_op_bits_base_vd_valid ? _GEN_25571 : _GEN_24555; // @[sequencer-master.scala 354:41]
  wire  _GEN_25620 = io_op_bits_base_vd_valid ? _GEN_25572 : _GEN_24556; // @[sequencer-master.scala 354:41]
  wire  _GEN_25621 = io_op_bits_base_vd_valid ? _GEN_25573 : _GEN_24557; // @[sequencer-master.scala 354:41]
  wire  _GEN_25622 = io_op_bits_base_vd_valid ? _GEN_25574 : _GEN_24558; // @[sequencer-master.scala 354:41]
  wire  _GEN_25623 = io_op_bits_base_vd_valid ? _GEN_25575 : _GEN_24559; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25624 = io_op_bits_base_vd_valid ? _GEN_25576 : _GEN_24560; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25625 = io_op_bits_base_vd_valid ? _GEN_25577 : _GEN_24561; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25626 = io_op_bits_base_vd_valid ? _GEN_25578 : _GEN_24562; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25627 = io_op_bits_base_vd_valid ? _GEN_25579 : _GEN_24563; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25628 = io_op_bits_base_vd_valid ? _GEN_25580 : _GEN_24564; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25629 = io_op_bits_base_vd_valid ? _GEN_25581 : _GEN_24565; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25630 = io_op_bits_base_vd_valid ? _GEN_25582 : _GEN_24566; // @[sequencer-master.scala 354:41]
  wire [1:0] _GEN_25631 = io_op_bits_base_vd_valid ? _GEN_25583 : _GEN_24567; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25632 = io_op_bits_base_vd_valid ? _GEN_25584 : _GEN_24568; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25633 = io_op_bits_base_vd_valid ? _GEN_25585 : _GEN_24569; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25634 = io_op_bits_base_vd_valid ? _GEN_25586 : _GEN_24570; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25635 = io_op_bits_base_vd_valid ? _GEN_25587 : _GEN_24571; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25636 = io_op_bits_base_vd_valid ? _GEN_25588 : _GEN_24572; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25637 = io_op_bits_base_vd_valid ? _GEN_25589 : _GEN_24573; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25638 = io_op_bits_base_vd_valid ? _GEN_25590 : _GEN_24574; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_25639 = io_op_bits_base_vd_valid ? _GEN_25591 : _GEN_24575; // @[sequencer-master.scala 354:41]
  wire  _GEN_25640 = _GEN_36426 | _GEN_25424; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25641 = _GEN_36427 | _GEN_25425; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25642 = _GEN_36428 | _GEN_25426; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25643 = _GEN_36429 | _GEN_25427; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25644 = _GEN_36430 | _GEN_25428; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25645 = _GEN_36431 | _GEN_25429; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25646 = _GEN_36432 | _GEN_25430; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25647 = _GEN_36433 | _GEN_25431; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25648 = _T_1442 ? _GEN_25640 : _GEN_25424; // @[sequencer-master.scala 154:24]
  wire  _GEN_25649 = _T_1442 ? _GEN_25641 : _GEN_25425; // @[sequencer-master.scala 154:24]
  wire  _GEN_25650 = _T_1442 ? _GEN_25642 : _GEN_25426; // @[sequencer-master.scala 154:24]
  wire  _GEN_25651 = _T_1442 ? _GEN_25643 : _GEN_25427; // @[sequencer-master.scala 154:24]
  wire  _GEN_25652 = _T_1442 ? _GEN_25644 : _GEN_25428; // @[sequencer-master.scala 154:24]
  wire  _GEN_25653 = _T_1442 ? _GEN_25645 : _GEN_25429; // @[sequencer-master.scala 154:24]
  wire  _GEN_25654 = _T_1442 ? _GEN_25646 : _GEN_25430; // @[sequencer-master.scala 154:24]
  wire  _GEN_25655 = _T_1442 ? _GEN_25647 : _GEN_25431; // @[sequencer-master.scala 154:24]
  wire  _GEN_25656 = _GEN_36426 | _GEN_25440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25657 = _GEN_36427 | _GEN_25441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25658 = _GEN_36428 | _GEN_25442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25659 = _GEN_36429 | _GEN_25443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25660 = _GEN_36430 | _GEN_25444; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25661 = _GEN_36431 | _GEN_25445; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25662 = _GEN_36432 | _GEN_25446; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25663 = _GEN_36433 | _GEN_25447; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25664 = _T_1464 ? _GEN_25656 : _GEN_25440; // @[sequencer-master.scala 154:24]
  wire  _GEN_25665 = _T_1464 ? _GEN_25657 : _GEN_25441; // @[sequencer-master.scala 154:24]
  wire  _GEN_25666 = _T_1464 ? _GEN_25658 : _GEN_25442; // @[sequencer-master.scala 154:24]
  wire  _GEN_25667 = _T_1464 ? _GEN_25659 : _GEN_25443; // @[sequencer-master.scala 154:24]
  wire  _GEN_25668 = _T_1464 ? _GEN_25660 : _GEN_25444; // @[sequencer-master.scala 154:24]
  wire  _GEN_25669 = _T_1464 ? _GEN_25661 : _GEN_25445; // @[sequencer-master.scala 154:24]
  wire  _GEN_25670 = _T_1464 ? _GEN_25662 : _GEN_25446; // @[sequencer-master.scala 154:24]
  wire  _GEN_25671 = _T_1464 ? _GEN_25663 : _GEN_25447; // @[sequencer-master.scala 154:24]
  wire  _GEN_25672 = _GEN_36426 | _GEN_25456; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25673 = _GEN_36427 | _GEN_25457; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25674 = _GEN_36428 | _GEN_25458; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25675 = _GEN_36429 | _GEN_25459; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25676 = _GEN_36430 | _GEN_25460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25677 = _GEN_36431 | _GEN_25461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25678 = _GEN_36432 | _GEN_25462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25679 = _GEN_36433 | _GEN_25463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25680 = _T_1486 ? _GEN_25672 : _GEN_25456; // @[sequencer-master.scala 154:24]
  wire  _GEN_25681 = _T_1486 ? _GEN_25673 : _GEN_25457; // @[sequencer-master.scala 154:24]
  wire  _GEN_25682 = _T_1486 ? _GEN_25674 : _GEN_25458; // @[sequencer-master.scala 154:24]
  wire  _GEN_25683 = _T_1486 ? _GEN_25675 : _GEN_25459; // @[sequencer-master.scala 154:24]
  wire  _GEN_25684 = _T_1486 ? _GEN_25676 : _GEN_25460; // @[sequencer-master.scala 154:24]
  wire  _GEN_25685 = _T_1486 ? _GEN_25677 : _GEN_25461; // @[sequencer-master.scala 154:24]
  wire  _GEN_25686 = _T_1486 ? _GEN_25678 : _GEN_25462; // @[sequencer-master.scala 154:24]
  wire  _GEN_25687 = _T_1486 ? _GEN_25679 : _GEN_25463; // @[sequencer-master.scala 154:24]
  wire  _GEN_25688 = _GEN_36426 | _GEN_25472; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25689 = _GEN_36427 | _GEN_25473; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25690 = _GEN_36428 | _GEN_25474; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25691 = _GEN_36429 | _GEN_25475; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25692 = _GEN_36430 | _GEN_25476; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25693 = _GEN_36431 | _GEN_25477; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25694 = _GEN_36432 | _GEN_25478; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25695 = _GEN_36433 | _GEN_25479; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25696 = _T_1508 ? _GEN_25688 : _GEN_25472; // @[sequencer-master.scala 154:24]
  wire  _GEN_25697 = _T_1508 ? _GEN_25689 : _GEN_25473; // @[sequencer-master.scala 154:24]
  wire  _GEN_25698 = _T_1508 ? _GEN_25690 : _GEN_25474; // @[sequencer-master.scala 154:24]
  wire  _GEN_25699 = _T_1508 ? _GEN_25691 : _GEN_25475; // @[sequencer-master.scala 154:24]
  wire  _GEN_25700 = _T_1508 ? _GEN_25692 : _GEN_25476; // @[sequencer-master.scala 154:24]
  wire  _GEN_25701 = _T_1508 ? _GEN_25693 : _GEN_25477; // @[sequencer-master.scala 154:24]
  wire  _GEN_25702 = _T_1508 ? _GEN_25694 : _GEN_25478; // @[sequencer-master.scala 154:24]
  wire  _GEN_25703 = _T_1508 ? _GEN_25695 : _GEN_25479; // @[sequencer-master.scala 154:24]
  wire  _GEN_25704 = _GEN_36426 | _GEN_25488; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25705 = _GEN_36427 | _GEN_25489; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25706 = _GEN_36428 | _GEN_25490; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25707 = _GEN_36429 | _GEN_25491; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25708 = _GEN_36430 | _GEN_25492; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25709 = _GEN_36431 | _GEN_25493; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25710 = _GEN_36432 | _GEN_25494; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25711 = _GEN_36433 | _GEN_25495; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25712 = _T_1530 ? _GEN_25704 : _GEN_25488; // @[sequencer-master.scala 154:24]
  wire  _GEN_25713 = _T_1530 ? _GEN_25705 : _GEN_25489; // @[sequencer-master.scala 154:24]
  wire  _GEN_25714 = _T_1530 ? _GEN_25706 : _GEN_25490; // @[sequencer-master.scala 154:24]
  wire  _GEN_25715 = _T_1530 ? _GEN_25707 : _GEN_25491; // @[sequencer-master.scala 154:24]
  wire  _GEN_25716 = _T_1530 ? _GEN_25708 : _GEN_25492; // @[sequencer-master.scala 154:24]
  wire  _GEN_25717 = _T_1530 ? _GEN_25709 : _GEN_25493; // @[sequencer-master.scala 154:24]
  wire  _GEN_25718 = _T_1530 ? _GEN_25710 : _GEN_25494; // @[sequencer-master.scala 154:24]
  wire  _GEN_25719 = _T_1530 ? _GEN_25711 : _GEN_25495; // @[sequencer-master.scala 154:24]
  wire  _GEN_25720 = _GEN_36426 | _GEN_25504; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25721 = _GEN_36427 | _GEN_25505; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25722 = _GEN_36428 | _GEN_25506; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25723 = _GEN_36429 | _GEN_25507; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25724 = _GEN_36430 | _GEN_25508; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25725 = _GEN_36431 | _GEN_25509; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25726 = _GEN_36432 | _GEN_25510; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25727 = _GEN_36433 | _GEN_25511; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25728 = _T_1552 ? _GEN_25720 : _GEN_25504; // @[sequencer-master.scala 154:24]
  wire  _GEN_25729 = _T_1552 ? _GEN_25721 : _GEN_25505; // @[sequencer-master.scala 154:24]
  wire  _GEN_25730 = _T_1552 ? _GEN_25722 : _GEN_25506; // @[sequencer-master.scala 154:24]
  wire  _GEN_25731 = _T_1552 ? _GEN_25723 : _GEN_25507; // @[sequencer-master.scala 154:24]
  wire  _GEN_25732 = _T_1552 ? _GEN_25724 : _GEN_25508; // @[sequencer-master.scala 154:24]
  wire  _GEN_25733 = _T_1552 ? _GEN_25725 : _GEN_25509; // @[sequencer-master.scala 154:24]
  wire  _GEN_25734 = _T_1552 ? _GEN_25726 : _GEN_25510; // @[sequencer-master.scala 154:24]
  wire  _GEN_25735 = _T_1552 ? _GEN_25727 : _GEN_25511; // @[sequencer-master.scala 154:24]
  wire  _GEN_25736 = _GEN_36426 | _GEN_25520; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25737 = _GEN_36427 | _GEN_25521; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25738 = _GEN_36428 | _GEN_25522; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25739 = _GEN_36429 | _GEN_25523; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25740 = _GEN_36430 | _GEN_25524; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25741 = _GEN_36431 | _GEN_25525; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25742 = _GEN_36432 | _GEN_25526; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25743 = _GEN_36433 | _GEN_25527; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25744 = _T_1574 ? _GEN_25736 : _GEN_25520; // @[sequencer-master.scala 154:24]
  wire  _GEN_25745 = _T_1574 ? _GEN_25737 : _GEN_25521; // @[sequencer-master.scala 154:24]
  wire  _GEN_25746 = _T_1574 ? _GEN_25738 : _GEN_25522; // @[sequencer-master.scala 154:24]
  wire  _GEN_25747 = _T_1574 ? _GEN_25739 : _GEN_25523; // @[sequencer-master.scala 154:24]
  wire  _GEN_25748 = _T_1574 ? _GEN_25740 : _GEN_25524; // @[sequencer-master.scala 154:24]
  wire  _GEN_25749 = _T_1574 ? _GEN_25741 : _GEN_25525; // @[sequencer-master.scala 154:24]
  wire  _GEN_25750 = _T_1574 ? _GEN_25742 : _GEN_25526; // @[sequencer-master.scala 154:24]
  wire  _GEN_25751 = _T_1574 ? _GEN_25743 : _GEN_25527; // @[sequencer-master.scala 154:24]
  wire  _GEN_25752 = _GEN_36426 | _GEN_25536; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25753 = _GEN_36427 | _GEN_25537; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25754 = _GEN_36428 | _GEN_25538; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25755 = _GEN_36429 | _GEN_25539; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25756 = _GEN_36430 | _GEN_25540; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25757 = _GEN_36431 | _GEN_25541; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25758 = _GEN_36432 | _GEN_25542; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25759 = _GEN_36433 | _GEN_25543; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25760 = _T_1596 ? _GEN_25752 : _GEN_25536; // @[sequencer-master.scala 154:24]
  wire  _GEN_25761 = _T_1596 ? _GEN_25753 : _GEN_25537; // @[sequencer-master.scala 154:24]
  wire  _GEN_25762 = _T_1596 ? _GEN_25754 : _GEN_25538; // @[sequencer-master.scala 154:24]
  wire  _GEN_25763 = _T_1596 ? _GEN_25755 : _GEN_25539; // @[sequencer-master.scala 154:24]
  wire  _GEN_25764 = _T_1596 ? _GEN_25756 : _GEN_25540; // @[sequencer-master.scala 154:24]
  wire  _GEN_25765 = _T_1596 ? _GEN_25757 : _GEN_25541; // @[sequencer-master.scala 154:24]
  wire  _GEN_25766 = _T_1596 ? _GEN_25758 : _GEN_25542; // @[sequencer-master.scala 154:24]
  wire  _GEN_25767 = _T_1596 ? _GEN_25759 : _GEN_25543; // @[sequencer-master.scala 154:24]
  wire [1:0] _e_T_1647_rports_1 = {{1'd0}, _T_1639}; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25768 = 3'h0 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25024; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25769 = 3'h1 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25025; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25770 = 3'h2 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25026; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25771 = 3'h3 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25027; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25772 = 3'h4 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25028; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25773 = 3'h5 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25029; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25774 = 3'h6 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25030; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_25775 = 3'h7 == _T_1647 ? _e_T_1647_rports_1 : _GEN_25031; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_25776 = 3'h0 == _T_1647 ? 4'h0 : _GEN_25032; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25777 = 3'h1 == _T_1647 ? 4'h0 : _GEN_25033; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25778 = 3'h2 == _T_1647 ? 4'h0 : _GEN_25034; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25779 = 3'h3 == _T_1647 ? 4'h0 : _GEN_25035; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25780 = 3'h4 == _T_1647 ? 4'h0 : _GEN_25036; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25781 = 3'h5 == _T_1647 ? 4'h0 : _GEN_25037; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25782 = 3'h6 == _T_1647 ? 4'h0 : _GEN_25038; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_25783 = 3'h7 == _T_1647 ? 4'h0 : _GEN_25039; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_25784 = 3'h0 == _T_1647 ? 3'h0 : _GEN_25040; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25785 = 3'h1 == _T_1647 ? 3'h0 : _GEN_25041; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25786 = 3'h2 == _T_1647 ? 3'h0 : _GEN_25042; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25787 = 3'h3 == _T_1647 ? 3'h0 : _GEN_25043; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25788 = 3'h4 == _T_1647 ? 3'h0 : _GEN_25044; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25789 = 3'h5 == _T_1647 ? 3'h0 : _GEN_25045; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25790 = 3'h6 == _T_1647 ? 3'h0 : _GEN_25046; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_25791 = 3'h7 == _T_1647 ? 3'h0 : _GEN_25047; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_25792 = _GEN_36426 & _GEN_34121 | _GEN_25648; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25793 = _GEN_36426 & _GEN_34122 | _GEN_25664; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25794 = _GEN_36426 & _GEN_34123 | _GEN_25680; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25795 = _GEN_36426 & _GEN_34124 | _GEN_25696; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25796 = _GEN_36426 & _GEN_34125 | _GEN_25712; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25797 = _GEN_36426 & _GEN_34126 | _GEN_25728; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25798 = _GEN_36426 & _GEN_34127 | _GEN_25744; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25799 = _GEN_36426 & _GEN_34128 | _GEN_25760; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25800 = _GEN_36427 & _GEN_34121 | _GEN_25649; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25801 = _GEN_36427 & _GEN_34122 | _GEN_25665; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25802 = _GEN_36427 & _GEN_34123 | _GEN_25681; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25803 = _GEN_36427 & _GEN_34124 | _GEN_25697; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25804 = _GEN_36427 & _GEN_34125 | _GEN_25713; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25805 = _GEN_36427 & _GEN_34126 | _GEN_25729; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25806 = _GEN_36427 & _GEN_34127 | _GEN_25745; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25807 = _GEN_36427 & _GEN_34128 | _GEN_25761; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25808 = _GEN_36428 & _GEN_34121 | _GEN_25650; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25809 = _GEN_36428 & _GEN_34122 | _GEN_25666; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25810 = _GEN_36428 & _GEN_34123 | _GEN_25682; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25811 = _GEN_36428 & _GEN_34124 | _GEN_25698; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25812 = _GEN_36428 & _GEN_34125 | _GEN_25714; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25813 = _GEN_36428 & _GEN_34126 | _GEN_25730; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25814 = _GEN_36428 & _GEN_34127 | _GEN_25746; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25815 = _GEN_36428 & _GEN_34128 | _GEN_25762; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25816 = _GEN_36429 & _GEN_34121 | _GEN_25651; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25817 = _GEN_36429 & _GEN_34122 | _GEN_25667; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25818 = _GEN_36429 & _GEN_34123 | _GEN_25683; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25819 = _GEN_36429 & _GEN_34124 | _GEN_25699; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25820 = _GEN_36429 & _GEN_34125 | _GEN_25715; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25821 = _GEN_36429 & _GEN_34126 | _GEN_25731; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25822 = _GEN_36429 & _GEN_34127 | _GEN_25747; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25823 = _GEN_36429 & _GEN_34128 | _GEN_25763; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25824 = _GEN_36430 & _GEN_34121 | _GEN_25652; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25825 = _GEN_36430 & _GEN_34122 | _GEN_25668; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25826 = _GEN_36430 & _GEN_34123 | _GEN_25684; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25827 = _GEN_36430 & _GEN_34124 | _GEN_25700; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25828 = _GEN_36430 & _GEN_34125 | _GEN_25716; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25829 = _GEN_36430 & _GEN_34126 | _GEN_25732; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25830 = _GEN_36430 & _GEN_34127 | _GEN_25748; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25831 = _GEN_36430 & _GEN_34128 | _GEN_25764; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25832 = _GEN_36431 & _GEN_34121 | _GEN_25653; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25833 = _GEN_36431 & _GEN_34122 | _GEN_25669; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25834 = _GEN_36431 & _GEN_34123 | _GEN_25685; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25835 = _GEN_36431 & _GEN_34124 | _GEN_25701; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25836 = _GEN_36431 & _GEN_34125 | _GEN_25717; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25837 = _GEN_36431 & _GEN_34126 | _GEN_25733; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25838 = _GEN_36431 & _GEN_34127 | _GEN_25749; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25839 = _GEN_36431 & _GEN_34128 | _GEN_25765; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25840 = _GEN_36432 & _GEN_34121 | _GEN_25654; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25841 = _GEN_36432 & _GEN_34122 | _GEN_25670; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25842 = _GEN_36432 & _GEN_34123 | _GEN_25686; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25843 = _GEN_36432 & _GEN_34124 | _GEN_25702; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25844 = _GEN_36432 & _GEN_34125 | _GEN_25718; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25845 = _GEN_36432 & _GEN_34126 | _GEN_25734; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25846 = _GEN_36432 & _GEN_34127 | _GEN_25750; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25847 = _GEN_36432 & _GEN_34128 | _GEN_25766; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25848 = _GEN_36433 & _GEN_34121 | _GEN_25655; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25849 = _GEN_36433 & _GEN_34122 | _GEN_25671; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25850 = _GEN_36433 & _GEN_34123 | _GEN_25687; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25851 = _GEN_36433 & _GEN_34124 | _GEN_25703; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25852 = _GEN_36433 & _GEN_34125 | _GEN_25719; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25853 = _GEN_36433 & _GEN_34126 | _GEN_25735; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25854 = _GEN_36433 & _GEN_34127 | _GEN_25751; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25855 = _GEN_36433 & _GEN_34128 | _GEN_25767; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_25856 = io_op_bits_active_vstx ? _GEN_25048 : _GEN_23518; // @[sequencer-master.scala 652:39]
  wire  _GEN_25857 = io_op_bits_active_vstx ? _GEN_25049 : _GEN_23519; // @[sequencer-master.scala 652:39]
  wire  _GEN_25858 = io_op_bits_active_vstx ? _GEN_25050 : _GEN_23520; // @[sequencer-master.scala 652:39]
  wire  _GEN_25859 = io_op_bits_active_vstx ? _GEN_25051 : _GEN_23521; // @[sequencer-master.scala 652:39]
  wire  _GEN_25860 = io_op_bits_active_vstx ? _GEN_25052 : _GEN_23522; // @[sequencer-master.scala 652:39]
  wire  _GEN_25861 = io_op_bits_active_vstx ? _GEN_25053 : _GEN_23523; // @[sequencer-master.scala 652:39]
  wire  _GEN_25862 = io_op_bits_active_vstx ? _GEN_25054 : _GEN_23524; // @[sequencer-master.scala 652:39]
  wire  _GEN_25863 = io_op_bits_active_vstx ? _GEN_25055 : _GEN_23525; // @[sequencer-master.scala 652:39]
  wire  _GEN_25872 = io_op_bits_active_vstx ? _GEN_25384 : _GEN_23534; // @[sequencer-master.scala 652:39]
  wire  _GEN_25873 = io_op_bits_active_vstx ? _GEN_25385 : _GEN_23535; // @[sequencer-master.scala 652:39]
  wire  _GEN_25874 = io_op_bits_active_vstx ? _GEN_25386 : _GEN_23536; // @[sequencer-master.scala 652:39]
  wire  _GEN_25875 = io_op_bits_active_vstx ? _GEN_25387 : _GEN_23537; // @[sequencer-master.scala 652:39]
  wire  _GEN_25876 = io_op_bits_active_vstx ? _GEN_25388 : _GEN_23538; // @[sequencer-master.scala 652:39]
  wire  _GEN_25877 = io_op_bits_active_vstx ? _GEN_25389 : _GEN_23539; // @[sequencer-master.scala 652:39]
  wire  _GEN_25878 = io_op_bits_active_vstx ? _GEN_25390 : _GEN_23540; // @[sequencer-master.scala 652:39]
  wire  _GEN_25879 = io_op_bits_active_vstx ? _GEN_25391 : _GEN_23541; // @[sequencer-master.scala 652:39]
  wire  _GEN_25880 = io_op_bits_active_vstx ? _GEN_25600 : _GEN_23542; // @[sequencer-master.scala 652:39]
  wire  _GEN_25881 = io_op_bits_active_vstx ? _GEN_25601 : _GEN_23543; // @[sequencer-master.scala 652:39]
  wire  _GEN_25882 = io_op_bits_active_vstx ? _GEN_25602 : _GEN_23544; // @[sequencer-master.scala 652:39]
  wire  _GEN_25883 = io_op_bits_active_vstx ? _GEN_25603 : _GEN_23545; // @[sequencer-master.scala 652:39]
  wire  _GEN_25884 = io_op_bits_active_vstx ? _GEN_25604 : _GEN_23546; // @[sequencer-master.scala 652:39]
  wire  _GEN_25885 = io_op_bits_active_vstx ? _GEN_25605 : _GEN_23547; // @[sequencer-master.scala 652:39]
  wire  _GEN_25886 = io_op_bits_active_vstx ? _GEN_25606 : _GEN_23548; // @[sequencer-master.scala 652:39]
  wire  _GEN_25887 = io_op_bits_active_vstx ? _GEN_25607 : _GEN_23549; // @[sequencer-master.scala 652:39]
  wire  _GEN_25888 = io_op_bits_active_vstx ? _GEN_25080 : _GEN_23550; // @[sequencer-master.scala 652:39]
  wire  _GEN_25889 = io_op_bits_active_vstx ? _GEN_25081 : _GEN_23551; // @[sequencer-master.scala 652:39]
  wire  _GEN_25890 = io_op_bits_active_vstx ? _GEN_25082 : _GEN_23552; // @[sequencer-master.scala 652:39]
  wire  _GEN_25891 = io_op_bits_active_vstx ? _GEN_25083 : _GEN_23553; // @[sequencer-master.scala 652:39]
  wire  _GEN_25892 = io_op_bits_active_vstx ? _GEN_25084 : _GEN_23554; // @[sequencer-master.scala 652:39]
  wire  _GEN_25893 = io_op_bits_active_vstx ? _GEN_25085 : _GEN_23555; // @[sequencer-master.scala 652:39]
  wire  _GEN_25894 = io_op_bits_active_vstx ? _GEN_25086 : _GEN_23556; // @[sequencer-master.scala 652:39]
  wire  _GEN_25895 = io_op_bits_active_vstx ? _GEN_25087 : _GEN_23557; // @[sequencer-master.scala 652:39]
  wire  _GEN_25896 = io_op_bits_active_vstx ? _GEN_25088 : _GEN_23558; // @[sequencer-master.scala 652:39]
  wire  _GEN_25897 = io_op_bits_active_vstx ? _GEN_25089 : _GEN_23559; // @[sequencer-master.scala 652:39]
  wire  _GEN_25898 = io_op_bits_active_vstx ? _GEN_25090 : _GEN_23560; // @[sequencer-master.scala 652:39]
  wire  _GEN_25899 = io_op_bits_active_vstx ? _GEN_25091 : _GEN_23561; // @[sequencer-master.scala 652:39]
  wire  _GEN_25900 = io_op_bits_active_vstx ? _GEN_25092 : _GEN_23562; // @[sequencer-master.scala 652:39]
  wire  _GEN_25901 = io_op_bits_active_vstx ? _GEN_25093 : _GEN_23563; // @[sequencer-master.scala 652:39]
  wire  _GEN_25902 = io_op_bits_active_vstx ? _GEN_25094 : _GEN_23564; // @[sequencer-master.scala 652:39]
  wire  _GEN_25903 = io_op_bits_active_vstx ? _GEN_25095 : _GEN_23565; // @[sequencer-master.scala 652:39]
  wire  _GEN_25904 = io_op_bits_active_vstx ? _GEN_25096 : _GEN_23566; // @[sequencer-master.scala 652:39]
  wire  _GEN_25905 = io_op_bits_active_vstx ? _GEN_25097 : _GEN_23567; // @[sequencer-master.scala 652:39]
  wire  _GEN_25906 = io_op_bits_active_vstx ? _GEN_25098 : _GEN_23568; // @[sequencer-master.scala 652:39]
  wire  _GEN_25907 = io_op_bits_active_vstx ? _GEN_25099 : _GEN_23569; // @[sequencer-master.scala 652:39]
  wire  _GEN_25908 = io_op_bits_active_vstx ? _GEN_25100 : _GEN_23570; // @[sequencer-master.scala 652:39]
  wire  _GEN_25909 = io_op_bits_active_vstx ? _GEN_25101 : _GEN_23571; // @[sequencer-master.scala 652:39]
  wire  _GEN_25910 = io_op_bits_active_vstx ? _GEN_25102 : _GEN_23572; // @[sequencer-master.scala 652:39]
  wire  _GEN_25911 = io_op_bits_active_vstx ? _GEN_25103 : _GEN_23573; // @[sequencer-master.scala 652:39]
  wire  _GEN_25912 = io_op_bits_active_vstx ? _GEN_25104 : _GEN_23574; // @[sequencer-master.scala 652:39]
  wire  _GEN_25913 = io_op_bits_active_vstx ? _GEN_25105 : _GEN_23575; // @[sequencer-master.scala 652:39]
  wire  _GEN_25914 = io_op_bits_active_vstx ? _GEN_25106 : _GEN_23576; // @[sequencer-master.scala 652:39]
  wire  _GEN_25915 = io_op_bits_active_vstx ? _GEN_25107 : _GEN_23577; // @[sequencer-master.scala 652:39]
  wire  _GEN_25916 = io_op_bits_active_vstx ? _GEN_25108 : _GEN_23578; // @[sequencer-master.scala 652:39]
  wire  _GEN_25917 = io_op_bits_active_vstx ? _GEN_25109 : _GEN_23579; // @[sequencer-master.scala 652:39]
  wire  _GEN_25918 = io_op_bits_active_vstx ? _GEN_25110 : _GEN_23580; // @[sequencer-master.scala 652:39]
  wire  _GEN_25919 = io_op_bits_active_vstx ? _GEN_25111 : _GEN_23581; // @[sequencer-master.scala 652:39]
  wire  _GEN_25920 = io_op_bits_active_vstx ? _GEN_25792 : _GEN_23582; // @[sequencer-master.scala 652:39]
  wire  _GEN_25921 = io_op_bits_active_vstx ? _GEN_25800 : _GEN_23583; // @[sequencer-master.scala 652:39]
  wire  _GEN_25922 = io_op_bits_active_vstx ? _GEN_25808 : _GEN_23584; // @[sequencer-master.scala 652:39]
  wire  _GEN_25923 = io_op_bits_active_vstx ? _GEN_25816 : _GEN_23585; // @[sequencer-master.scala 652:39]
  wire  _GEN_25924 = io_op_bits_active_vstx ? _GEN_25824 : _GEN_23586; // @[sequencer-master.scala 652:39]
  wire  _GEN_25925 = io_op_bits_active_vstx ? _GEN_25832 : _GEN_23587; // @[sequencer-master.scala 652:39]
  wire  _GEN_25926 = io_op_bits_active_vstx ? _GEN_25840 : _GEN_23588; // @[sequencer-master.scala 652:39]
  wire  _GEN_25927 = io_op_bits_active_vstx ? _GEN_25848 : _GEN_23589; // @[sequencer-master.scala 652:39]
  wire  _GEN_25928 = io_op_bits_active_vstx ? _GEN_25120 : _GEN_23590; // @[sequencer-master.scala 652:39]
  wire  _GEN_25929 = io_op_bits_active_vstx ? _GEN_25121 : _GEN_23591; // @[sequencer-master.scala 652:39]
  wire  _GEN_25930 = io_op_bits_active_vstx ? _GEN_25122 : _GEN_23592; // @[sequencer-master.scala 652:39]
  wire  _GEN_25931 = io_op_bits_active_vstx ? _GEN_25123 : _GEN_23593; // @[sequencer-master.scala 652:39]
  wire  _GEN_25932 = io_op_bits_active_vstx ? _GEN_25124 : _GEN_23594; // @[sequencer-master.scala 652:39]
  wire  _GEN_25933 = io_op_bits_active_vstx ? _GEN_25125 : _GEN_23595; // @[sequencer-master.scala 652:39]
  wire  _GEN_25934 = io_op_bits_active_vstx ? _GEN_25126 : _GEN_23596; // @[sequencer-master.scala 652:39]
  wire  _GEN_25935 = io_op_bits_active_vstx ? _GEN_25127 : _GEN_23597; // @[sequencer-master.scala 652:39]
  wire  _GEN_25936 = io_op_bits_active_vstx ? _GEN_25128 : _GEN_23598; // @[sequencer-master.scala 652:39]
  wire  _GEN_25937 = io_op_bits_active_vstx ? _GEN_25129 : _GEN_23599; // @[sequencer-master.scala 652:39]
  wire  _GEN_25938 = io_op_bits_active_vstx ? _GEN_25130 : _GEN_23600; // @[sequencer-master.scala 652:39]
  wire  _GEN_25939 = io_op_bits_active_vstx ? _GEN_25131 : _GEN_23601; // @[sequencer-master.scala 652:39]
  wire  _GEN_25940 = io_op_bits_active_vstx ? _GEN_25132 : _GEN_23602; // @[sequencer-master.scala 652:39]
  wire  _GEN_25941 = io_op_bits_active_vstx ? _GEN_25133 : _GEN_23603; // @[sequencer-master.scala 652:39]
  wire  _GEN_25942 = io_op_bits_active_vstx ? _GEN_25134 : _GEN_23604; // @[sequencer-master.scala 652:39]
  wire  _GEN_25943 = io_op_bits_active_vstx ? _GEN_25135 : _GEN_23605; // @[sequencer-master.scala 652:39]
  wire  _GEN_25944 = io_op_bits_active_vstx ? _GEN_25793 : _GEN_23606; // @[sequencer-master.scala 652:39]
  wire  _GEN_25945 = io_op_bits_active_vstx ? _GEN_25801 : _GEN_23607; // @[sequencer-master.scala 652:39]
  wire  _GEN_25946 = io_op_bits_active_vstx ? _GEN_25809 : _GEN_23608; // @[sequencer-master.scala 652:39]
  wire  _GEN_25947 = io_op_bits_active_vstx ? _GEN_25817 : _GEN_23609; // @[sequencer-master.scala 652:39]
  wire  _GEN_25948 = io_op_bits_active_vstx ? _GEN_25825 : _GEN_23610; // @[sequencer-master.scala 652:39]
  wire  _GEN_25949 = io_op_bits_active_vstx ? _GEN_25833 : _GEN_23611; // @[sequencer-master.scala 652:39]
  wire  _GEN_25950 = io_op_bits_active_vstx ? _GEN_25841 : _GEN_23612; // @[sequencer-master.scala 652:39]
  wire  _GEN_25951 = io_op_bits_active_vstx ? _GEN_25849 : _GEN_23613; // @[sequencer-master.scala 652:39]
  wire  _GEN_25952 = io_op_bits_active_vstx ? _GEN_25144 : _GEN_23614; // @[sequencer-master.scala 652:39]
  wire  _GEN_25953 = io_op_bits_active_vstx ? _GEN_25145 : _GEN_23615; // @[sequencer-master.scala 652:39]
  wire  _GEN_25954 = io_op_bits_active_vstx ? _GEN_25146 : _GEN_23616; // @[sequencer-master.scala 652:39]
  wire  _GEN_25955 = io_op_bits_active_vstx ? _GEN_25147 : _GEN_23617; // @[sequencer-master.scala 652:39]
  wire  _GEN_25956 = io_op_bits_active_vstx ? _GEN_25148 : _GEN_23618; // @[sequencer-master.scala 652:39]
  wire  _GEN_25957 = io_op_bits_active_vstx ? _GEN_25149 : _GEN_23619; // @[sequencer-master.scala 652:39]
  wire  _GEN_25958 = io_op_bits_active_vstx ? _GEN_25150 : _GEN_23620; // @[sequencer-master.scala 652:39]
  wire  _GEN_25959 = io_op_bits_active_vstx ? _GEN_25151 : _GEN_23621; // @[sequencer-master.scala 652:39]
  wire  _GEN_25960 = io_op_bits_active_vstx ? _GEN_25152 : _GEN_23622; // @[sequencer-master.scala 652:39]
  wire  _GEN_25961 = io_op_bits_active_vstx ? _GEN_25153 : _GEN_23623; // @[sequencer-master.scala 652:39]
  wire  _GEN_25962 = io_op_bits_active_vstx ? _GEN_25154 : _GEN_23624; // @[sequencer-master.scala 652:39]
  wire  _GEN_25963 = io_op_bits_active_vstx ? _GEN_25155 : _GEN_23625; // @[sequencer-master.scala 652:39]
  wire  _GEN_25964 = io_op_bits_active_vstx ? _GEN_25156 : _GEN_23626; // @[sequencer-master.scala 652:39]
  wire  _GEN_25965 = io_op_bits_active_vstx ? _GEN_25157 : _GEN_23627; // @[sequencer-master.scala 652:39]
  wire  _GEN_25966 = io_op_bits_active_vstx ? _GEN_25158 : _GEN_23628; // @[sequencer-master.scala 652:39]
  wire  _GEN_25967 = io_op_bits_active_vstx ? _GEN_25159 : _GEN_23629; // @[sequencer-master.scala 652:39]
  wire  _GEN_25968 = io_op_bits_active_vstx ? _GEN_25794 : _GEN_23630; // @[sequencer-master.scala 652:39]
  wire  _GEN_25969 = io_op_bits_active_vstx ? _GEN_25802 : _GEN_23631; // @[sequencer-master.scala 652:39]
  wire  _GEN_25970 = io_op_bits_active_vstx ? _GEN_25810 : _GEN_23632; // @[sequencer-master.scala 652:39]
  wire  _GEN_25971 = io_op_bits_active_vstx ? _GEN_25818 : _GEN_23633; // @[sequencer-master.scala 652:39]
  wire  _GEN_25972 = io_op_bits_active_vstx ? _GEN_25826 : _GEN_23634; // @[sequencer-master.scala 652:39]
  wire  _GEN_25973 = io_op_bits_active_vstx ? _GEN_25834 : _GEN_23635; // @[sequencer-master.scala 652:39]
  wire  _GEN_25974 = io_op_bits_active_vstx ? _GEN_25842 : _GEN_23636; // @[sequencer-master.scala 652:39]
  wire  _GEN_25975 = io_op_bits_active_vstx ? _GEN_25850 : _GEN_23637; // @[sequencer-master.scala 652:39]
  wire  _GEN_25976 = io_op_bits_active_vstx ? _GEN_25168 : _GEN_23638; // @[sequencer-master.scala 652:39]
  wire  _GEN_25977 = io_op_bits_active_vstx ? _GEN_25169 : _GEN_23639; // @[sequencer-master.scala 652:39]
  wire  _GEN_25978 = io_op_bits_active_vstx ? _GEN_25170 : _GEN_23640; // @[sequencer-master.scala 652:39]
  wire  _GEN_25979 = io_op_bits_active_vstx ? _GEN_25171 : _GEN_23641; // @[sequencer-master.scala 652:39]
  wire  _GEN_25980 = io_op_bits_active_vstx ? _GEN_25172 : _GEN_23642; // @[sequencer-master.scala 652:39]
  wire  _GEN_25981 = io_op_bits_active_vstx ? _GEN_25173 : _GEN_23643; // @[sequencer-master.scala 652:39]
  wire  _GEN_25982 = io_op_bits_active_vstx ? _GEN_25174 : _GEN_23644; // @[sequencer-master.scala 652:39]
  wire  _GEN_25983 = io_op_bits_active_vstx ? _GEN_25175 : _GEN_23645; // @[sequencer-master.scala 652:39]
  wire  _GEN_25984 = io_op_bits_active_vstx ? _GEN_25176 : _GEN_23646; // @[sequencer-master.scala 652:39]
  wire  _GEN_25985 = io_op_bits_active_vstx ? _GEN_25177 : _GEN_23647; // @[sequencer-master.scala 652:39]
  wire  _GEN_25986 = io_op_bits_active_vstx ? _GEN_25178 : _GEN_23648; // @[sequencer-master.scala 652:39]
  wire  _GEN_25987 = io_op_bits_active_vstx ? _GEN_25179 : _GEN_23649; // @[sequencer-master.scala 652:39]
  wire  _GEN_25988 = io_op_bits_active_vstx ? _GEN_25180 : _GEN_23650; // @[sequencer-master.scala 652:39]
  wire  _GEN_25989 = io_op_bits_active_vstx ? _GEN_25181 : _GEN_23651; // @[sequencer-master.scala 652:39]
  wire  _GEN_25990 = io_op_bits_active_vstx ? _GEN_25182 : _GEN_23652; // @[sequencer-master.scala 652:39]
  wire  _GEN_25991 = io_op_bits_active_vstx ? _GEN_25183 : _GEN_23653; // @[sequencer-master.scala 652:39]
  wire  _GEN_25992 = io_op_bits_active_vstx ? _GEN_25795 : _GEN_23654; // @[sequencer-master.scala 652:39]
  wire  _GEN_25993 = io_op_bits_active_vstx ? _GEN_25803 : _GEN_23655; // @[sequencer-master.scala 652:39]
  wire  _GEN_25994 = io_op_bits_active_vstx ? _GEN_25811 : _GEN_23656; // @[sequencer-master.scala 652:39]
  wire  _GEN_25995 = io_op_bits_active_vstx ? _GEN_25819 : _GEN_23657; // @[sequencer-master.scala 652:39]
  wire  _GEN_25996 = io_op_bits_active_vstx ? _GEN_25827 : _GEN_23658; // @[sequencer-master.scala 652:39]
  wire  _GEN_25997 = io_op_bits_active_vstx ? _GEN_25835 : _GEN_23659; // @[sequencer-master.scala 652:39]
  wire  _GEN_25998 = io_op_bits_active_vstx ? _GEN_25843 : _GEN_23660; // @[sequencer-master.scala 652:39]
  wire  _GEN_25999 = io_op_bits_active_vstx ? _GEN_25851 : _GEN_23661; // @[sequencer-master.scala 652:39]
  wire  _GEN_26000 = io_op_bits_active_vstx ? _GEN_25192 : _GEN_23662; // @[sequencer-master.scala 652:39]
  wire  _GEN_26001 = io_op_bits_active_vstx ? _GEN_25193 : _GEN_23663; // @[sequencer-master.scala 652:39]
  wire  _GEN_26002 = io_op_bits_active_vstx ? _GEN_25194 : _GEN_23664; // @[sequencer-master.scala 652:39]
  wire  _GEN_26003 = io_op_bits_active_vstx ? _GEN_25195 : _GEN_23665; // @[sequencer-master.scala 652:39]
  wire  _GEN_26004 = io_op_bits_active_vstx ? _GEN_25196 : _GEN_23666; // @[sequencer-master.scala 652:39]
  wire  _GEN_26005 = io_op_bits_active_vstx ? _GEN_25197 : _GEN_23667; // @[sequencer-master.scala 652:39]
  wire  _GEN_26006 = io_op_bits_active_vstx ? _GEN_25198 : _GEN_23668; // @[sequencer-master.scala 652:39]
  wire  _GEN_26007 = io_op_bits_active_vstx ? _GEN_25199 : _GEN_23669; // @[sequencer-master.scala 652:39]
  wire  _GEN_26008 = io_op_bits_active_vstx ? _GEN_25200 : _GEN_23670; // @[sequencer-master.scala 652:39]
  wire  _GEN_26009 = io_op_bits_active_vstx ? _GEN_25201 : _GEN_23671; // @[sequencer-master.scala 652:39]
  wire  _GEN_26010 = io_op_bits_active_vstx ? _GEN_25202 : _GEN_23672; // @[sequencer-master.scala 652:39]
  wire  _GEN_26011 = io_op_bits_active_vstx ? _GEN_25203 : _GEN_23673; // @[sequencer-master.scala 652:39]
  wire  _GEN_26012 = io_op_bits_active_vstx ? _GEN_25204 : _GEN_23674; // @[sequencer-master.scala 652:39]
  wire  _GEN_26013 = io_op_bits_active_vstx ? _GEN_25205 : _GEN_23675; // @[sequencer-master.scala 652:39]
  wire  _GEN_26014 = io_op_bits_active_vstx ? _GEN_25206 : _GEN_23676; // @[sequencer-master.scala 652:39]
  wire  _GEN_26015 = io_op_bits_active_vstx ? _GEN_25207 : _GEN_23677; // @[sequencer-master.scala 652:39]
  wire  _GEN_26016 = io_op_bits_active_vstx ? _GEN_25796 : _GEN_23678; // @[sequencer-master.scala 652:39]
  wire  _GEN_26017 = io_op_bits_active_vstx ? _GEN_25804 : _GEN_23679; // @[sequencer-master.scala 652:39]
  wire  _GEN_26018 = io_op_bits_active_vstx ? _GEN_25812 : _GEN_23680; // @[sequencer-master.scala 652:39]
  wire  _GEN_26019 = io_op_bits_active_vstx ? _GEN_25820 : _GEN_23681; // @[sequencer-master.scala 652:39]
  wire  _GEN_26020 = io_op_bits_active_vstx ? _GEN_25828 : _GEN_23682; // @[sequencer-master.scala 652:39]
  wire  _GEN_26021 = io_op_bits_active_vstx ? _GEN_25836 : _GEN_23683; // @[sequencer-master.scala 652:39]
  wire  _GEN_26022 = io_op_bits_active_vstx ? _GEN_25844 : _GEN_23684; // @[sequencer-master.scala 652:39]
  wire  _GEN_26023 = io_op_bits_active_vstx ? _GEN_25852 : _GEN_23685; // @[sequencer-master.scala 652:39]
  wire  _GEN_26024 = io_op_bits_active_vstx ? _GEN_25216 : _GEN_23686; // @[sequencer-master.scala 652:39]
  wire  _GEN_26025 = io_op_bits_active_vstx ? _GEN_25217 : _GEN_23687; // @[sequencer-master.scala 652:39]
  wire  _GEN_26026 = io_op_bits_active_vstx ? _GEN_25218 : _GEN_23688; // @[sequencer-master.scala 652:39]
  wire  _GEN_26027 = io_op_bits_active_vstx ? _GEN_25219 : _GEN_23689; // @[sequencer-master.scala 652:39]
  wire  _GEN_26028 = io_op_bits_active_vstx ? _GEN_25220 : _GEN_23690; // @[sequencer-master.scala 652:39]
  wire  _GEN_26029 = io_op_bits_active_vstx ? _GEN_25221 : _GEN_23691; // @[sequencer-master.scala 652:39]
  wire  _GEN_26030 = io_op_bits_active_vstx ? _GEN_25222 : _GEN_23692; // @[sequencer-master.scala 652:39]
  wire  _GEN_26031 = io_op_bits_active_vstx ? _GEN_25223 : _GEN_23693; // @[sequencer-master.scala 652:39]
  wire  _GEN_26032 = io_op_bits_active_vstx ? _GEN_25224 : _GEN_23694; // @[sequencer-master.scala 652:39]
  wire  _GEN_26033 = io_op_bits_active_vstx ? _GEN_25225 : _GEN_23695; // @[sequencer-master.scala 652:39]
  wire  _GEN_26034 = io_op_bits_active_vstx ? _GEN_25226 : _GEN_23696; // @[sequencer-master.scala 652:39]
  wire  _GEN_26035 = io_op_bits_active_vstx ? _GEN_25227 : _GEN_23697; // @[sequencer-master.scala 652:39]
  wire  _GEN_26036 = io_op_bits_active_vstx ? _GEN_25228 : _GEN_23698; // @[sequencer-master.scala 652:39]
  wire  _GEN_26037 = io_op_bits_active_vstx ? _GEN_25229 : _GEN_23699; // @[sequencer-master.scala 652:39]
  wire  _GEN_26038 = io_op_bits_active_vstx ? _GEN_25230 : _GEN_23700; // @[sequencer-master.scala 652:39]
  wire  _GEN_26039 = io_op_bits_active_vstx ? _GEN_25231 : _GEN_23701; // @[sequencer-master.scala 652:39]
  wire  _GEN_26040 = io_op_bits_active_vstx ? _GEN_25797 : _GEN_23702; // @[sequencer-master.scala 652:39]
  wire  _GEN_26041 = io_op_bits_active_vstx ? _GEN_25805 : _GEN_23703; // @[sequencer-master.scala 652:39]
  wire  _GEN_26042 = io_op_bits_active_vstx ? _GEN_25813 : _GEN_23704; // @[sequencer-master.scala 652:39]
  wire  _GEN_26043 = io_op_bits_active_vstx ? _GEN_25821 : _GEN_23705; // @[sequencer-master.scala 652:39]
  wire  _GEN_26044 = io_op_bits_active_vstx ? _GEN_25829 : _GEN_23706; // @[sequencer-master.scala 652:39]
  wire  _GEN_26045 = io_op_bits_active_vstx ? _GEN_25837 : _GEN_23707; // @[sequencer-master.scala 652:39]
  wire  _GEN_26046 = io_op_bits_active_vstx ? _GEN_25845 : _GEN_23708; // @[sequencer-master.scala 652:39]
  wire  _GEN_26047 = io_op_bits_active_vstx ? _GEN_25853 : _GEN_23709; // @[sequencer-master.scala 652:39]
  wire  _GEN_26048 = io_op_bits_active_vstx ? _GEN_25240 : _GEN_23710; // @[sequencer-master.scala 652:39]
  wire  _GEN_26049 = io_op_bits_active_vstx ? _GEN_25241 : _GEN_23711; // @[sequencer-master.scala 652:39]
  wire  _GEN_26050 = io_op_bits_active_vstx ? _GEN_25242 : _GEN_23712; // @[sequencer-master.scala 652:39]
  wire  _GEN_26051 = io_op_bits_active_vstx ? _GEN_25243 : _GEN_23713; // @[sequencer-master.scala 652:39]
  wire  _GEN_26052 = io_op_bits_active_vstx ? _GEN_25244 : _GEN_23714; // @[sequencer-master.scala 652:39]
  wire  _GEN_26053 = io_op_bits_active_vstx ? _GEN_25245 : _GEN_23715; // @[sequencer-master.scala 652:39]
  wire  _GEN_26054 = io_op_bits_active_vstx ? _GEN_25246 : _GEN_23716; // @[sequencer-master.scala 652:39]
  wire  _GEN_26055 = io_op_bits_active_vstx ? _GEN_25247 : _GEN_23717; // @[sequencer-master.scala 652:39]
  wire  _GEN_26056 = io_op_bits_active_vstx ? _GEN_25248 : _GEN_23718; // @[sequencer-master.scala 652:39]
  wire  _GEN_26057 = io_op_bits_active_vstx ? _GEN_25249 : _GEN_23719; // @[sequencer-master.scala 652:39]
  wire  _GEN_26058 = io_op_bits_active_vstx ? _GEN_25250 : _GEN_23720; // @[sequencer-master.scala 652:39]
  wire  _GEN_26059 = io_op_bits_active_vstx ? _GEN_25251 : _GEN_23721; // @[sequencer-master.scala 652:39]
  wire  _GEN_26060 = io_op_bits_active_vstx ? _GEN_25252 : _GEN_23722; // @[sequencer-master.scala 652:39]
  wire  _GEN_26061 = io_op_bits_active_vstx ? _GEN_25253 : _GEN_23723; // @[sequencer-master.scala 652:39]
  wire  _GEN_26062 = io_op_bits_active_vstx ? _GEN_25254 : _GEN_23724; // @[sequencer-master.scala 652:39]
  wire  _GEN_26063 = io_op_bits_active_vstx ? _GEN_25255 : _GEN_23725; // @[sequencer-master.scala 652:39]
  wire  _GEN_26064 = io_op_bits_active_vstx ? _GEN_25798 : _GEN_23726; // @[sequencer-master.scala 652:39]
  wire  _GEN_26065 = io_op_bits_active_vstx ? _GEN_25806 : _GEN_23727; // @[sequencer-master.scala 652:39]
  wire  _GEN_26066 = io_op_bits_active_vstx ? _GEN_25814 : _GEN_23728; // @[sequencer-master.scala 652:39]
  wire  _GEN_26067 = io_op_bits_active_vstx ? _GEN_25822 : _GEN_23729; // @[sequencer-master.scala 652:39]
  wire  _GEN_26068 = io_op_bits_active_vstx ? _GEN_25830 : _GEN_23730; // @[sequencer-master.scala 652:39]
  wire  _GEN_26069 = io_op_bits_active_vstx ? _GEN_25838 : _GEN_23731; // @[sequencer-master.scala 652:39]
  wire  _GEN_26070 = io_op_bits_active_vstx ? _GEN_25846 : _GEN_23732; // @[sequencer-master.scala 652:39]
  wire  _GEN_26071 = io_op_bits_active_vstx ? _GEN_25854 : _GEN_23733; // @[sequencer-master.scala 652:39]
  wire  _GEN_26072 = io_op_bits_active_vstx ? _GEN_25264 : _GEN_23734; // @[sequencer-master.scala 652:39]
  wire  _GEN_26073 = io_op_bits_active_vstx ? _GEN_25265 : _GEN_23735; // @[sequencer-master.scala 652:39]
  wire  _GEN_26074 = io_op_bits_active_vstx ? _GEN_25266 : _GEN_23736; // @[sequencer-master.scala 652:39]
  wire  _GEN_26075 = io_op_bits_active_vstx ? _GEN_25267 : _GEN_23737; // @[sequencer-master.scala 652:39]
  wire  _GEN_26076 = io_op_bits_active_vstx ? _GEN_25268 : _GEN_23738; // @[sequencer-master.scala 652:39]
  wire  _GEN_26077 = io_op_bits_active_vstx ? _GEN_25269 : _GEN_23739; // @[sequencer-master.scala 652:39]
  wire  _GEN_26078 = io_op_bits_active_vstx ? _GEN_25270 : _GEN_23740; // @[sequencer-master.scala 652:39]
  wire  _GEN_26079 = io_op_bits_active_vstx ? _GEN_25271 : _GEN_23741; // @[sequencer-master.scala 652:39]
  wire  _GEN_26080 = io_op_bits_active_vstx ? _GEN_25272 : _GEN_23742; // @[sequencer-master.scala 652:39]
  wire  _GEN_26081 = io_op_bits_active_vstx ? _GEN_25273 : _GEN_23743; // @[sequencer-master.scala 652:39]
  wire  _GEN_26082 = io_op_bits_active_vstx ? _GEN_25274 : _GEN_23744; // @[sequencer-master.scala 652:39]
  wire  _GEN_26083 = io_op_bits_active_vstx ? _GEN_25275 : _GEN_23745; // @[sequencer-master.scala 652:39]
  wire  _GEN_26084 = io_op_bits_active_vstx ? _GEN_25276 : _GEN_23746; // @[sequencer-master.scala 652:39]
  wire  _GEN_26085 = io_op_bits_active_vstx ? _GEN_25277 : _GEN_23747; // @[sequencer-master.scala 652:39]
  wire  _GEN_26086 = io_op_bits_active_vstx ? _GEN_25278 : _GEN_23748; // @[sequencer-master.scala 652:39]
  wire  _GEN_26087 = io_op_bits_active_vstx ? _GEN_25279 : _GEN_23749; // @[sequencer-master.scala 652:39]
  wire  _GEN_26088 = io_op_bits_active_vstx ? _GEN_25799 : _GEN_23750; // @[sequencer-master.scala 652:39]
  wire  _GEN_26089 = io_op_bits_active_vstx ? _GEN_25807 : _GEN_23751; // @[sequencer-master.scala 652:39]
  wire  _GEN_26090 = io_op_bits_active_vstx ? _GEN_25815 : _GEN_23752; // @[sequencer-master.scala 652:39]
  wire  _GEN_26091 = io_op_bits_active_vstx ? _GEN_25823 : _GEN_23753; // @[sequencer-master.scala 652:39]
  wire  _GEN_26092 = io_op_bits_active_vstx ? _GEN_25831 : _GEN_23754; // @[sequencer-master.scala 652:39]
  wire  _GEN_26093 = io_op_bits_active_vstx ? _GEN_25839 : _GEN_23755; // @[sequencer-master.scala 652:39]
  wire  _GEN_26094 = io_op_bits_active_vstx ? _GEN_25847 : _GEN_23756; // @[sequencer-master.scala 652:39]
  wire  _GEN_26095 = io_op_bits_active_vstx ? _GEN_25855 : _GEN_23757; // @[sequencer-master.scala 652:39]
  wire  _GEN_26096 = io_op_bits_active_vstx ? _GEN_25288 : _GEN_23758; // @[sequencer-master.scala 652:39]
  wire  _GEN_26097 = io_op_bits_active_vstx ? _GEN_25289 : _GEN_23759; // @[sequencer-master.scala 652:39]
  wire  _GEN_26098 = io_op_bits_active_vstx ? _GEN_25290 : _GEN_23760; // @[sequencer-master.scala 652:39]
  wire  _GEN_26099 = io_op_bits_active_vstx ? _GEN_25291 : _GEN_23761; // @[sequencer-master.scala 652:39]
  wire  _GEN_26100 = io_op_bits_active_vstx ? _GEN_25292 : _GEN_23762; // @[sequencer-master.scala 652:39]
  wire  _GEN_26101 = io_op_bits_active_vstx ? _GEN_25293 : _GEN_23763; // @[sequencer-master.scala 652:39]
  wire  _GEN_26102 = io_op_bits_active_vstx ? _GEN_25294 : _GEN_23764; // @[sequencer-master.scala 652:39]
  wire  _GEN_26103 = io_op_bits_active_vstx ? _GEN_25295 : _GEN_23765; // @[sequencer-master.scala 652:39]
  wire  _GEN_26104 = io_op_bits_active_vstx ? _GEN_25296 : _GEN_23766; // @[sequencer-master.scala 652:39]
  wire  _GEN_26105 = io_op_bits_active_vstx ? _GEN_25297 : _GEN_23767; // @[sequencer-master.scala 652:39]
  wire  _GEN_26106 = io_op_bits_active_vstx ? _GEN_25298 : _GEN_23768; // @[sequencer-master.scala 652:39]
  wire  _GEN_26107 = io_op_bits_active_vstx ? _GEN_25299 : _GEN_23769; // @[sequencer-master.scala 652:39]
  wire  _GEN_26108 = io_op_bits_active_vstx ? _GEN_25300 : _GEN_23770; // @[sequencer-master.scala 652:39]
  wire  _GEN_26109 = io_op_bits_active_vstx ? _GEN_25301 : _GEN_23771; // @[sequencer-master.scala 652:39]
  wire  _GEN_26110 = io_op_bits_active_vstx ? _GEN_25302 : _GEN_23772; // @[sequencer-master.scala 652:39]
  wire  _GEN_26111 = io_op_bits_active_vstx ? _GEN_25303 : _GEN_23773; // @[sequencer-master.scala 652:39]
  wire  _GEN_26112 = io_op_bits_active_vstx ? _GEN_25304 : _GEN_23774; // @[sequencer-master.scala 652:39]
  wire  _GEN_26113 = io_op_bits_active_vstx ? _GEN_25305 : _GEN_23775; // @[sequencer-master.scala 652:39]
  wire  _GEN_26114 = io_op_bits_active_vstx ? _GEN_25306 : _GEN_23776; // @[sequencer-master.scala 652:39]
  wire  _GEN_26115 = io_op_bits_active_vstx ? _GEN_25307 : _GEN_23777; // @[sequencer-master.scala 652:39]
  wire  _GEN_26116 = io_op_bits_active_vstx ? _GEN_25308 : _GEN_23778; // @[sequencer-master.scala 652:39]
  wire  _GEN_26117 = io_op_bits_active_vstx ? _GEN_25309 : _GEN_23779; // @[sequencer-master.scala 652:39]
  wire  _GEN_26118 = io_op_bits_active_vstx ? _GEN_25310 : _GEN_23780; // @[sequencer-master.scala 652:39]
  wire  _GEN_26119 = io_op_bits_active_vstx ? _GEN_25311 : _GEN_23781; // @[sequencer-master.scala 652:39]
  wire  _GEN_26128 = io_op_bits_active_vstx ? _GEN_24240 : _GEN_23790; // @[sequencer-master.scala 652:39]
  wire  _GEN_26129 = io_op_bits_active_vstx ? _GEN_24241 : _GEN_23791; // @[sequencer-master.scala 652:39]
  wire  _GEN_26130 = io_op_bits_active_vstx ? _GEN_24242 : _GEN_23792; // @[sequencer-master.scala 652:39]
  wire  _GEN_26131 = io_op_bits_active_vstx ? _GEN_24243 : _GEN_23793; // @[sequencer-master.scala 652:39]
  wire  _GEN_26132 = io_op_bits_active_vstx ? _GEN_24244 : _GEN_23794; // @[sequencer-master.scala 652:39]
  wire  _GEN_26133 = io_op_bits_active_vstx ? _GEN_24245 : _GEN_23795; // @[sequencer-master.scala 652:39]
  wire  _GEN_26134 = io_op_bits_active_vstx ? _GEN_24246 : _GEN_23796; // @[sequencer-master.scala 652:39]
  wire  _GEN_26135 = io_op_bits_active_vstx ? _GEN_24247 : _GEN_23797; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26136 = io_op_bits_active_vstx ? _GEN_25328 : _GEN_23798; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26137 = io_op_bits_active_vstx ? _GEN_25329 : _GEN_23799; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26138 = io_op_bits_active_vstx ? _GEN_25330 : _GEN_23800; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26139 = io_op_bits_active_vstx ? _GEN_25331 : _GEN_23801; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26140 = io_op_bits_active_vstx ? _GEN_25332 : _GEN_23802; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26141 = io_op_bits_active_vstx ? _GEN_25333 : _GEN_23803; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26142 = io_op_bits_active_vstx ? _GEN_25334 : _GEN_23804; // @[sequencer-master.scala 652:39]
  wire [9:0] _GEN_26143 = io_op_bits_active_vstx ? _GEN_25335 : _GEN_23805; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26144 = io_op_bits_active_vstx ? _GEN_25376 : _GEN_23806; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26145 = io_op_bits_active_vstx ? _GEN_25377 : _GEN_23807; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26146 = io_op_bits_active_vstx ? _GEN_25378 : _GEN_23808; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26147 = io_op_bits_active_vstx ? _GEN_25379 : _GEN_23809; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26148 = io_op_bits_active_vstx ? _GEN_25380 : _GEN_23810; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26149 = io_op_bits_active_vstx ? _GEN_25381 : _GEN_23811; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26150 = io_op_bits_active_vstx ? _GEN_25382 : _GEN_23812; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26151 = io_op_bits_active_vstx ? _GEN_25383 : _GEN_23813; // @[sequencer-master.scala 652:39]
  wire  _GEN_26152 = io_op_bits_active_vstx ? _GEN_25392 : _GEN_23814; // @[sequencer-master.scala 652:39]
  wire  _GEN_26153 = io_op_bits_active_vstx ? _GEN_25393 : _GEN_23815; // @[sequencer-master.scala 652:39]
  wire  _GEN_26154 = io_op_bits_active_vstx ? _GEN_25394 : _GEN_23816; // @[sequencer-master.scala 652:39]
  wire  _GEN_26155 = io_op_bits_active_vstx ? _GEN_25395 : _GEN_23817; // @[sequencer-master.scala 652:39]
  wire  _GEN_26156 = io_op_bits_active_vstx ? _GEN_25396 : _GEN_23818; // @[sequencer-master.scala 652:39]
  wire  _GEN_26157 = io_op_bits_active_vstx ? _GEN_25397 : _GEN_23819; // @[sequencer-master.scala 652:39]
  wire  _GEN_26158 = io_op_bits_active_vstx ? _GEN_25398 : _GEN_23820; // @[sequencer-master.scala 652:39]
  wire  _GEN_26159 = io_op_bits_active_vstx ? _GEN_25399 : _GEN_23821; // @[sequencer-master.scala 652:39]
  wire  _GEN_26160 = io_op_bits_active_vstx ? _GEN_25400 : _GEN_23822; // @[sequencer-master.scala 652:39]
  wire  _GEN_26161 = io_op_bits_active_vstx ? _GEN_25401 : _GEN_23823; // @[sequencer-master.scala 652:39]
  wire  _GEN_26162 = io_op_bits_active_vstx ? _GEN_25402 : _GEN_23824; // @[sequencer-master.scala 652:39]
  wire  _GEN_26163 = io_op_bits_active_vstx ? _GEN_25403 : _GEN_23825; // @[sequencer-master.scala 652:39]
  wire  _GEN_26164 = io_op_bits_active_vstx ? _GEN_25404 : _GEN_23826; // @[sequencer-master.scala 652:39]
  wire  _GEN_26165 = io_op_bits_active_vstx ? _GEN_25405 : _GEN_23827; // @[sequencer-master.scala 652:39]
  wire  _GEN_26166 = io_op_bits_active_vstx ? _GEN_25406 : _GEN_23828; // @[sequencer-master.scala 652:39]
  wire  _GEN_26167 = io_op_bits_active_vstx ? _GEN_25407 : _GEN_23829; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26168 = io_op_bits_active_vstx ? _GEN_25408 : _GEN_23830; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26169 = io_op_bits_active_vstx ? _GEN_25409 : _GEN_23831; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26170 = io_op_bits_active_vstx ? _GEN_25410 : _GEN_23832; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26171 = io_op_bits_active_vstx ? _GEN_25411 : _GEN_23833; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26172 = io_op_bits_active_vstx ? _GEN_25412 : _GEN_23834; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26173 = io_op_bits_active_vstx ? _GEN_25413 : _GEN_23835; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26174 = io_op_bits_active_vstx ? _GEN_25414 : _GEN_23836; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26175 = io_op_bits_active_vstx ? _GEN_25415 : _GEN_23837; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26176 = io_op_bits_active_vstx ? _GEN_25592 : _GEN_23838; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26177 = io_op_bits_active_vstx ? _GEN_25593 : _GEN_23839; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26178 = io_op_bits_active_vstx ? _GEN_25594 : _GEN_23840; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26179 = io_op_bits_active_vstx ? _GEN_25595 : _GEN_23841; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26180 = io_op_bits_active_vstx ? _GEN_25596 : _GEN_23842; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26181 = io_op_bits_active_vstx ? _GEN_25597 : _GEN_23843; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26182 = io_op_bits_active_vstx ? _GEN_25598 : _GEN_23844; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26183 = io_op_bits_active_vstx ? _GEN_25599 : _GEN_23845; // @[sequencer-master.scala 652:39]
  wire  _GEN_26184 = io_op_bits_active_vstx ? _GEN_25608 : _GEN_23846; // @[sequencer-master.scala 652:39]
  wire  _GEN_26185 = io_op_bits_active_vstx ? _GEN_25609 : _GEN_23847; // @[sequencer-master.scala 652:39]
  wire  _GEN_26186 = io_op_bits_active_vstx ? _GEN_25610 : _GEN_23848; // @[sequencer-master.scala 652:39]
  wire  _GEN_26187 = io_op_bits_active_vstx ? _GEN_25611 : _GEN_23849; // @[sequencer-master.scala 652:39]
  wire  _GEN_26188 = io_op_bits_active_vstx ? _GEN_25612 : _GEN_23850; // @[sequencer-master.scala 652:39]
  wire  _GEN_26189 = io_op_bits_active_vstx ? _GEN_25613 : _GEN_23851; // @[sequencer-master.scala 652:39]
  wire  _GEN_26190 = io_op_bits_active_vstx ? _GEN_25614 : _GEN_23852; // @[sequencer-master.scala 652:39]
  wire  _GEN_26191 = io_op_bits_active_vstx ? _GEN_25615 : _GEN_23853; // @[sequencer-master.scala 652:39]
  wire  _GEN_26192 = io_op_bits_active_vstx ? _GEN_25616 : _GEN_23854; // @[sequencer-master.scala 652:39]
  wire  _GEN_26193 = io_op_bits_active_vstx ? _GEN_25617 : _GEN_23855; // @[sequencer-master.scala 652:39]
  wire  _GEN_26194 = io_op_bits_active_vstx ? _GEN_25618 : _GEN_23856; // @[sequencer-master.scala 652:39]
  wire  _GEN_26195 = io_op_bits_active_vstx ? _GEN_25619 : _GEN_23857; // @[sequencer-master.scala 652:39]
  wire  _GEN_26196 = io_op_bits_active_vstx ? _GEN_25620 : _GEN_23858; // @[sequencer-master.scala 652:39]
  wire  _GEN_26197 = io_op_bits_active_vstx ? _GEN_25621 : _GEN_23859; // @[sequencer-master.scala 652:39]
  wire  _GEN_26198 = io_op_bits_active_vstx ? _GEN_25622 : _GEN_23860; // @[sequencer-master.scala 652:39]
  wire  _GEN_26199 = io_op_bits_active_vstx ? _GEN_25623 : _GEN_23861; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26200 = io_op_bits_active_vstx ? _GEN_25624 : _GEN_23862; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26201 = io_op_bits_active_vstx ? _GEN_25625 : _GEN_23863; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26202 = io_op_bits_active_vstx ? _GEN_25626 : _GEN_23864; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26203 = io_op_bits_active_vstx ? _GEN_25627 : _GEN_23865; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26204 = io_op_bits_active_vstx ? _GEN_25628 : _GEN_23866; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26205 = io_op_bits_active_vstx ? _GEN_25629 : _GEN_23867; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26206 = io_op_bits_active_vstx ? _GEN_25630 : _GEN_23868; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26207 = io_op_bits_active_vstx ? _GEN_25631 : _GEN_23869; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26208 = io_op_bits_active_vstx ? _GEN_25632 : _GEN_23870; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26209 = io_op_bits_active_vstx ? _GEN_25633 : _GEN_23871; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26210 = io_op_bits_active_vstx ? _GEN_25634 : _GEN_23872; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26211 = io_op_bits_active_vstx ? _GEN_25635 : _GEN_23873; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26212 = io_op_bits_active_vstx ? _GEN_25636 : _GEN_23874; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26213 = io_op_bits_active_vstx ? _GEN_25637 : _GEN_23875; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26214 = io_op_bits_active_vstx ? _GEN_25638 : _GEN_23876; // @[sequencer-master.scala 652:39]
  wire [7:0] _GEN_26215 = io_op_bits_active_vstx ? _GEN_25639 : _GEN_23877; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26224 = io_op_bits_active_vstx ? _GEN_25768 : _GEN_23886; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26225 = io_op_bits_active_vstx ? _GEN_25769 : _GEN_23887; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26226 = io_op_bits_active_vstx ? _GEN_25770 : _GEN_23888; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26227 = io_op_bits_active_vstx ? _GEN_25771 : _GEN_23889; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26228 = io_op_bits_active_vstx ? _GEN_25772 : _GEN_23890; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26229 = io_op_bits_active_vstx ? _GEN_25773 : _GEN_23891; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26230 = io_op_bits_active_vstx ? _GEN_25774 : _GEN_23892; // @[sequencer-master.scala 652:39]
  wire [1:0] _GEN_26231 = io_op_bits_active_vstx ? _GEN_25775 : _GEN_23893; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26232 = io_op_bits_active_vstx ? _GEN_25776 : _GEN_23894; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26233 = io_op_bits_active_vstx ? _GEN_25777 : _GEN_23895; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26234 = io_op_bits_active_vstx ? _GEN_25778 : _GEN_23896; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26235 = io_op_bits_active_vstx ? _GEN_25779 : _GEN_23897; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26236 = io_op_bits_active_vstx ? _GEN_25780 : _GEN_23898; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26237 = io_op_bits_active_vstx ? _GEN_25781 : _GEN_23899; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26238 = io_op_bits_active_vstx ? _GEN_25782 : _GEN_23900; // @[sequencer-master.scala 652:39]
  wire [3:0] _GEN_26239 = io_op_bits_active_vstx ? _GEN_25783 : _GEN_23901; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26240 = io_op_bits_active_vstx ? _GEN_25784 : _GEN_23902; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26241 = io_op_bits_active_vstx ? _GEN_25785 : _GEN_23903; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26242 = io_op_bits_active_vstx ? _GEN_25786 : _GEN_23904; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26243 = io_op_bits_active_vstx ? _GEN_25787 : _GEN_23905; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26244 = io_op_bits_active_vstx ? _GEN_25788 : _GEN_23906; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26245 = io_op_bits_active_vstx ? _GEN_25789 : _GEN_23907; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26246 = io_op_bits_active_vstx ? _GEN_25790 : _GEN_23908; // @[sequencer-master.scala 652:39]
  wire [2:0] _GEN_26247 = io_op_bits_active_vstx ? _GEN_25791 : _GEN_23909; // @[sequencer-master.scala 652:39]
  wire  _GEN_26248 = io_op_bits_active_vstx ? _GEN_25008 : _GEN_23910; // @[sequencer-master.scala 652:39]
  wire  _GEN_26249 = io_op_bits_active_vstx ? _GEN_25009 : _GEN_23911; // @[sequencer-master.scala 652:39]
  wire  _GEN_26250 = io_op_bits_active_vstx ? _GEN_25010 : _GEN_23912; // @[sequencer-master.scala 652:39]
  wire  _GEN_26251 = io_op_bits_active_vstx ? _GEN_25011 : _GEN_23913; // @[sequencer-master.scala 652:39]
  wire  _GEN_26252 = io_op_bits_active_vstx ? _GEN_25012 : _GEN_23914; // @[sequencer-master.scala 652:39]
  wire  _GEN_26253 = io_op_bits_active_vstx ? _GEN_25013 : _GEN_23915; // @[sequencer-master.scala 652:39]
  wire  _GEN_26254 = io_op_bits_active_vstx ? _GEN_25014 : _GEN_23916; // @[sequencer-master.scala 652:39]
  wire  _GEN_26255 = io_op_bits_active_vstx ? _GEN_25015 : _GEN_23917; // @[sequencer-master.scala 652:39]
  wire  _GEN_26256 = io_op_bits_active_vstx ? _GEN_25320 : _GEN_21460; // @[sequencer-master.scala 652:39]
  wire  _GEN_26257 = io_op_bits_active_vstx ? _GEN_25321 : _GEN_21461; // @[sequencer-master.scala 652:39]
  wire  _GEN_26258 = io_op_bits_active_vstx ? _GEN_25322 : _GEN_21462; // @[sequencer-master.scala 652:39]
  wire  _GEN_26259 = io_op_bits_active_vstx ? _GEN_25323 : _GEN_21463; // @[sequencer-master.scala 652:39]
  wire  _GEN_26260 = io_op_bits_active_vstx ? _GEN_25324 : _GEN_21464; // @[sequencer-master.scala 652:39]
  wire  _GEN_26261 = io_op_bits_active_vstx ? _GEN_25325 : _GEN_21465; // @[sequencer-master.scala 652:39]
  wire  _GEN_26262 = io_op_bits_active_vstx ? _GEN_25326 : _GEN_21466; // @[sequencer-master.scala 652:39]
  wire  _GEN_26263 = io_op_bits_active_vstx ? _GEN_25327 : _GEN_21467; // @[sequencer-master.scala 652:39]
  wire  _GEN_26264 = io_op_bits_active_vstx | _GEN_23966; // @[sequencer-master.scala 652:39 sequencer-master.scala 265:41]
  wire [2:0] _GEN_26265 = io_op_bits_active_vstx ? _T_1649 : _GEN_23967; // @[sequencer-master.scala 652:39 sequencer-master.scala 265:66]
  wire  _GEN_26282 = 3'h0 == tail ? 1'h0 : _GEN_25872; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26283 = 3'h1 == tail ? 1'h0 : _GEN_25873; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26284 = 3'h2 == tail ? 1'h0 : _GEN_25874; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26285 = 3'h3 == tail ? 1'h0 : _GEN_25875; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26286 = 3'h4 == tail ? 1'h0 : _GEN_25876; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26287 = 3'h5 == tail ? 1'h0 : _GEN_25877; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26288 = 3'h6 == tail ? 1'h0 : _GEN_25878; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26289 = 3'h7 == tail ? 1'h0 : _GEN_25879; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26290 = 3'h0 == tail ? 1'h0 : _GEN_25880; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26291 = 3'h1 == tail ? 1'h0 : _GEN_25881; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26292 = 3'h2 == tail ? 1'h0 : _GEN_25882; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26293 = 3'h3 == tail ? 1'h0 : _GEN_25883; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26294 = 3'h4 == tail ? 1'h0 : _GEN_25884; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26295 = 3'h5 == tail ? 1'h0 : _GEN_25885; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26296 = 3'h6 == tail ? 1'h0 : _GEN_25886; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26297 = 3'h7 == tail ? 1'h0 : _GEN_25887; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26298 = 3'h0 == tail ? 1'h0 : _GEN_25888; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26299 = 3'h1 == tail ? 1'h0 : _GEN_25889; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26300 = 3'h2 == tail ? 1'h0 : _GEN_25890; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26301 = 3'h3 == tail ? 1'h0 : _GEN_25891; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26302 = 3'h4 == tail ? 1'h0 : _GEN_25892; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26303 = 3'h5 == tail ? 1'h0 : _GEN_25893; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26304 = 3'h6 == tail ? 1'h0 : _GEN_25894; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26305 = 3'h7 == tail ? 1'h0 : _GEN_25895; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26306 = 3'h0 == tail ? 1'h0 : _GEN_25896; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26307 = 3'h1 == tail ? 1'h0 : _GEN_25897; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26308 = 3'h2 == tail ? 1'h0 : _GEN_25898; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26309 = 3'h3 == tail ? 1'h0 : _GEN_25899; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26310 = 3'h4 == tail ? 1'h0 : _GEN_25900; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26311 = 3'h5 == tail ? 1'h0 : _GEN_25901; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26312 = 3'h6 == tail ? 1'h0 : _GEN_25902; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26313 = 3'h7 == tail ? 1'h0 : _GEN_25903; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26314 = 3'h0 == tail ? 1'h0 : _GEN_25904; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26315 = 3'h1 == tail ? 1'h0 : _GEN_25905; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26316 = 3'h2 == tail ? 1'h0 : _GEN_25906; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26317 = 3'h3 == tail ? 1'h0 : _GEN_25907; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26318 = 3'h4 == tail ? 1'h0 : _GEN_25908; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26319 = 3'h5 == tail ? 1'h0 : _GEN_25909; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26320 = 3'h6 == tail ? 1'h0 : _GEN_25910; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26321 = 3'h7 == tail ? 1'h0 : _GEN_25911; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26330 = 3'h0 == tail ? 1'h0 : _GEN_25920; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26331 = 3'h1 == tail ? 1'h0 : _GEN_25921; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26332 = 3'h2 == tail ? 1'h0 : _GEN_25922; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26333 = 3'h3 == tail ? 1'h0 : _GEN_25923; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26334 = 3'h4 == tail ? 1'h0 : _GEN_25924; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26335 = 3'h5 == tail ? 1'h0 : _GEN_25925; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26336 = 3'h6 == tail ? 1'h0 : _GEN_25926; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26337 = 3'h7 == tail ? 1'h0 : _GEN_25927; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26338 = 3'h0 == tail ? 1'h0 : _GEN_25928; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26339 = 3'h1 == tail ? 1'h0 : _GEN_25929; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26340 = 3'h2 == tail ? 1'h0 : _GEN_25930; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26341 = 3'h3 == tail ? 1'h0 : _GEN_25931; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26342 = 3'h4 == tail ? 1'h0 : _GEN_25932; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26343 = 3'h5 == tail ? 1'h0 : _GEN_25933; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26344 = 3'h6 == tail ? 1'h0 : _GEN_25934; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26345 = 3'h7 == tail ? 1'h0 : _GEN_25935; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26346 = 3'h0 == tail ? 1'h0 : _GEN_25936; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26347 = 3'h1 == tail ? 1'h0 : _GEN_25937; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26348 = 3'h2 == tail ? 1'h0 : _GEN_25938; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26349 = 3'h3 == tail ? 1'h0 : _GEN_25939; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26350 = 3'h4 == tail ? 1'h0 : _GEN_25940; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26351 = 3'h5 == tail ? 1'h0 : _GEN_25941; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26352 = 3'h6 == tail ? 1'h0 : _GEN_25942; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26353 = 3'h7 == tail ? 1'h0 : _GEN_25943; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26354 = 3'h0 == tail ? 1'h0 : _GEN_25944; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26355 = 3'h1 == tail ? 1'h0 : _GEN_25945; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26356 = 3'h2 == tail ? 1'h0 : _GEN_25946; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26357 = 3'h3 == tail ? 1'h0 : _GEN_25947; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26358 = 3'h4 == tail ? 1'h0 : _GEN_25948; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26359 = 3'h5 == tail ? 1'h0 : _GEN_25949; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26360 = 3'h6 == tail ? 1'h0 : _GEN_25950; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26361 = 3'h7 == tail ? 1'h0 : _GEN_25951; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26362 = 3'h0 == tail ? 1'h0 : _GEN_25952; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26363 = 3'h1 == tail ? 1'h0 : _GEN_25953; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26364 = 3'h2 == tail ? 1'h0 : _GEN_25954; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26365 = 3'h3 == tail ? 1'h0 : _GEN_25955; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26366 = 3'h4 == tail ? 1'h0 : _GEN_25956; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26367 = 3'h5 == tail ? 1'h0 : _GEN_25957; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26368 = 3'h6 == tail ? 1'h0 : _GEN_25958; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26369 = 3'h7 == tail ? 1'h0 : _GEN_25959; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26370 = 3'h0 == tail ? 1'h0 : _GEN_25960; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26371 = 3'h1 == tail ? 1'h0 : _GEN_25961; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26372 = 3'h2 == tail ? 1'h0 : _GEN_25962; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26373 = 3'h3 == tail ? 1'h0 : _GEN_25963; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26374 = 3'h4 == tail ? 1'h0 : _GEN_25964; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26375 = 3'h5 == tail ? 1'h0 : _GEN_25965; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26376 = 3'h6 == tail ? 1'h0 : _GEN_25966; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26377 = 3'h7 == tail ? 1'h0 : _GEN_25967; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26378 = 3'h0 == tail ? 1'h0 : _GEN_25968; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26379 = 3'h1 == tail ? 1'h0 : _GEN_25969; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26380 = 3'h2 == tail ? 1'h0 : _GEN_25970; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26381 = 3'h3 == tail ? 1'h0 : _GEN_25971; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26382 = 3'h4 == tail ? 1'h0 : _GEN_25972; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26383 = 3'h5 == tail ? 1'h0 : _GEN_25973; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26384 = 3'h6 == tail ? 1'h0 : _GEN_25974; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26385 = 3'h7 == tail ? 1'h0 : _GEN_25975; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26386 = 3'h0 == tail ? 1'h0 : _GEN_25976; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26387 = 3'h1 == tail ? 1'h0 : _GEN_25977; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26388 = 3'h2 == tail ? 1'h0 : _GEN_25978; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26389 = 3'h3 == tail ? 1'h0 : _GEN_25979; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26390 = 3'h4 == tail ? 1'h0 : _GEN_25980; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26391 = 3'h5 == tail ? 1'h0 : _GEN_25981; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26392 = 3'h6 == tail ? 1'h0 : _GEN_25982; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26393 = 3'h7 == tail ? 1'h0 : _GEN_25983; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26394 = 3'h0 == tail ? 1'h0 : _GEN_25984; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26395 = 3'h1 == tail ? 1'h0 : _GEN_25985; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26396 = 3'h2 == tail ? 1'h0 : _GEN_25986; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26397 = 3'h3 == tail ? 1'h0 : _GEN_25987; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26398 = 3'h4 == tail ? 1'h0 : _GEN_25988; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26399 = 3'h5 == tail ? 1'h0 : _GEN_25989; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26400 = 3'h6 == tail ? 1'h0 : _GEN_25990; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26401 = 3'h7 == tail ? 1'h0 : _GEN_25991; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26402 = 3'h0 == tail ? 1'h0 : _GEN_25992; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26403 = 3'h1 == tail ? 1'h0 : _GEN_25993; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26404 = 3'h2 == tail ? 1'h0 : _GEN_25994; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26405 = 3'h3 == tail ? 1'h0 : _GEN_25995; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26406 = 3'h4 == tail ? 1'h0 : _GEN_25996; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26407 = 3'h5 == tail ? 1'h0 : _GEN_25997; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26408 = 3'h6 == tail ? 1'h0 : _GEN_25998; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26409 = 3'h7 == tail ? 1'h0 : _GEN_25999; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26410 = 3'h0 == tail ? 1'h0 : _GEN_26000; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26411 = 3'h1 == tail ? 1'h0 : _GEN_26001; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26412 = 3'h2 == tail ? 1'h0 : _GEN_26002; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26413 = 3'h3 == tail ? 1'h0 : _GEN_26003; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26414 = 3'h4 == tail ? 1'h0 : _GEN_26004; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26415 = 3'h5 == tail ? 1'h0 : _GEN_26005; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26416 = 3'h6 == tail ? 1'h0 : _GEN_26006; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26417 = 3'h7 == tail ? 1'h0 : _GEN_26007; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26418 = 3'h0 == tail ? 1'h0 : _GEN_26008; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26419 = 3'h1 == tail ? 1'h0 : _GEN_26009; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26420 = 3'h2 == tail ? 1'h0 : _GEN_26010; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26421 = 3'h3 == tail ? 1'h0 : _GEN_26011; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26422 = 3'h4 == tail ? 1'h0 : _GEN_26012; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26423 = 3'h5 == tail ? 1'h0 : _GEN_26013; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26424 = 3'h6 == tail ? 1'h0 : _GEN_26014; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26425 = 3'h7 == tail ? 1'h0 : _GEN_26015; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26426 = 3'h0 == tail ? 1'h0 : _GEN_26016; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26427 = 3'h1 == tail ? 1'h0 : _GEN_26017; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26428 = 3'h2 == tail ? 1'h0 : _GEN_26018; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26429 = 3'h3 == tail ? 1'h0 : _GEN_26019; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26430 = 3'h4 == tail ? 1'h0 : _GEN_26020; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26431 = 3'h5 == tail ? 1'h0 : _GEN_26021; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26432 = 3'h6 == tail ? 1'h0 : _GEN_26022; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26433 = 3'h7 == tail ? 1'h0 : _GEN_26023; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26434 = 3'h0 == tail ? 1'h0 : _GEN_26024; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26435 = 3'h1 == tail ? 1'h0 : _GEN_26025; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26436 = 3'h2 == tail ? 1'h0 : _GEN_26026; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26437 = 3'h3 == tail ? 1'h0 : _GEN_26027; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26438 = 3'h4 == tail ? 1'h0 : _GEN_26028; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26439 = 3'h5 == tail ? 1'h0 : _GEN_26029; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26440 = 3'h6 == tail ? 1'h0 : _GEN_26030; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26441 = 3'h7 == tail ? 1'h0 : _GEN_26031; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26442 = 3'h0 == tail ? 1'h0 : _GEN_26032; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26443 = 3'h1 == tail ? 1'h0 : _GEN_26033; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26444 = 3'h2 == tail ? 1'h0 : _GEN_26034; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26445 = 3'h3 == tail ? 1'h0 : _GEN_26035; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26446 = 3'h4 == tail ? 1'h0 : _GEN_26036; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26447 = 3'h5 == tail ? 1'h0 : _GEN_26037; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26448 = 3'h6 == tail ? 1'h0 : _GEN_26038; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26449 = 3'h7 == tail ? 1'h0 : _GEN_26039; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26450 = 3'h0 == tail ? 1'h0 : _GEN_26040; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26451 = 3'h1 == tail ? 1'h0 : _GEN_26041; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26452 = 3'h2 == tail ? 1'h0 : _GEN_26042; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26453 = 3'h3 == tail ? 1'h0 : _GEN_26043; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26454 = 3'h4 == tail ? 1'h0 : _GEN_26044; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26455 = 3'h5 == tail ? 1'h0 : _GEN_26045; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26456 = 3'h6 == tail ? 1'h0 : _GEN_26046; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26457 = 3'h7 == tail ? 1'h0 : _GEN_26047; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26458 = 3'h0 == tail ? 1'h0 : _GEN_26048; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26459 = 3'h1 == tail ? 1'h0 : _GEN_26049; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26460 = 3'h2 == tail ? 1'h0 : _GEN_26050; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26461 = 3'h3 == tail ? 1'h0 : _GEN_26051; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26462 = 3'h4 == tail ? 1'h0 : _GEN_26052; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26463 = 3'h5 == tail ? 1'h0 : _GEN_26053; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26464 = 3'h6 == tail ? 1'h0 : _GEN_26054; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26465 = 3'h7 == tail ? 1'h0 : _GEN_26055; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26466 = 3'h0 == tail ? 1'h0 : _GEN_26056; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26467 = 3'h1 == tail ? 1'h0 : _GEN_26057; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26468 = 3'h2 == tail ? 1'h0 : _GEN_26058; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26469 = 3'h3 == tail ? 1'h0 : _GEN_26059; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26470 = 3'h4 == tail ? 1'h0 : _GEN_26060; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26471 = 3'h5 == tail ? 1'h0 : _GEN_26061; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26472 = 3'h6 == tail ? 1'h0 : _GEN_26062; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26473 = 3'h7 == tail ? 1'h0 : _GEN_26063; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26474 = 3'h0 == tail ? 1'h0 : _GEN_26064; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26475 = 3'h1 == tail ? 1'h0 : _GEN_26065; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26476 = 3'h2 == tail ? 1'h0 : _GEN_26066; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26477 = 3'h3 == tail ? 1'h0 : _GEN_26067; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26478 = 3'h4 == tail ? 1'h0 : _GEN_26068; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26479 = 3'h5 == tail ? 1'h0 : _GEN_26069; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26480 = 3'h6 == tail ? 1'h0 : _GEN_26070; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26481 = 3'h7 == tail ? 1'h0 : _GEN_26071; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26482 = 3'h0 == tail ? 1'h0 : _GEN_26072; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26483 = 3'h1 == tail ? 1'h0 : _GEN_26073; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26484 = 3'h2 == tail ? 1'h0 : _GEN_26074; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26485 = 3'h3 == tail ? 1'h0 : _GEN_26075; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26486 = 3'h4 == tail ? 1'h0 : _GEN_26076; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26487 = 3'h5 == tail ? 1'h0 : _GEN_26077; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26488 = 3'h6 == tail ? 1'h0 : _GEN_26078; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26489 = 3'h7 == tail ? 1'h0 : _GEN_26079; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26490 = 3'h0 == tail ? 1'h0 : _GEN_26080; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26491 = 3'h1 == tail ? 1'h0 : _GEN_26081; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26492 = 3'h2 == tail ? 1'h0 : _GEN_26082; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26493 = 3'h3 == tail ? 1'h0 : _GEN_26083; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26494 = 3'h4 == tail ? 1'h0 : _GEN_26084; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26495 = 3'h5 == tail ? 1'h0 : _GEN_26085; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26496 = 3'h6 == tail ? 1'h0 : _GEN_26086; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26497 = 3'h7 == tail ? 1'h0 : _GEN_26087; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26498 = 3'h0 == tail ? 1'h0 : _GEN_26088; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26499 = 3'h1 == tail ? 1'h0 : _GEN_26089; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26500 = 3'h2 == tail ? 1'h0 : _GEN_26090; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26501 = 3'h3 == tail ? 1'h0 : _GEN_26091; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26502 = 3'h4 == tail ? 1'h0 : _GEN_26092; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26503 = 3'h5 == tail ? 1'h0 : _GEN_26093; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26504 = 3'h6 == tail ? 1'h0 : _GEN_26094; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26505 = 3'h7 == tail ? 1'h0 : _GEN_26095; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26506 = 3'h0 == tail ? 1'h0 : _GEN_26096; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26507 = 3'h1 == tail ? 1'h0 : _GEN_26097; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26508 = 3'h2 == tail ? 1'h0 : _GEN_26098; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26509 = 3'h3 == tail ? 1'h0 : _GEN_26099; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26510 = 3'h4 == tail ? 1'h0 : _GEN_26100; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26511 = 3'h5 == tail ? 1'h0 : _GEN_26101; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26512 = 3'h6 == tail ? 1'h0 : _GEN_26102; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26513 = 3'h7 == tail ? 1'h0 : _GEN_26103; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26514 = 3'h0 == tail ? 1'h0 : _GEN_26104; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26515 = 3'h1 == tail ? 1'h0 : _GEN_26105; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26516 = 3'h2 == tail ? 1'h0 : _GEN_26106; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26517 = 3'h3 == tail ? 1'h0 : _GEN_26107; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26518 = 3'h4 == tail ? 1'h0 : _GEN_26108; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26519 = 3'h5 == tail ? 1'h0 : _GEN_26109; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26520 = 3'h6 == tail ? 1'h0 : _GEN_26110; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26521 = 3'h7 == tail ? 1'h0 : _GEN_26111; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26522 = 3'h0 == tail ? 1'h0 : _GEN_26112; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26523 = 3'h1 == tail ? 1'h0 : _GEN_26113; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26524 = 3'h2 == tail ? 1'h0 : _GEN_26114; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26525 = 3'h3 == tail ? 1'h0 : _GEN_26115; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26526 = 3'h4 == tail ? 1'h0 : _GEN_26116; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26527 = 3'h5 == tail ? 1'h0 : _GEN_26117; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26528 = 3'h6 == tail ? 1'h0 : _GEN_26118; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26529 = 3'h7 == tail ? 1'h0 : _GEN_26119; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_26538 = _GEN_32729 | e_0_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26539 = _GEN_32730 | e_1_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26540 = _GEN_32731 | e_2_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26541 = _GEN_32732 | e_3_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26542 = _GEN_32733 | e_4_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26543 = _GEN_32734 | e_5_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26544 = _GEN_32735 | e_6_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire  _GEN_26545 = _GEN_32736 | e_7_active_vpu; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26 sequencer-master.scala 109:14]
  wire [9:0] _GEN_26546 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_26136; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26547 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_26137; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26548 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_26138; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26549 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_26139; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26550 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_26140; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26551 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_26141; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26552 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_26142; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_26553 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_26143; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_26554 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_26144; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26555 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_26145; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26556 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_26146; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26557 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_26147; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26558 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_26148; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26559 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_26149; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26560 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_26150; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_26561 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_26151; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26562 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_26282; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26563 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_26283; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26564 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_26284; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26565 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_26285; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26566 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_26286; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26567 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_26287; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26568 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_26288; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26569 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_26289; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26570 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_26152; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26571 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_26153; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26572 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_26154; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26573 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_26155; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26574 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_26156; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26575 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_26157; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26576 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_26158; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26577 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_26159; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26578 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_26160; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26579 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_26161; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26580 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_26162; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26581 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_26163; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26582 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_26164; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26583 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_26165; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26584 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_26166; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_26585 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_26167; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_26586 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_26168; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26587 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_26169; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26588 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_26170; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26589 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_26171; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26590 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_26172; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26591 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_26173; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26592 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_26174; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_26593 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_26175; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_26594 = io_op_bits_base_vp_valid ? _GEN_26554 : _GEN_26144; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26595 = io_op_bits_base_vp_valid ? _GEN_26555 : _GEN_26145; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26596 = io_op_bits_base_vp_valid ? _GEN_26556 : _GEN_26146; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26597 = io_op_bits_base_vp_valid ? _GEN_26557 : _GEN_26147; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26598 = io_op_bits_base_vp_valid ? _GEN_26558 : _GEN_26148; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26599 = io_op_bits_base_vp_valid ? _GEN_26559 : _GEN_26149; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26600 = io_op_bits_base_vp_valid ? _GEN_26560 : _GEN_26150; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_26601 = io_op_bits_base_vp_valid ? _GEN_26561 : _GEN_26151; // @[sequencer-master.scala 320:41]
  wire  _GEN_26602 = io_op_bits_base_vp_valid ? _GEN_26562 : _GEN_26282; // @[sequencer-master.scala 320:41]
  wire  _GEN_26603 = io_op_bits_base_vp_valid ? _GEN_26563 : _GEN_26283; // @[sequencer-master.scala 320:41]
  wire  _GEN_26604 = io_op_bits_base_vp_valid ? _GEN_26564 : _GEN_26284; // @[sequencer-master.scala 320:41]
  wire  _GEN_26605 = io_op_bits_base_vp_valid ? _GEN_26565 : _GEN_26285; // @[sequencer-master.scala 320:41]
  wire  _GEN_26606 = io_op_bits_base_vp_valid ? _GEN_26566 : _GEN_26286; // @[sequencer-master.scala 320:41]
  wire  _GEN_26607 = io_op_bits_base_vp_valid ? _GEN_26567 : _GEN_26287; // @[sequencer-master.scala 320:41]
  wire  _GEN_26608 = io_op_bits_base_vp_valid ? _GEN_26568 : _GEN_26288; // @[sequencer-master.scala 320:41]
  wire  _GEN_26609 = io_op_bits_base_vp_valid ? _GEN_26569 : _GEN_26289; // @[sequencer-master.scala 320:41]
  wire  _GEN_26610 = io_op_bits_base_vp_valid ? _GEN_26570 : _GEN_26152; // @[sequencer-master.scala 320:41]
  wire  _GEN_26611 = io_op_bits_base_vp_valid ? _GEN_26571 : _GEN_26153; // @[sequencer-master.scala 320:41]
  wire  _GEN_26612 = io_op_bits_base_vp_valid ? _GEN_26572 : _GEN_26154; // @[sequencer-master.scala 320:41]
  wire  _GEN_26613 = io_op_bits_base_vp_valid ? _GEN_26573 : _GEN_26155; // @[sequencer-master.scala 320:41]
  wire  _GEN_26614 = io_op_bits_base_vp_valid ? _GEN_26574 : _GEN_26156; // @[sequencer-master.scala 320:41]
  wire  _GEN_26615 = io_op_bits_base_vp_valid ? _GEN_26575 : _GEN_26157; // @[sequencer-master.scala 320:41]
  wire  _GEN_26616 = io_op_bits_base_vp_valid ? _GEN_26576 : _GEN_26158; // @[sequencer-master.scala 320:41]
  wire  _GEN_26617 = io_op_bits_base_vp_valid ? _GEN_26577 : _GEN_26159; // @[sequencer-master.scala 320:41]
  wire  _GEN_26618 = io_op_bits_base_vp_valid ? _GEN_26578 : _GEN_26160; // @[sequencer-master.scala 320:41]
  wire  _GEN_26619 = io_op_bits_base_vp_valid ? _GEN_26579 : _GEN_26161; // @[sequencer-master.scala 320:41]
  wire  _GEN_26620 = io_op_bits_base_vp_valid ? _GEN_26580 : _GEN_26162; // @[sequencer-master.scala 320:41]
  wire  _GEN_26621 = io_op_bits_base_vp_valid ? _GEN_26581 : _GEN_26163; // @[sequencer-master.scala 320:41]
  wire  _GEN_26622 = io_op_bits_base_vp_valid ? _GEN_26582 : _GEN_26164; // @[sequencer-master.scala 320:41]
  wire  _GEN_26623 = io_op_bits_base_vp_valid ? _GEN_26583 : _GEN_26165; // @[sequencer-master.scala 320:41]
  wire  _GEN_26624 = io_op_bits_base_vp_valid ? _GEN_26584 : _GEN_26166; // @[sequencer-master.scala 320:41]
  wire  _GEN_26625 = io_op_bits_base_vp_valid ? _GEN_26585 : _GEN_26167; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26626 = io_op_bits_base_vp_valid ? _GEN_26586 : _GEN_26168; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26627 = io_op_bits_base_vp_valid ? _GEN_26587 : _GEN_26169; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26628 = io_op_bits_base_vp_valid ? _GEN_26588 : _GEN_26170; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26629 = io_op_bits_base_vp_valid ? _GEN_26589 : _GEN_26171; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26630 = io_op_bits_base_vp_valid ? _GEN_26590 : _GEN_26172; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26631 = io_op_bits_base_vp_valid ? _GEN_26591 : _GEN_26173; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26632 = io_op_bits_base_vp_valid ? _GEN_26592 : _GEN_26174; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_26633 = io_op_bits_base_vp_valid ? _GEN_26593 : _GEN_26175; // @[sequencer-master.scala 320:41]
  wire  _GEN_26634 = _GEN_32729 | _GEN_26330; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26635 = _GEN_32730 | _GEN_26331; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26636 = _GEN_32731 | _GEN_26332; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26637 = _GEN_32732 | _GEN_26333; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26638 = _GEN_32733 | _GEN_26334; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26639 = _GEN_32734 | _GEN_26335; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26640 = _GEN_32735 | _GEN_26336; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26641 = _GEN_32736 | _GEN_26337; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26642 = _T_26 ? _GEN_26634 : _GEN_26330; // @[sequencer-master.scala 154:24]
  wire  _GEN_26643 = _T_26 ? _GEN_26635 : _GEN_26331; // @[sequencer-master.scala 154:24]
  wire  _GEN_26644 = _T_26 ? _GEN_26636 : _GEN_26332; // @[sequencer-master.scala 154:24]
  wire  _GEN_26645 = _T_26 ? _GEN_26637 : _GEN_26333; // @[sequencer-master.scala 154:24]
  wire  _GEN_26646 = _T_26 ? _GEN_26638 : _GEN_26334; // @[sequencer-master.scala 154:24]
  wire  _GEN_26647 = _T_26 ? _GEN_26639 : _GEN_26335; // @[sequencer-master.scala 154:24]
  wire  _GEN_26648 = _T_26 ? _GEN_26640 : _GEN_26336; // @[sequencer-master.scala 154:24]
  wire  _GEN_26649 = _T_26 ? _GEN_26641 : _GEN_26337; // @[sequencer-master.scala 154:24]
  wire  _GEN_26650 = _GEN_32729 | _GEN_26354; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26651 = _GEN_32730 | _GEN_26355; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26652 = _GEN_32731 | _GEN_26356; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26653 = _GEN_32732 | _GEN_26357; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26654 = _GEN_32733 | _GEN_26358; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26655 = _GEN_32734 | _GEN_26359; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26656 = _GEN_32735 | _GEN_26360; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26657 = _GEN_32736 | _GEN_26361; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26658 = _T_48 ? _GEN_26650 : _GEN_26354; // @[sequencer-master.scala 154:24]
  wire  _GEN_26659 = _T_48 ? _GEN_26651 : _GEN_26355; // @[sequencer-master.scala 154:24]
  wire  _GEN_26660 = _T_48 ? _GEN_26652 : _GEN_26356; // @[sequencer-master.scala 154:24]
  wire  _GEN_26661 = _T_48 ? _GEN_26653 : _GEN_26357; // @[sequencer-master.scala 154:24]
  wire  _GEN_26662 = _T_48 ? _GEN_26654 : _GEN_26358; // @[sequencer-master.scala 154:24]
  wire  _GEN_26663 = _T_48 ? _GEN_26655 : _GEN_26359; // @[sequencer-master.scala 154:24]
  wire  _GEN_26664 = _T_48 ? _GEN_26656 : _GEN_26360; // @[sequencer-master.scala 154:24]
  wire  _GEN_26665 = _T_48 ? _GEN_26657 : _GEN_26361; // @[sequencer-master.scala 154:24]
  wire  _GEN_26666 = _GEN_32729 | _GEN_26378; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26667 = _GEN_32730 | _GEN_26379; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26668 = _GEN_32731 | _GEN_26380; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26669 = _GEN_32732 | _GEN_26381; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26670 = _GEN_32733 | _GEN_26382; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26671 = _GEN_32734 | _GEN_26383; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26672 = _GEN_32735 | _GEN_26384; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26673 = _GEN_32736 | _GEN_26385; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26674 = _T_70 ? _GEN_26666 : _GEN_26378; // @[sequencer-master.scala 154:24]
  wire  _GEN_26675 = _T_70 ? _GEN_26667 : _GEN_26379; // @[sequencer-master.scala 154:24]
  wire  _GEN_26676 = _T_70 ? _GEN_26668 : _GEN_26380; // @[sequencer-master.scala 154:24]
  wire  _GEN_26677 = _T_70 ? _GEN_26669 : _GEN_26381; // @[sequencer-master.scala 154:24]
  wire  _GEN_26678 = _T_70 ? _GEN_26670 : _GEN_26382; // @[sequencer-master.scala 154:24]
  wire  _GEN_26679 = _T_70 ? _GEN_26671 : _GEN_26383; // @[sequencer-master.scala 154:24]
  wire  _GEN_26680 = _T_70 ? _GEN_26672 : _GEN_26384; // @[sequencer-master.scala 154:24]
  wire  _GEN_26681 = _T_70 ? _GEN_26673 : _GEN_26385; // @[sequencer-master.scala 154:24]
  wire  _GEN_26682 = _GEN_32729 | _GEN_26402; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26683 = _GEN_32730 | _GEN_26403; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26684 = _GEN_32731 | _GEN_26404; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26685 = _GEN_32732 | _GEN_26405; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26686 = _GEN_32733 | _GEN_26406; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26687 = _GEN_32734 | _GEN_26407; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26688 = _GEN_32735 | _GEN_26408; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26689 = _GEN_32736 | _GEN_26409; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26690 = _T_92 ? _GEN_26682 : _GEN_26402; // @[sequencer-master.scala 154:24]
  wire  _GEN_26691 = _T_92 ? _GEN_26683 : _GEN_26403; // @[sequencer-master.scala 154:24]
  wire  _GEN_26692 = _T_92 ? _GEN_26684 : _GEN_26404; // @[sequencer-master.scala 154:24]
  wire  _GEN_26693 = _T_92 ? _GEN_26685 : _GEN_26405; // @[sequencer-master.scala 154:24]
  wire  _GEN_26694 = _T_92 ? _GEN_26686 : _GEN_26406; // @[sequencer-master.scala 154:24]
  wire  _GEN_26695 = _T_92 ? _GEN_26687 : _GEN_26407; // @[sequencer-master.scala 154:24]
  wire  _GEN_26696 = _T_92 ? _GEN_26688 : _GEN_26408; // @[sequencer-master.scala 154:24]
  wire  _GEN_26697 = _T_92 ? _GEN_26689 : _GEN_26409; // @[sequencer-master.scala 154:24]
  wire  _GEN_26698 = _GEN_32729 | _GEN_26426; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26699 = _GEN_32730 | _GEN_26427; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26700 = _GEN_32731 | _GEN_26428; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26701 = _GEN_32732 | _GEN_26429; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26702 = _GEN_32733 | _GEN_26430; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26703 = _GEN_32734 | _GEN_26431; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26704 = _GEN_32735 | _GEN_26432; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26705 = _GEN_32736 | _GEN_26433; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26706 = _T_114 ? _GEN_26698 : _GEN_26426; // @[sequencer-master.scala 154:24]
  wire  _GEN_26707 = _T_114 ? _GEN_26699 : _GEN_26427; // @[sequencer-master.scala 154:24]
  wire  _GEN_26708 = _T_114 ? _GEN_26700 : _GEN_26428; // @[sequencer-master.scala 154:24]
  wire  _GEN_26709 = _T_114 ? _GEN_26701 : _GEN_26429; // @[sequencer-master.scala 154:24]
  wire  _GEN_26710 = _T_114 ? _GEN_26702 : _GEN_26430; // @[sequencer-master.scala 154:24]
  wire  _GEN_26711 = _T_114 ? _GEN_26703 : _GEN_26431; // @[sequencer-master.scala 154:24]
  wire  _GEN_26712 = _T_114 ? _GEN_26704 : _GEN_26432; // @[sequencer-master.scala 154:24]
  wire  _GEN_26713 = _T_114 ? _GEN_26705 : _GEN_26433; // @[sequencer-master.scala 154:24]
  wire  _GEN_26714 = _GEN_32729 | _GEN_26450; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26715 = _GEN_32730 | _GEN_26451; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26716 = _GEN_32731 | _GEN_26452; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26717 = _GEN_32732 | _GEN_26453; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26718 = _GEN_32733 | _GEN_26454; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26719 = _GEN_32734 | _GEN_26455; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26720 = _GEN_32735 | _GEN_26456; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26721 = _GEN_32736 | _GEN_26457; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26722 = _T_136 ? _GEN_26714 : _GEN_26450; // @[sequencer-master.scala 154:24]
  wire  _GEN_26723 = _T_136 ? _GEN_26715 : _GEN_26451; // @[sequencer-master.scala 154:24]
  wire  _GEN_26724 = _T_136 ? _GEN_26716 : _GEN_26452; // @[sequencer-master.scala 154:24]
  wire  _GEN_26725 = _T_136 ? _GEN_26717 : _GEN_26453; // @[sequencer-master.scala 154:24]
  wire  _GEN_26726 = _T_136 ? _GEN_26718 : _GEN_26454; // @[sequencer-master.scala 154:24]
  wire  _GEN_26727 = _T_136 ? _GEN_26719 : _GEN_26455; // @[sequencer-master.scala 154:24]
  wire  _GEN_26728 = _T_136 ? _GEN_26720 : _GEN_26456; // @[sequencer-master.scala 154:24]
  wire  _GEN_26729 = _T_136 ? _GEN_26721 : _GEN_26457; // @[sequencer-master.scala 154:24]
  wire  _GEN_26730 = _GEN_32729 | _GEN_26474; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26731 = _GEN_32730 | _GEN_26475; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26732 = _GEN_32731 | _GEN_26476; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26733 = _GEN_32732 | _GEN_26477; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26734 = _GEN_32733 | _GEN_26478; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26735 = _GEN_32734 | _GEN_26479; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26736 = _GEN_32735 | _GEN_26480; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26737 = _GEN_32736 | _GEN_26481; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26738 = _T_158 ? _GEN_26730 : _GEN_26474; // @[sequencer-master.scala 154:24]
  wire  _GEN_26739 = _T_158 ? _GEN_26731 : _GEN_26475; // @[sequencer-master.scala 154:24]
  wire  _GEN_26740 = _T_158 ? _GEN_26732 : _GEN_26476; // @[sequencer-master.scala 154:24]
  wire  _GEN_26741 = _T_158 ? _GEN_26733 : _GEN_26477; // @[sequencer-master.scala 154:24]
  wire  _GEN_26742 = _T_158 ? _GEN_26734 : _GEN_26478; // @[sequencer-master.scala 154:24]
  wire  _GEN_26743 = _T_158 ? _GEN_26735 : _GEN_26479; // @[sequencer-master.scala 154:24]
  wire  _GEN_26744 = _T_158 ? _GEN_26736 : _GEN_26480; // @[sequencer-master.scala 154:24]
  wire  _GEN_26745 = _T_158 ? _GEN_26737 : _GEN_26481; // @[sequencer-master.scala 154:24]
  wire  _GEN_26746 = _GEN_32729 | _GEN_26498; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26747 = _GEN_32730 | _GEN_26499; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26748 = _GEN_32731 | _GEN_26500; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26749 = _GEN_32732 | _GEN_26501; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26750 = _GEN_32733 | _GEN_26502; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26751 = _GEN_32734 | _GEN_26503; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26752 = _GEN_32735 | _GEN_26504; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26753 = _GEN_32736 | _GEN_26505; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_26754 = _T_180 ? _GEN_26746 : _GEN_26498; // @[sequencer-master.scala 154:24]
  wire  _GEN_26755 = _T_180 ? _GEN_26747 : _GEN_26499; // @[sequencer-master.scala 154:24]
  wire  _GEN_26756 = _T_180 ? _GEN_26748 : _GEN_26500; // @[sequencer-master.scala 154:24]
  wire  _GEN_26757 = _T_180 ? _GEN_26749 : _GEN_26501; // @[sequencer-master.scala 154:24]
  wire  _GEN_26758 = _T_180 ? _GEN_26750 : _GEN_26502; // @[sequencer-master.scala 154:24]
  wire  _GEN_26759 = _T_180 ? _GEN_26751 : _GEN_26503; // @[sequencer-master.scala 154:24]
  wire  _GEN_26760 = _T_180 ? _GEN_26752 : _GEN_26504; // @[sequencer-master.scala 154:24]
  wire  _GEN_26761 = _T_180 ? _GEN_26753 : _GEN_26505; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_26762 = 3'h0 == tail ? 2'h0 : _GEN_26224; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26763 = 3'h1 == tail ? 2'h0 : _GEN_26225; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26764 = 3'h2 == tail ? 2'h0 : _GEN_26226; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26765 = 3'h3 == tail ? 2'h0 : _GEN_26227; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26766 = 3'h4 == tail ? 2'h0 : _GEN_26228; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26767 = 3'h5 == tail ? 2'h0 : _GEN_26229; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26768 = 3'h6 == tail ? 2'h0 : _GEN_26230; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_26769 = 3'h7 == tail ? 2'h0 : _GEN_26231; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_26770 = 3'h0 == tail ? 4'h0 : _GEN_26232; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26771 = 3'h1 == tail ? 4'h0 : _GEN_26233; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26772 = 3'h2 == tail ? 4'h0 : _GEN_26234; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26773 = 3'h3 == tail ? 4'h0 : _GEN_26235; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26774 = 3'h4 == tail ? 4'h0 : _GEN_26236; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26775 = 3'h5 == tail ? 4'h0 : _GEN_26237; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26776 = 3'h6 == tail ? 4'h0 : _GEN_26238; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_26777 = 3'h7 == tail ? 4'h0 : _GEN_26239; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_26778 = 3'h0 == tail ? 3'h0 : _GEN_26240; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26779 = 3'h1 == tail ? 3'h0 : _GEN_26241; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26780 = 3'h2 == tail ? 3'h0 : _GEN_26242; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26781 = 3'h3 == tail ? 3'h0 : _GEN_26243; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26782 = 3'h4 == tail ? 3'h0 : _GEN_26244; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26783 = 3'h5 == tail ? 3'h0 : _GEN_26245; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26784 = 3'h6 == tail ? 3'h0 : _GEN_26246; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_26785 = 3'h7 == tail ? 3'h0 : _GEN_26247; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_26802 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26602; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26803 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26603; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26804 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26604; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26805 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26605; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26806 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26606; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26807 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26607; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26808 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26608; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26809 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26609; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_26810 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26290; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26811 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26291; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26812 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26292; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26813 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26293; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26814 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26294; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26815 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26295; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26816 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26296; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26817 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26297; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_26818 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26298; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26819 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26299; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26820 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26300; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26821 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26301; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26822 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26302; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26823 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26303; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26824 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26304; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26825 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26305; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_26826 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26306; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26827 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26307; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26828 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26308; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26829 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26309; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26830 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26310; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26831 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26311; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26832 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26312; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26833 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26313; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_26834 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26314; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26835 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26315; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26836 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26316; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26837 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26317; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26838 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26318; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26839 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26319; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26840 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26320; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26841 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26321; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_26850 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26642; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26851 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26643; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26852 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26644; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26853 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26645; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26854 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26646; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26855 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26647; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26856 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26648; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26857 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26649; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26858 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26338; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26859 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26339; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26860 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26340; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26861 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26341; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26862 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26342; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26863 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26343; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26864 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26344; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26865 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26345; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26866 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26346; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26867 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26347; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26868 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26348; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26869 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26349; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26870 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26350; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26871 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26351; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26872 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26352; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26873 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26353; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26874 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26658; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26875 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26659; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26876 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26660; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26877 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26661; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26878 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26662; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26879 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26663; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26880 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26664; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26881 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26665; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26882 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26362; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26883 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26363; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26884 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26364; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26885 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26365; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26886 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26366; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26887 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26367; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26888 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26368; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26889 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26369; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26890 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26370; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26891 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26371; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26892 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26372; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26893 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26373; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26894 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26374; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26895 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26375; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26896 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26376; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26897 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26377; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26898 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26674; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26899 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26675; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26900 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26676; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26901 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26677; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26902 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26678; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26903 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26679; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26904 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26680; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26905 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26681; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26906 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26386; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26907 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26387; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26908 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26388; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26909 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26389; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26910 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26390; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26911 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26391; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26912 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26392; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26913 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26393; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26914 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26394; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26915 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26395; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26916 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26396; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26917 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26397; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26918 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26398; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26919 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26399; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26920 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26400; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26921 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26401; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26922 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26690; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26923 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26691; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26924 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26692; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26925 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26693; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26926 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26694; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26927 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26695; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26928 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26696; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26929 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26697; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26930 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26410; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26931 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26411; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26932 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26412; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26933 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26413; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26934 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26414; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26935 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26415; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26936 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26416; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26937 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26417; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26938 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26418; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26939 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26419; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26940 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26420; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26941 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26421; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26942 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26422; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26943 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26423; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26944 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26424; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26945 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26425; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26946 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26706; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26947 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26707; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26948 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26708; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26949 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26709; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26950 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26710; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26951 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26711; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26952 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26712; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26953 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26713; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26954 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26434; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26955 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26435; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26956 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26436; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26957 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26437; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26958 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26438; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26959 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26439; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26960 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26440; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26961 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26441; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26962 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26442; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26963 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26443; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26964 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26444; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26965 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26445; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26966 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26446; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26967 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26447; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26968 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26448; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26969 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26449; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26970 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26722; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26971 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26723; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26972 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26724; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26973 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26725; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26974 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26726; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26975 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26727; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26976 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26728; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26977 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26729; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26978 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26458; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26979 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26459; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26980 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26460; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26981 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26461; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26982 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26462; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26983 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26463; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26984 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26464; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26985 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26465; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_26986 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26466; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26987 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26467; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26988 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26468; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26989 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26469; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26990 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26470; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26991 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26471; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26992 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26472; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26993 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26473; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_26994 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26738; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26995 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26739; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26996 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26740; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26997 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26741; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26998 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26742; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_26999 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26743; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27000 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26744; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27001 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26745; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27002 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26482; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27003 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26483; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27004 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26484; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27005 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26485; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27006 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26486; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27007 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26487; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27008 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26488; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27009 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26489; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27010 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26490; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27011 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26491; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27012 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26492; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27013 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26493; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27014 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26494; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27015 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26495; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27016 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26496; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27017 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26497; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27018 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26754; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27019 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26755; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27020 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26756; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27021 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26757; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27022 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26758; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27023 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26759; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27024 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26760; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27025 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26761; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27026 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26506; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27027 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26507; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27028 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26508; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27029 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26509; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27030 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26510; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27031 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26511; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27032 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26512; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27033 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26513; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27034 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26514; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27035 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26515; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27036 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26516; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27037 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26517; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27038 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26518; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27039 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26519; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27040 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26520; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27041 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26521; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27042 = 3'h0 == _T_1645 ? 1'h0 : _GEN_26522; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27043 = 3'h1 == _T_1645 ? 1'h0 : _GEN_26523; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27044 = 3'h2 == _T_1645 ? 1'h0 : _GEN_26524; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27045 = 3'h3 == _T_1645 ? 1'h0 : _GEN_26525; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27046 = 3'h4 == _T_1645 ? 1'h0 : _GEN_26526; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27047 = 3'h5 == _T_1645 ? 1'h0 : _GEN_26527; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27048 = 3'h6 == _T_1645 ? 1'h0 : _GEN_26528; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27049 = 3'h7 == _T_1645 ? 1'h0 : _GEN_26529; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27058 = _GEN_34121 | _GEN_26248; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27059 = _GEN_34122 | _GEN_26249; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27060 = _GEN_34123 | _GEN_26250; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27061 = _GEN_34124 | _GEN_26251; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27062 = _GEN_34125 | _GEN_26252; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27063 = _GEN_34126 | _GEN_26253; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27064 = _GEN_34127 | _GEN_26254; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27065 = _GEN_34128 | _GEN_26255; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_27066 = 3'h0 == _T_1645 ? io_op_bits_fn_union : _GEN_26546; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27067 = 3'h1 == _T_1645 ? io_op_bits_fn_union : _GEN_26547; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27068 = 3'h2 == _T_1645 ? io_op_bits_fn_union : _GEN_26548; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27069 = 3'h3 == _T_1645 ? io_op_bits_fn_union : _GEN_26549; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27070 = 3'h4 == _T_1645 ? io_op_bits_fn_union : _GEN_26550; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27071 = 3'h5 == _T_1645 ? io_op_bits_fn_union : _GEN_26551; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27072 = 3'h6 == _T_1645 ? io_op_bits_fn_union : _GEN_26552; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27073 = 3'h7 == _T_1645 ? io_op_bits_fn_union : _GEN_26553; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [1:0] _GEN_27074 = 3'h0 == _T_1645 ? 2'h0 : _GEN_26762; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27075 = 3'h1 == _T_1645 ? 2'h0 : _GEN_26763; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27076 = 3'h2 == _T_1645 ? 2'h0 : _GEN_26764; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27077 = 3'h3 == _T_1645 ? 2'h0 : _GEN_26765; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27078 = 3'h4 == _T_1645 ? 2'h0 : _GEN_26766; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27079 = 3'h5 == _T_1645 ? 2'h0 : _GEN_26767; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27080 = 3'h6 == _T_1645 ? 2'h0 : _GEN_26768; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27081 = 3'h7 == _T_1645 ? 2'h0 : _GEN_26769; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_27082 = 3'h0 == _T_1645 ? 4'h0 : _GEN_26770; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27083 = 3'h1 == _T_1645 ? 4'h0 : _GEN_26771; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27084 = 3'h2 == _T_1645 ? 4'h0 : _GEN_26772; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27085 = 3'h3 == _T_1645 ? 4'h0 : _GEN_26773; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27086 = 3'h4 == _T_1645 ? 4'h0 : _GEN_26774; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27087 = 3'h5 == _T_1645 ? 4'h0 : _GEN_26775; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27088 = 3'h6 == _T_1645 ? 4'h0 : _GEN_26776; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_27089 = 3'h7 == _T_1645 ? 4'h0 : _GEN_26777; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_27090 = 3'h0 == _T_1645 ? 3'h0 : _GEN_26778; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27091 = 3'h1 == _T_1645 ? 3'h0 : _GEN_26779; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27092 = 3'h2 == _T_1645 ? 3'h0 : _GEN_26780; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27093 = 3'h3 == _T_1645 ? 3'h0 : _GEN_26781; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27094 = 3'h4 == _T_1645 ? 3'h0 : _GEN_26782; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27095 = 3'h5 == _T_1645 ? 3'h0 : _GEN_26783; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27096 = 3'h6 == _T_1645 ? 3'h0 : _GEN_26784; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_27097 = 3'h7 == _T_1645 ? 3'h0 : _GEN_26785; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_27098 = _GEN_34121 | _GEN_26858; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27099 = _GEN_34122 | _GEN_26859; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27100 = _GEN_34123 | _GEN_26860; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27101 = _GEN_34124 | _GEN_26861; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27102 = _GEN_34125 | _GEN_26862; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27103 = _GEN_34126 | _GEN_26863; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27104 = _GEN_34127 | _GEN_26864; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27105 = _GEN_34128 | _GEN_26865; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27106 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27098 : _GEN_26858; // @[sequencer-master.scala 161:86]
  wire  _GEN_27107 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27099 : _GEN_26859; // @[sequencer-master.scala 161:86]
  wire  _GEN_27108 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27100 : _GEN_26860; // @[sequencer-master.scala 161:86]
  wire  _GEN_27109 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27101 : _GEN_26861; // @[sequencer-master.scala 161:86]
  wire  _GEN_27110 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27102 : _GEN_26862; // @[sequencer-master.scala 161:86]
  wire  _GEN_27111 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27103 : _GEN_26863; // @[sequencer-master.scala 161:86]
  wire  _GEN_27112 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27104 : _GEN_26864; // @[sequencer-master.scala 161:86]
  wire  _GEN_27113 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27105 : _GEN_26865; // @[sequencer-master.scala 161:86]
  wire  _GEN_27114 = _GEN_34121 | _GEN_26882; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27115 = _GEN_34122 | _GEN_26883; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27116 = _GEN_34123 | _GEN_26884; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27117 = _GEN_34124 | _GEN_26885; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27118 = _GEN_34125 | _GEN_26886; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27119 = _GEN_34126 | _GEN_26887; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27120 = _GEN_34127 | _GEN_26888; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27121 = _GEN_34128 | _GEN_26889; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27122 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27114 : _GEN_26882; // @[sequencer-master.scala 161:86]
  wire  _GEN_27123 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27115 : _GEN_26883; // @[sequencer-master.scala 161:86]
  wire  _GEN_27124 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27116 : _GEN_26884; // @[sequencer-master.scala 161:86]
  wire  _GEN_27125 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27117 : _GEN_26885; // @[sequencer-master.scala 161:86]
  wire  _GEN_27126 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27118 : _GEN_26886; // @[sequencer-master.scala 161:86]
  wire  _GEN_27127 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27119 : _GEN_26887; // @[sequencer-master.scala 161:86]
  wire  _GEN_27128 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27120 : _GEN_26888; // @[sequencer-master.scala 161:86]
  wire  _GEN_27129 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27121 : _GEN_26889; // @[sequencer-master.scala 161:86]
  wire  _GEN_27130 = _GEN_34121 | _GEN_26906; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27131 = _GEN_34122 | _GEN_26907; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27132 = _GEN_34123 | _GEN_26908; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27133 = _GEN_34124 | _GEN_26909; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27134 = _GEN_34125 | _GEN_26910; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27135 = _GEN_34126 | _GEN_26911; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27136 = _GEN_34127 | _GEN_26912; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27137 = _GEN_34128 | _GEN_26913; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27138 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27130 : _GEN_26906; // @[sequencer-master.scala 161:86]
  wire  _GEN_27139 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27131 : _GEN_26907; // @[sequencer-master.scala 161:86]
  wire  _GEN_27140 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27132 : _GEN_26908; // @[sequencer-master.scala 161:86]
  wire  _GEN_27141 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27133 : _GEN_26909; // @[sequencer-master.scala 161:86]
  wire  _GEN_27142 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27134 : _GEN_26910; // @[sequencer-master.scala 161:86]
  wire  _GEN_27143 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27135 : _GEN_26911; // @[sequencer-master.scala 161:86]
  wire  _GEN_27144 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27136 : _GEN_26912; // @[sequencer-master.scala 161:86]
  wire  _GEN_27145 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27137 : _GEN_26913; // @[sequencer-master.scala 161:86]
  wire  _GEN_27146 = _GEN_34121 | _GEN_26930; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27147 = _GEN_34122 | _GEN_26931; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27148 = _GEN_34123 | _GEN_26932; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27149 = _GEN_34124 | _GEN_26933; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27150 = _GEN_34125 | _GEN_26934; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27151 = _GEN_34126 | _GEN_26935; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27152 = _GEN_34127 | _GEN_26936; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27153 = _GEN_34128 | _GEN_26937; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27154 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27146 : _GEN_26930; // @[sequencer-master.scala 161:86]
  wire  _GEN_27155 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27147 : _GEN_26931; // @[sequencer-master.scala 161:86]
  wire  _GEN_27156 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27148 : _GEN_26932; // @[sequencer-master.scala 161:86]
  wire  _GEN_27157 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27149 : _GEN_26933; // @[sequencer-master.scala 161:86]
  wire  _GEN_27158 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27150 : _GEN_26934; // @[sequencer-master.scala 161:86]
  wire  _GEN_27159 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27151 : _GEN_26935; // @[sequencer-master.scala 161:86]
  wire  _GEN_27160 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27152 : _GEN_26936; // @[sequencer-master.scala 161:86]
  wire  _GEN_27161 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27153 : _GEN_26937; // @[sequencer-master.scala 161:86]
  wire  _GEN_27162 = _GEN_34121 | _GEN_26954; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27163 = _GEN_34122 | _GEN_26955; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27164 = _GEN_34123 | _GEN_26956; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27165 = _GEN_34124 | _GEN_26957; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27166 = _GEN_34125 | _GEN_26958; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27167 = _GEN_34126 | _GEN_26959; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27168 = _GEN_34127 | _GEN_26960; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27169 = _GEN_34128 | _GEN_26961; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27170 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27162 : _GEN_26954; // @[sequencer-master.scala 161:86]
  wire  _GEN_27171 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27163 : _GEN_26955; // @[sequencer-master.scala 161:86]
  wire  _GEN_27172 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27164 : _GEN_26956; // @[sequencer-master.scala 161:86]
  wire  _GEN_27173 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27165 : _GEN_26957; // @[sequencer-master.scala 161:86]
  wire  _GEN_27174 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27166 : _GEN_26958; // @[sequencer-master.scala 161:86]
  wire  _GEN_27175 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27167 : _GEN_26959; // @[sequencer-master.scala 161:86]
  wire  _GEN_27176 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27168 : _GEN_26960; // @[sequencer-master.scala 161:86]
  wire  _GEN_27177 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27169 : _GEN_26961; // @[sequencer-master.scala 161:86]
  wire  _GEN_27178 = _GEN_34121 | _GEN_26978; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27179 = _GEN_34122 | _GEN_26979; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27180 = _GEN_34123 | _GEN_26980; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27181 = _GEN_34124 | _GEN_26981; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27182 = _GEN_34125 | _GEN_26982; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27183 = _GEN_34126 | _GEN_26983; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27184 = _GEN_34127 | _GEN_26984; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27185 = _GEN_34128 | _GEN_26985; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27186 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27178 : _GEN_26978; // @[sequencer-master.scala 161:86]
  wire  _GEN_27187 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27179 : _GEN_26979; // @[sequencer-master.scala 161:86]
  wire  _GEN_27188 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27180 : _GEN_26980; // @[sequencer-master.scala 161:86]
  wire  _GEN_27189 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27181 : _GEN_26981; // @[sequencer-master.scala 161:86]
  wire  _GEN_27190 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27182 : _GEN_26982; // @[sequencer-master.scala 161:86]
  wire  _GEN_27191 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27183 : _GEN_26983; // @[sequencer-master.scala 161:86]
  wire  _GEN_27192 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27184 : _GEN_26984; // @[sequencer-master.scala 161:86]
  wire  _GEN_27193 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27185 : _GEN_26985; // @[sequencer-master.scala 161:86]
  wire  _GEN_27194 = _GEN_34121 | _GEN_27002; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27195 = _GEN_34122 | _GEN_27003; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27196 = _GEN_34123 | _GEN_27004; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27197 = _GEN_34124 | _GEN_27005; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27198 = _GEN_34125 | _GEN_27006; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27199 = _GEN_34126 | _GEN_27007; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27200 = _GEN_34127 | _GEN_27008; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27201 = _GEN_34128 | _GEN_27009; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27202 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27194 : _GEN_27002; // @[sequencer-master.scala 161:86]
  wire  _GEN_27203 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27195 : _GEN_27003; // @[sequencer-master.scala 161:86]
  wire  _GEN_27204 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27196 : _GEN_27004; // @[sequencer-master.scala 161:86]
  wire  _GEN_27205 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27197 : _GEN_27005; // @[sequencer-master.scala 161:86]
  wire  _GEN_27206 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27198 : _GEN_27006; // @[sequencer-master.scala 161:86]
  wire  _GEN_27207 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27199 : _GEN_27007; // @[sequencer-master.scala 161:86]
  wire  _GEN_27208 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27200 : _GEN_27008; // @[sequencer-master.scala 161:86]
  wire  _GEN_27209 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27201 : _GEN_27009; // @[sequencer-master.scala 161:86]
  wire  _GEN_27210 = _GEN_34121 | _GEN_27026; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27211 = _GEN_34122 | _GEN_27027; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27212 = _GEN_34123 | _GEN_27028; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27213 = _GEN_34124 | _GEN_27029; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27214 = _GEN_34125 | _GEN_27030; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27215 = _GEN_34126 | _GEN_27031; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27216 = _GEN_34127 | _GEN_27032; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27217 = _GEN_34128 | _GEN_27033; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27218 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27210 : _GEN_27026; // @[sequencer-master.scala 161:86]
  wire  _GEN_27219 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27211 : _GEN_27027; // @[sequencer-master.scala 161:86]
  wire  _GEN_27220 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27212 : _GEN_27028; // @[sequencer-master.scala 161:86]
  wire  _GEN_27221 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27213 : _GEN_27029; // @[sequencer-master.scala 161:86]
  wire  _GEN_27222 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27214 : _GEN_27030; // @[sequencer-master.scala 161:86]
  wire  _GEN_27223 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27215 : _GEN_27031; // @[sequencer-master.scala 161:86]
  wire  _GEN_27224 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27216 : _GEN_27032; // @[sequencer-master.scala 161:86]
  wire  _GEN_27225 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27217 : _GEN_27033; // @[sequencer-master.scala 161:86]
  wire  _GEN_27226 = _GEN_34121 | _GEN_26866; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27227 = _GEN_34122 | _GEN_26867; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27228 = _GEN_34123 | _GEN_26868; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27229 = _GEN_34124 | _GEN_26869; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27230 = _GEN_34125 | _GEN_26870; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27231 = _GEN_34126 | _GEN_26871; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27232 = _GEN_34127 | _GEN_26872; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27233 = _GEN_34128 | _GEN_26873; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27234 = _T_1442 ? _GEN_27226 : _GEN_26866; // @[sequencer-master.scala 168:32]
  wire  _GEN_27235 = _T_1442 ? _GEN_27227 : _GEN_26867; // @[sequencer-master.scala 168:32]
  wire  _GEN_27236 = _T_1442 ? _GEN_27228 : _GEN_26868; // @[sequencer-master.scala 168:32]
  wire  _GEN_27237 = _T_1442 ? _GEN_27229 : _GEN_26869; // @[sequencer-master.scala 168:32]
  wire  _GEN_27238 = _T_1442 ? _GEN_27230 : _GEN_26870; // @[sequencer-master.scala 168:32]
  wire  _GEN_27239 = _T_1442 ? _GEN_27231 : _GEN_26871; // @[sequencer-master.scala 168:32]
  wire  _GEN_27240 = _T_1442 ? _GEN_27232 : _GEN_26872; // @[sequencer-master.scala 168:32]
  wire  _GEN_27241 = _T_1442 ? _GEN_27233 : _GEN_26873; // @[sequencer-master.scala 168:32]
  wire  _GEN_27242 = _GEN_34121 | _GEN_26890; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27243 = _GEN_34122 | _GEN_26891; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27244 = _GEN_34123 | _GEN_26892; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27245 = _GEN_34124 | _GEN_26893; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27246 = _GEN_34125 | _GEN_26894; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27247 = _GEN_34126 | _GEN_26895; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27248 = _GEN_34127 | _GEN_26896; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27249 = _GEN_34128 | _GEN_26897; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27250 = _T_1464 ? _GEN_27242 : _GEN_26890; // @[sequencer-master.scala 168:32]
  wire  _GEN_27251 = _T_1464 ? _GEN_27243 : _GEN_26891; // @[sequencer-master.scala 168:32]
  wire  _GEN_27252 = _T_1464 ? _GEN_27244 : _GEN_26892; // @[sequencer-master.scala 168:32]
  wire  _GEN_27253 = _T_1464 ? _GEN_27245 : _GEN_26893; // @[sequencer-master.scala 168:32]
  wire  _GEN_27254 = _T_1464 ? _GEN_27246 : _GEN_26894; // @[sequencer-master.scala 168:32]
  wire  _GEN_27255 = _T_1464 ? _GEN_27247 : _GEN_26895; // @[sequencer-master.scala 168:32]
  wire  _GEN_27256 = _T_1464 ? _GEN_27248 : _GEN_26896; // @[sequencer-master.scala 168:32]
  wire  _GEN_27257 = _T_1464 ? _GEN_27249 : _GEN_26897; // @[sequencer-master.scala 168:32]
  wire  _GEN_27258 = _GEN_34121 | _GEN_26914; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27259 = _GEN_34122 | _GEN_26915; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27260 = _GEN_34123 | _GEN_26916; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27261 = _GEN_34124 | _GEN_26917; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27262 = _GEN_34125 | _GEN_26918; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27263 = _GEN_34126 | _GEN_26919; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27264 = _GEN_34127 | _GEN_26920; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27265 = _GEN_34128 | _GEN_26921; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27266 = _T_1486 ? _GEN_27258 : _GEN_26914; // @[sequencer-master.scala 168:32]
  wire  _GEN_27267 = _T_1486 ? _GEN_27259 : _GEN_26915; // @[sequencer-master.scala 168:32]
  wire  _GEN_27268 = _T_1486 ? _GEN_27260 : _GEN_26916; // @[sequencer-master.scala 168:32]
  wire  _GEN_27269 = _T_1486 ? _GEN_27261 : _GEN_26917; // @[sequencer-master.scala 168:32]
  wire  _GEN_27270 = _T_1486 ? _GEN_27262 : _GEN_26918; // @[sequencer-master.scala 168:32]
  wire  _GEN_27271 = _T_1486 ? _GEN_27263 : _GEN_26919; // @[sequencer-master.scala 168:32]
  wire  _GEN_27272 = _T_1486 ? _GEN_27264 : _GEN_26920; // @[sequencer-master.scala 168:32]
  wire  _GEN_27273 = _T_1486 ? _GEN_27265 : _GEN_26921; // @[sequencer-master.scala 168:32]
  wire  _GEN_27274 = _GEN_34121 | _GEN_26938; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27275 = _GEN_34122 | _GEN_26939; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27276 = _GEN_34123 | _GEN_26940; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27277 = _GEN_34124 | _GEN_26941; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27278 = _GEN_34125 | _GEN_26942; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27279 = _GEN_34126 | _GEN_26943; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27280 = _GEN_34127 | _GEN_26944; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27281 = _GEN_34128 | _GEN_26945; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27282 = _T_1508 ? _GEN_27274 : _GEN_26938; // @[sequencer-master.scala 168:32]
  wire  _GEN_27283 = _T_1508 ? _GEN_27275 : _GEN_26939; // @[sequencer-master.scala 168:32]
  wire  _GEN_27284 = _T_1508 ? _GEN_27276 : _GEN_26940; // @[sequencer-master.scala 168:32]
  wire  _GEN_27285 = _T_1508 ? _GEN_27277 : _GEN_26941; // @[sequencer-master.scala 168:32]
  wire  _GEN_27286 = _T_1508 ? _GEN_27278 : _GEN_26942; // @[sequencer-master.scala 168:32]
  wire  _GEN_27287 = _T_1508 ? _GEN_27279 : _GEN_26943; // @[sequencer-master.scala 168:32]
  wire  _GEN_27288 = _T_1508 ? _GEN_27280 : _GEN_26944; // @[sequencer-master.scala 168:32]
  wire  _GEN_27289 = _T_1508 ? _GEN_27281 : _GEN_26945; // @[sequencer-master.scala 168:32]
  wire  _GEN_27290 = _GEN_34121 | _GEN_26962; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27291 = _GEN_34122 | _GEN_26963; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27292 = _GEN_34123 | _GEN_26964; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27293 = _GEN_34124 | _GEN_26965; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27294 = _GEN_34125 | _GEN_26966; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27295 = _GEN_34126 | _GEN_26967; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27296 = _GEN_34127 | _GEN_26968; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27297 = _GEN_34128 | _GEN_26969; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27298 = _T_1530 ? _GEN_27290 : _GEN_26962; // @[sequencer-master.scala 168:32]
  wire  _GEN_27299 = _T_1530 ? _GEN_27291 : _GEN_26963; // @[sequencer-master.scala 168:32]
  wire  _GEN_27300 = _T_1530 ? _GEN_27292 : _GEN_26964; // @[sequencer-master.scala 168:32]
  wire  _GEN_27301 = _T_1530 ? _GEN_27293 : _GEN_26965; // @[sequencer-master.scala 168:32]
  wire  _GEN_27302 = _T_1530 ? _GEN_27294 : _GEN_26966; // @[sequencer-master.scala 168:32]
  wire  _GEN_27303 = _T_1530 ? _GEN_27295 : _GEN_26967; // @[sequencer-master.scala 168:32]
  wire  _GEN_27304 = _T_1530 ? _GEN_27296 : _GEN_26968; // @[sequencer-master.scala 168:32]
  wire  _GEN_27305 = _T_1530 ? _GEN_27297 : _GEN_26969; // @[sequencer-master.scala 168:32]
  wire  _GEN_27306 = _GEN_34121 | _GEN_26986; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27307 = _GEN_34122 | _GEN_26987; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27308 = _GEN_34123 | _GEN_26988; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27309 = _GEN_34124 | _GEN_26989; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27310 = _GEN_34125 | _GEN_26990; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27311 = _GEN_34126 | _GEN_26991; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27312 = _GEN_34127 | _GEN_26992; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27313 = _GEN_34128 | _GEN_26993; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27314 = _T_1552 ? _GEN_27306 : _GEN_26986; // @[sequencer-master.scala 168:32]
  wire  _GEN_27315 = _T_1552 ? _GEN_27307 : _GEN_26987; // @[sequencer-master.scala 168:32]
  wire  _GEN_27316 = _T_1552 ? _GEN_27308 : _GEN_26988; // @[sequencer-master.scala 168:32]
  wire  _GEN_27317 = _T_1552 ? _GEN_27309 : _GEN_26989; // @[sequencer-master.scala 168:32]
  wire  _GEN_27318 = _T_1552 ? _GEN_27310 : _GEN_26990; // @[sequencer-master.scala 168:32]
  wire  _GEN_27319 = _T_1552 ? _GEN_27311 : _GEN_26991; // @[sequencer-master.scala 168:32]
  wire  _GEN_27320 = _T_1552 ? _GEN_27312 : _GEN_26992; // @[sequencer-master.scala 168:32]
  wire  _GEN_27321 = _T_1552 ? _GEN_27313 : _GEN_26993; // @[sequencer-master.scala 168:32]
  wire  _GEN_27322 = _GEN_34121 | _GEN_27010; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27323 = _GEN_34122 | _GEN_27011; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27324 = _GEN_34123 | _GEN_27012; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27325 = _GEN_34124 | _GEN_27013; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27326 = _GEN_34125 | _GEN_27014; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27327 = _GEN_34126 | _GEN_27015; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27328 = _GEN_34127 | _GEN_27016; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27329 = _GEN_34128 | _GEN_27017; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27330 = _T_1574 ? _GEN_27322 : _GEN_27010; // @[sequencer-master.scala 168:32]
  wire  _GEN_27331 = _T_1574 ? _GEN_27323 : _GEN_27011; // @[sequencer-master.scala 168:32]
  wire  _GEN_27332 = _T_1574 ? _GEN_27324 : _GEN_27012; // @[sequencer-master.scala 168:32]
  wire  _GEN_27333 = _T_1574 ? _GEN_27325 : _GEN_27013; // @[sequencer-master.scala 168:32]
  wire  _GEN_27334 = _T_1574 ? _GEN_27326 : _GEN_27014; // @[sequencer-master.scala 168:32]
  wire  _GEN_27335 = _T_1574 ? _GEN_27327 : _GEN_27015; // @[sequencer-master.scala 168:32]
  wire  _GEN_27336 = _T_1574 ? _GEN_27328 : _GEN_27016; // @[sequencer-master.scala 168:32]
  wire  _GEN_27337 = _T_1574 ? _GEN_27329 : _GEN_27017; // @[sequencer-master.scala 168:32]
  wire  _GEN_27338 = _GEN_34121 | _GEN_27034; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27339 = _GEN_34122 | _GEN_27035; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27340 = _GEN_34123 | _GEN_27036; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27341 = _GEN_34124 | _GEN_27037; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27342 = _GEN_34125 | _GEN_27038; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27343 = _GEN_34126 | _GEN_27039; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27344 = _GEN_34127 | _GEN_27040; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27345 = _GEN_34128 | _GEN_27041; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27346 = _T_1596 ? _GEN_27338 : _GEN_27034; // @[sequencer-master.scala 168:32]
  wire  _GEN_27347 = _T_1596 ? _GEN_27339 : _GEN_27035; // @[sequencer-master.scala 168:32]
  wire  _GEN_27348 = _T_1596 ? _GEN_27340 : _GEN_27036; // @[sequencer-master.scala 168:32]
  wire  _GEN_27349 = _T_1596 ? _GEN_27341 : _GEN_27037; // @[sequencer-master.scala 168:32]
  wire  _GEN_27350 = _T_1596 ? _GEN_27342 : _GEN_27038; // @[sequencer-master.scala 168:32]
  wire  _GEN_27351 = _T_1596 ? _GEN_27343 : _GEN_27039; // @[sequencer-master.scala 168:32]
  wire  _GEN_27352 = _T_1596 ? _GEN_27344 : _GEN_27040; // @[sequencer-master.scala 168:32]
  wire  _GEN_27353 = _T_1596 ? _GEN_27345 : _GEN_27041; // @[sequencer-master.scala 168:32]
  wire  _GEN_27354 = 3'h0 == _T_1647 | (3'h0 == _T_1645 | (_GEN_32729 | _GEN_25856)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27355 = 3'h1 == _T_1647 | (3'h1 == _T_1645 | (_GEN_32730 | _GEN_25857)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27356 = 3'h2 == _T_1647 | (3'h2 == _T_1645 | (_GEN_32731 | _GEN_25858)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27357 = 3'h3 == _T_1647 | (3'h3 == _T_1645 | (_GEN_32732 | _GEN_25859)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27358 = 3'h4 == _T_1647 | (3'h4 == _T_1645 | (_GEN_32733 | _GEN_25860)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27359 = 3'h5 == _T_1647 | (3'h5 == _T_1645 | (_GEN_32734 | _GEN_25861)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27360 = 3'h6 == _T_1647 | (3'h6 == _T_1645 | (_GEN_32735 | _GEN_25862)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27361 = 3'h7 == _T_1647 | (3'h7 == _T_1645 | (_GEN_32736 | _GEN_25863)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_27370 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26802; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27371 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26803; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27372 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26804; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27373 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26805; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27374 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26806; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27375 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26807; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27376 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26808; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27377 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26809; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_27378 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26810; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27379 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26811; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27380 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26812; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27381 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26813; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27382 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26814; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27383 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26815; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27384 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26816; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27385 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26817; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_27386 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26818; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27387 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26819; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27388 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26820; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27389 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26821; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27390 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26822; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27391 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26823; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27392 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26824; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27393 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26825; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_27394 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26826; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27395 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26827; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27396 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26828; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27397 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26829; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27398 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26830; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27399 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26831; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27400 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26832; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27401 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26833; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_27402 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26834; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27403 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26835; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27404 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26836; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27405 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26837; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27406 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26838; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27407 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26839; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27408 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26840; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27409 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26841; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_27410 = _GEN_36426 | (_GEN_34121 | (_GEN_32729 | _GEN_25912)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27411 = _GEN_36427 | (_GEN_34122 | (_GEN_32730 | _GEN_25913)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27412 = _GEN_36428 | (_GEN_34123 | (_GEN_32731 | _GEN_25914)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27413 = _GEN_36429 | (_GEN_34124 | (_GEN_32732 | _GEN_25915)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27414 = _GEN_36430 | (_GEN_34125 | (_GEN_32733 | _GEN_25916)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27415 = _GEN_36431 | (_GEN_34126 | (_GEN_32734 | _GEN_25917)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27416 = _GEN_36432 | (_GEN_34127 | (_GEN_32735 | _GEN_25918)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27417 = _GEN_36433 | (_GEN_34128 | (_GEN_32736 | _GEN_25919)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_27418 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26850; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27419 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26851; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27420 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26852; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27421 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26853; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27422 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26854; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27423 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26855; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27424 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26856; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27425 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26857; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27426 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27106; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27427 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27107; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27428 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27108; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27429 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27109; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27430 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27110; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27431 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27111; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27432 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27112; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27433 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27113; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27434 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27234; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27435 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27235; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27436 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27236; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27437 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27237; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27438 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27238; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27439 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27239; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27440 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27240; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27441 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27241; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27442 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26874; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27443 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26875; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27444 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26876; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27445 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26877; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27446 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26878; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27447 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26879; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27448 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26880; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27449 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26881; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27450 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27122; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27451 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27123; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27452 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27124; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27453 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27125; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27454 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27126; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27455 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27127; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27456 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27128; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27457 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27129; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27458 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27250; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27459 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27251; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27460 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27252; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27461 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27253; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27462 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27254; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27463 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27255; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27464 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27256; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27465 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27257; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27466 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26898; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27467 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26899; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27468 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26900; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27469 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26901; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27470 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26902; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27471 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26903; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27472 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26904; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27473 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26905; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27474 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27138; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27475 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27139; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27476 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27140; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27477 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27141; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27478 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27142; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27479 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27143; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27480 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27144; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27481 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27145; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27482 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27266; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27483 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27267; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27484 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27268; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27485 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27269; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27486 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27270; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27487 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27271; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27488 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27272; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27489 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27273; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27490 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26922; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27491 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26923; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27492 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26924; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27493 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26925; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27494 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26926; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27495 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26927; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27496 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26928; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27497 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26929; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27498 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27154; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27499 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27155; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27500 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27156; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27501 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27157; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27502 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27158; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27503 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27159; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27504 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27160; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27505 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27161; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27506 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27282; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27507 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27283; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27508 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27284; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27509 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27285; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27510 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27286; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27511 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27287; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27512 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27288; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27513 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27289; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27514 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26946; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27515 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26947; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27516 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26948; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27517 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26949; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27518 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26950; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27519 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26951; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27520 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26952; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27521 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26953; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27522 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27170; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27523 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27171; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27524 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27172; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27525 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27173; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27526 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27174; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27527 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27175; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27528 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27176; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27529 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27177; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27530 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27298; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27531 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27299; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27532 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27300; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27533 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27301; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27534 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27302; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27535 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27303; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27536 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27304; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27537 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27305; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27538 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26970; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27539 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26971; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27540 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26972; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27541 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26973; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27542 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26974; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27543 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26975; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27544 = 3'h6 == _T_1647 ? 1'h0 : _GEN_26976; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27545 = 3'h7 == _T_1647 ? 1'h0 : _GEN_26977; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27546 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27186; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27547 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27187; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27548 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27188; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27549 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27189; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27550 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27190; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27551 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27191; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27552 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27192; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27553 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27193; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27554 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27314; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27555 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27315; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27556 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27316; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27557 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27317; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27558 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27318; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27559 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27319; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27560 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27320; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27561 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27321; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27562 = 3'h0 == _T_1647 ? 1'h0 : _GEN_26994; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27563 = 3'h1 == _T_1647 ? 1'h0 : _GEN_26995; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27564 = 3'h2 == _T_1647 ? 1'h0 : _GEN_26996; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27565 = 3'h3 == _T_1647 ? 1'h0 : _GEN_26997; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27566 = 3'h4 == _T_1647 ? 1'h0 : _GEN_26998; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27567 = 3'h5 == _T_1647 ? 1'h0 : _GEN_26999; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27568 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27000; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27569 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27001; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27570 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27202; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27571 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27203; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27572 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27204; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27573 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27205; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27574 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27206; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27575 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27207; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27576 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27208; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27577 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27209; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27578 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27330; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27579 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27331; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27580 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27332; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27581 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27333; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27582 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27334; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27583 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27335; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27584 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27336; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27585 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27337; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27586 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27018; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27587 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27019; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27588 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27020; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27589 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27021; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27590 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27022; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27591 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27023; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27592 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27024; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27593 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27025; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_27594 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27218; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27595 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27219; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27596 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27220; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27597 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27221; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27598 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27222; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27599 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27223; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27600 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27224; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27601 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27225; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_27602 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27346; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27603 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27347; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27604 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27348; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27605 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27349; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27606 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27350; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27607 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27351; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27608 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27352; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27609 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27353; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_27610 = 3'h0 == _T_1647 ? 1'h0 : _GEN_27042; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27611 = 3'h1 == _T_1647 ? 1'h0 : _GEN_27043; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27612 = 3'h2 == _T_1647 ? 1'h0 : _GEN_27044; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27613 = 3'h3 == _T_1647 ? 1'h0 : _GEN_27045; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27614 = 3'h4 == _T_1647 ? 1'h0 : _GEN_27046; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27615 = 3'h5 == _T_1647 ? 1'h0 : _GEN_27047; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27616 = 3'h6 == _T_1647 ? 1'h0 : _GEN_27048; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27617 = 3'h7 == _T_1647 ? 1'h0 : _GEN_27049; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_27626 = _GEN_36426 | _GEN_23918; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27627 = _GEN_36427 | _GEN_23919; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27628 = _GEN_36428 | _GEN_23920; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27629 = _GEN_36429 | _GEN_23921; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27630 = _GEN_36430 | _GEN_23922; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27631 = _GEN_36431 | _GEN_23923; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27632 = _GEN_36432 | _GEN_23924; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_27633 = _GEN_36433 | _GEN_23925; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_27634 = 3'h0 == _T_1647 ? io_op_bits_fn_union : _GEN_27066; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27635 = 3'h1 == _T_1647 ? io_op_bits_fn_union : _GEN_27067; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27636 = 3'h2 == _T_1647 ? io_op_bits_fn_union : _GEN_27068; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27637 = 3'h3 == _T_1647 ? io_op_bits_fn_union : _GEN_27069; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27638 = 3'h4 == _T_1647 ? io_op_bits_fn_union : _GEN_27070; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27639 = 3'h5 == _T_1647 ? io_op_bits_fn_union : _GEN_27071; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27640 = 3'h6 == _T_1647 ? io_op_bits_fn_union : _GEN_27072; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_27641 = 3'h7 == _T_1647 ? io_op_bits_fn_union : _GEN_27073; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire  _GEN_27650 = 3'h0 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27402; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27651 = 3'h1 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27403; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27652 = 3'h2 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27404; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27653 = 3'h3 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27405; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27654 = 3'h4 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27406; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27655 = 3'h5 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27407; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27656 = 3'h6 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27408; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire  _GEN_27657 = 3'h7 == _T_1647 ? io_op_bits_base_vd_valid : _GEN_27409; // @[sequencer-master.scala 363:24 sequencer-master.scala 363:24]
  wire [7:0] _GEN_27682 = 3'h0 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23958; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27683 = 3'h1 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23959; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27684 = 3'h2 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23960; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27685 = 3'h3 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23961; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27686 = 3'h4 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23962; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27687 = 3'h5 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23963; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27688 = 3'h6 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23964; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire [7:0] _GEN_27689 = 3'h7 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_23965; // @[sequencer-master.scala 364:41 sequencer-master.scala 364:41]
  wire  _GEN_27698 = io_op_bits_base_vd_valid ? _GEN_27650 : _GEN_27402; // @[sequencer-master.scala 362:41]
  wire  _GEN_27699 = io_op_bits_base_vd_valid ? _GEN_27651 : _GEN_27403; // @[sequencer-master.scala 362:41]
  wire  _GEN_27700 = io_op_bits_base_vd_valid ? _GEN_27652 : _GEN_27404; // @[sequencer-master.scala 362:41]
  wire  _GEN_27701 = io_op_bits_base_vd_valid ? _GEN_27653 : _GEN_27405; // @[sequencer-master.scala 362:41]
  wire  _GEN_27702 = io_op_bits_base_vd_valid ? _GEN_27654 : _GEN_27406; // @[sequencer-master.scala 362:41]
  wire  _GEN_27703 = io_op_bits_base_vd_valid ? _GEN_27655 : _GEN_27407; // @[sequencer-master.scala 362:41]
  wire  _GEN_27704 = io_op_bits_base_vd_valid ? _GEN_27656 : _GEN_27408; // @[sequencer-master.scala 362:41]
  wire  _GEN_27705 = io_op_bits_base_vd_valid ? _GEN_27657 : _GEN_27409; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27730 = io_op_bits_base_vd_valid ? _GEN_27682 : _GEN_23958; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27731 = io_op_bits_base_vd_valid ? _GEN_27683 : _GEN_23959; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27732 = io_op_bits_base_vd_valid ? _GEN_27684 : _GEN_23960; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27733 = io_op_bits_base_vd_valid ? _GEN_27685 : _GEN_23961; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27734 = io_op_bits_base_vd_valid ? _GEN_27686 : _GEN_23962; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27735 = io_op_bits_base_vd_valid ? _GEN_27687 : _GEN_23963; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27736 = io_op_bits_base_vd_valid ? _GEN_27688 : _GEN_23964; // @[sequencer-master.scala 362:41]
  wire [7:0] _GEN_27737 = io_op_bits_base_vd_valid ? _GEN_27689 : _GEN_23965; // @[sequencer-master.scala 362:41]
  wire  _GEN_27738 = _GEN_36426 | _GEN_27426; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27739 = _GEN_36427 | _GEN_27427; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27740 = _GEN_36428 | _GEN_27428; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27741 = _GEN_36429 | _GEN_27429; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27742 = _GEN_36430 | _GEN_27430; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27743 = _GEN_36431 | _GEN_27431; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27744 = _GEN_36432 | _GEN_27432; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27745 = _GEN_36433 | _GEN_27433; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27746 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27738 : _GEN_27426; // @[sequencer-master.scala 161:86]
  wire  _GEN_27747 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27739 : _GEN_27427; // @[sequencer-master.scala 161:86]
  wire  _GEN_27748 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27740 : _GEN_27428; // @[sequencer-master.scala 161:86]
  wire  _GEN_27749 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27741 : _GEN_27429; // @[sequencer-master.scala 161:86]
  wire  _GEN_27750 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27742 : _GEN_27430; // @[sequencer-master.scala 161:86]
  wire  _GEN_27751 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27743 : _GEN_27431; // @[sequencer-master.scala 161:86]
  wire  _GEN_27752 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27744 : _GEN_27432; // @[sequencer-master.scala 161:86]
  wire  _GEN_27753 = _T_734 | _T_911 | _T_1088 | _T_1265 ? _GEN_27745 : _GEN_27433; // @[sequencer-master.scala 161:86]
  wire  _GEN_27754 = _GEN_36426 | _GEN_27450; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27755 = _GEN_36427 | _GEN_27451; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27756 = _GEN_36428 | _GEN_27452; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27757 = _GEN_36429 | _GEN_27453; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27758 = _GEN_36430 | _GEN_27454; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27759 = _GEN_36431 | _GEN_27455; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27760 = _GEN_36432 | _GEN_27456; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27761 = _GEN_36433 | _GEN_27457; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27762 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27754 : _GEN_27450; // @[sequencer-master.scala 161:86]
  wire  _GEN_27763 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27755 : _GEN_27451; // @[sequencer-master.scala 161:86]
  wire  _GEN_27764 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27756 : _GEN_27452; // @[sequencer-master.scala 161:86]
  wire  _GEN_27765 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27757 : _GEN_27453; // @[sequencer-master.scala 161:86]
  wire  _GEN_27766 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27758 : _GEN_27454; // @[sequencer-master.scala 161:86]
  wire  _GEN_27767 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27759 : _GEN_27455; // @[sequencer-master.scala 161:86]
  wire  _GEN_27768 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27760 : _GEN_27456; // @[sequencer-master.scala 161:86]
  wire  _GEN_27769 = _T_756 | _T_933 | _T_1110 | _T_1287 ? _GEN_27761 : _GEN_27457; // @[sequencer-master.scala 161:86]
  wire  _GEN_27770 = _GEN_36426 | _GEN_27474; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27771 = _GEN_36427 | _GEN_27475; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27772 = _GEN_36428 | _GEN_27476; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27773 = _GEN_36429 | _GEN_27477; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27774 = _GEN_36430 | _GEN_27478; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27775 = _GEN_36431 | _GEN_27479; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27776 = _GEN_36432 | _GEN_27480; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27777 = _GEN_36433 | _GEN_27481; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27778 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27770 : _GEN_27474; // @[sequencer-master.scala 161:86]
  wire  _GEN_27779 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27771 : _GEN_27475; // @[sequencer-master.scala 161:86]
  wire  _GEN_27780 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27772 : _GEN_27476; // @[sequencer-master.scala 161:86]
  wire  _GEN_27781 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27773 : _GEN_27477; // @[sequencer-master.scala 161:86]
  wire  _GEN_27782 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27774 : _GEN_27478; // @[sequencer-master.scala 161:86]
  wire  _GEN_27783 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27775 : _GEN_27479; // @[sequencer-master.scala 161:86]
  wire  _GEN_27784 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27776 : _GEN_27480; // @[sequencer-master.scala 161:86]
  wire  _GEN_27785 = _T_778 | _T_955 | _T_1132 | _T_1309 ? _GEN_27777 : _GEN_27481; // @[sequencer-master.scala 161:86]
  wire  _GEN_27786 = _GEN_36426 | _GEN_27498; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27787 = _GEN_36427 | _GEN_27499; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27788 = _GEN_36428 | _GEN_27500; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27789 = _GEN_36429 | _GEN_27501; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27790 = _GEN_36430 | _GEN_27502; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27791 = _GEN_36431 | _GEN_27503; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27792 = _GEN_36432 | _GEN_27504; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27793 = _GEN_36433 | _GEN_27505; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27794 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27786 : _GEN_27498; // @[sequencer-master.scala 161:86]
  wire  _GEN_27795 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27787 : _GEN_27499; // @[sequencer-master.scala 161:86]
  wire  _GEN_27796 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27788 : _GEN_27500; // @[sequencer-master.scala 161:86]
  wire  _GEN_27797 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27789 : _GEN_27501; // @[sequencer-master.scala 161:86]
  wire  _GEN_27798 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27790 : _GEN_27502; // @[sequencer-master.scala 161:86]
  wire  _GEN_27799 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27791 : _GEN_27503; // @[sequencer-master.scala 161:86]
  wire  _GEN_27800 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27792 : _GEN_27504; // @[sequencer-master.scala 161:86]
  wire  _GEN_27801 = _T_800 | _T_977 | _T_1154 | _T_1331 ? _GEN_27793 : _GEN_27505; // @[sequencer-master.scala 161:86]
  wire  _GEN_27802 = _GEN_36426 | _GEN_27522; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27803 = _GEN_36427 | _GEN_27523; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27804 = _GEN_36428 | _GEN_27524; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27805 = _GEN_36429 | _GEN_27525; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27806 = _GEN_36430 | _GEN_27526; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27807 = _GEN_36431 | _GEN_27527; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27808 = _GEN_36432 | _GEN_27528; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27809 = _GEN_36433 | _GEN_27529; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27810 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27802 : _GEN_27522; // @[sequencer-master.scala 161:86]
  wire  _GEN_27811 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27803 : _GEN_27523; // @[sequencer-master.scala 161:86]
  wire  _GEN_27812 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27804 : _GEN_27524; // @[sequencer-master.scala 161:86]
  wire  _GEN_27813 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27805 : _GEN_27525; // @[sequencer-master.scala 161:86]
  wire  _GEN_27814 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27806 : _GEN_27526; // @[sequencer-master.scala 161:86]
  wire  _GEN_27815 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27807 : _GEN_27527; // @[sequencer-master.scala 161:86]
  wire  _GEN_27816 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27808 : _GEN_27528; // @[sequencer-master.scala 161:86]
  wire  _GEN_27817 = _T_822 | _T_999 | _T_1176 | _T_1353 ? _GEN_27809 : _GEN_27529; // @[sequencer-master.scala 161:86]
  wire  _GEN_27818 = _GEN_36426 | _GEN_27546; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27819 = _GEN_36427 | _GEN_27547; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27820 = _GEN_36428 | _GEN_27548; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27821 = _GEN_36429 | _GEN_27549; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27822 = _GEN_36430 | _GEN_27550; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27823 = _GEN_36431 | _GEN_27551; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27824 = _GEN_36432 | _GEN_27552; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27825 = _GEN_36433 | _GEN_27553; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27826 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27818 : _GEN_27546; // @[sequencer-master.scala 161:86]
  wire  _GEN_27827 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27819 : _GEN_27547; // @[sequencer-master.scala 161:86]
  wire  _GEN_27828 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27820 : _GEN_27548; // @[sequencer-master.scala 161:86]
  wire  _GEN_27829 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27821 : _GEN_27549; // @[sequencer-master.scala 161:86]
  wire  _GEN_27830 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27822 : _GEN_27550; // @[sequencer-master.scala 161:86]
  wire  _GEN_27831 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27823 : _GEN_27551; // @[sequencer-master.scala 161:86]
  wire  _GEN_27832 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27824 : _GEN_27552; // @[sequencer-master.scala 161:86]
  wire  _GEN_27833 = _T_844 | _T_1021 | _T_1198 | _T_1375 ? _GEN_27825 : _GEN_27553; // @[sequencer-master.scala 161:86]
  wire  _GEN_27834 = _GEN_36426 | _GEN_27570; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27835 = _GEN_36427 | _GEN_27571; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27836 = _GEN_36428 | _GEN_27572; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27837 = _GEN_36429 | _GEN_27573; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27838 = _GEN_36430 | _GEN_27574; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27839 = _GEN_36431 | _GEN_27575; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27840 = _GEN_36432 | _GEN_27576; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27841 = _GEN_36433 | _GEN_27577; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27842 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27834 : _GEN_27570; // @[sequencer-master.scala 161:86]
  wire  _GEN_27843 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27835 : _GEN_27571; // @[sequencer-master.scala 161:86]
  wire  _GEN_27844 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27836 : _GEN_27572; // @[sequencer-master.scala 161:86]
  wire  _GEN_27845 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27837 : _GEN_27573; // @[sequencer-master.scala 161:86]
  wire  _GEN_27846 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27838 : _GEN_27574; // @[sequencer-master.scala 161:86]
  wire  _GEN_27847 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27839 : _GEN_27575; // @[sequencer-master.scala 161:86]
  wire  _GEN_27848 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27840 : _GEN_27576; // @[sequencer-master.scala 161:86]
  wire  _GEN_27849 = _T_866 | _T_1043 | _T_1220 | _T_1397 ? _GEN_27841 : _GEN_27577; // @[sequencer-master.scala 161:86]
  wire  _GEN_27850 = _GEN_36426 | _GEN_27594; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27851 = _GEN_36427 | _GEN_27595; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27852 = _GEN_36428 | _GEN_27596; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27853 = _GEN_36429 | _GEN_27597; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27854 = _GEN_36430 | _GEN_27598; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27855 = _GEN_36431 | _GEN_27599; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27856 = _GEN_36432 | _GEN_27600; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27857 = _GEN_36433 | _GEN_27601; // @[sequencer-master.scala 132:52 sequencer-master.scala 132:52]
  wire  _GEN_27858 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27850 : _GEN_27594; // @[sequencer-master.scala 161:86]
  wire  _GEN_27859 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27851 : _GEN_27595; // @[sequencer-master.scala 161:86]
  wire  _GEN_27860 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27852 : _GEN_27596; // @[sequencer-master.scala 161:86]
  wire  _GEN_27861 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27853 : _GEN_27597; // @[sequencer-master.scala 161:86]
  wire  _GEN_27862 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27854 : _GEN_27598; // @[sequencer-master.scala 161:86]
  wire  _GEN_27863 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27855 : _GEN_27599; // @[sequencer-master.scala 161:86]
  wire  _GEN_27864 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27856 : _GEN_27600; // @[sequencer-master.scala 161:86]
  wire  _GEN_27865 = _T_888 | _T_1065 | _T_1242 | _T_1419 ? _GEN_27857 : _GEN_27601; // @[sequencer-master.scala 161:86]
  wire  _GEN_27866 = _GEN_36426 | _GEN_27434; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27867 = _GEN_36427 | _GEN_27435; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27868 = _GEN_36428 | _GEN_27436; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27869 = _GEN_36429 | _GEN_27437; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27870 = _GEN_36430 | _GEN_27438; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27871 = _GEN_36431 | _GEN_27439; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27872 = _GEN_36432 | _GEN_27440; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27873 = _GEN_36433 | _GEN_27441; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27874 = _T_1442 ? _GEN_27866 : _GEN_27434; // @[sequencer-master.scala 168:32]
  wire  _GEN_27875 = _T_1442 ? _GEN_27867 : _GEN_27435; // @[sequencer-master.scala 168:32]
  wire  _GEN_27876 = _T_1442 ? _GEN_27868 : _GEN_27436; // @[sequencer-master.scala 168:32]
  wire  _GEN_27877 = _T_1442 ? _GEN_27869 : _GEN_27437; // @[sequencer-master.scala 168:32]
  wire  _GEN_27878 = _T_1442 ? _GEN_27870 : _GEN_27438; // @[sequencer-master.scala 168:32]
  wire  _GEN_27879 = _T_1442 ? _GEN_27871 : _GEN_27439; // @[sequencer-master.scala 168:32]
  wire  _GEN_27880 = _T_1442 ? _GEN_27872 : _GEN_27440; // @[sequencer-master.scala 168:32]
  wire  _GEN_27881 = _T_1442 ? _GEN_27873 : _GEN_27441; // @[sequencer-master.scala 168:32]
  wire  _GEN_27882 = _GEN_36426 | _GEN_27458; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27883 = _GEN_36427 | _GEN_27459; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27884 = _GEN_36428 | _GEN_27460; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27885 = _GEN_36429 | _GEN_27461; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27886 = _GEN_36430 | _GEN_27462; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27887 = _GEN_36431 | _GEN_27463; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27888 = _GEN_36432 | _GEN_27464; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27889 = _GEN_36433 | _GEN_27465; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27890 = _T_1464 ? _GEN_27882 : _GEN_27458; // @[sequencer-master.scala 168:32]
  wire  _GEN_27891 = _T_1464 ? _GEN_27883 : _GEN_27459; // @[sequencer-master.scala 168:32]
  wire  _GEN_27892 = _T_1464 ? _GEN_27884 : _GEN_27460; // @[sequencer-master.scala 168:32]
  wire  _GEN_27893 = _T_1464 ? _GEN_27885 : _GEN_27461; // @[sequencer-master.scala 168:32]
  wire  _GEN_27894 = _T_1464 ? _GEN_27886 : _GEN_27462; // @[sequencer-master.scala 168:32]
  wire  _GEN_27895 = _T_1464 ? _GEN_27887 : _GEN_27463; // @[sequencer-master.scala 168:32]
  wire  _GEN_27896 = _T_1464 ? _GEN_27888 : _GEN_27464; // @[sequencer-master.scala 168:32]
  wire  _GEN_27897 = _T_1464 ? _GEN_27889 : _GEN_27465; // @[sequencer-master.scala 168:32]
  wire  _GEN_27898 = _GEN_36426 | _GEN_27482; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27899 = _GEN_36427 | _GEN_27483; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27900 = _GEN_36428 | _GEN_27484; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27901 = _GEN_36429 | _GEN_27485; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27902 = _GEN_36430 | _GEN_27486; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27903 = _GEN_36431 | _GEN_27487; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27904 = _GEN_36432 | _GEN_27488; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27905 = _GEN_36433 | _GEN_27489; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27906 = _T_1486 ? _GEN_27898 : _GEN_27482; // @[sequencer-master.scala 168:32]
  wire  _GEN_27907 = _T_1486 ? _GEN_27899 : _GEN_27483; // @[sequencer-master.scala 168:32]
  wire  _GEN_27908 = _T_1486 ? _GEN_27900 : _GEN_27484; // @[sequencer-master.scala 168:32]
  wire  _GEN_27909 = _T_1486 ? _GEN_27901 : _GEN_27485; // @[sequencer-master.scala 168:32]
  wire  _GEN_27910 = _T_1486 ? _GEN_27902 : _GEN_27486; // @[sequencer-master.scala 168:32]
  wire  _GEN_27911 = _T_1486 ? _GEN_27903 : _GEN_27487; // @[sequencer-master.scala 168:32]
  wire  _GEN_27912 = _T_1486 ? _GEN_27904 : _GEN_27488; // @[sequencer-master.scala 168:32]
  wire  _GEN_27913 = _T_1486 ? _GEN_27905 : _GEN_27489; // @[sequencer-master.scala 168:32]
  wire  _GEN_27914 = _GEN_36426 | _GEN_27506; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27915 = _GEN_36427 | _GEN_27507; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27916 = _GEN_36428 | _GEN_27508; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27917 = _GEN_36429 | _GEN_27509; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27918 = _GEN_36430 | _GEN_27510; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27919 = _GEN_36431 | _GEN_27511; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27920 = _GEN_36432 | _GEN_27512; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27921 = _GEN_36433 | _GEN_27513; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27922 = _T_1508 ? _GEN_27914 : _GEN_27506; // @[sequencer-master.scala 168:32]
  wire  _GEN_27923 = _T_1508 ? _GEN_27915 : _GEN_27507; // @[sequencer-master.scala 168:32]
  wire  _GEN_27924 = _T_1508 ? _GEN_27916 : _GEN_27508; // @[sequencer-master.scala 168:32]
  wire  _GEN_27925 = _T_1508 ? _GEN_27917 : _GEN_27509; // @[sequencer-master.scala 168:32]
  wire  _GEN_27926 = _T_1508 ? _GEN_27918 : _GEN_27510; // @[sequencer-master.scala 168:32]
  wire  _GEN_27927 = _T_1508 ? _GEN_27919 : _GEN_27511; // @[sequencer-master.scala 168:32]
  wire  _GEN_27928 = _T_1508 ? _GEN_27920 : _GEN_27512; // @[sequencer-master.scala 168:32]
  wire  _GEN_27929 = _T_1508 ? _GEN_27921 : _GEN_27513; // @[sequencer-master.scala 168:32]
  wire  _GEN_27930 = _GEN_36426 | _GEN_27530; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27931 = _GEN_36427 | _GEN_27531; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27932 = _GEN_36428 | _GEN_27532; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27933 = _GEN_36429 | _GEN_27533; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27934 = _GEN_36430 | _GEN_27534; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27935 = _GEN_36431 | _GEN_27535; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27936 = _GEN_36432 | _GEN_27536; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27937 = _GEN_36433 | _GEN_27537; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27938 = _T_1530 ? _GEN_27930 : _GEN_27530; // @[sequencer-master.scala 168:32]
  wire  _GEN_27939 = _T_1530 ? _GEN_27931 : _GEN_27531; // @[sequencer-master.scala 168:32]
  wire  _GEN_27940 = _T_1530 ? _GEN_27932 : _GEN_27532; // @[sequencer-master.scala 168:32]
  wire  _GEN_27941 = _T_1530 ? _GEN_27933 : _GEN_27533; // @[sequencer-master.scala 168:32]
  wire  _GEN_27942 = _T_1530 ? _GEN_27934 : _GEN_27534; // @[sequencer-master.scala 168:32]
  wire  _GEN_27943 = _T_1530 ? _GEN_27935 : _GEN_27535; // @[sequencer-master.scala 168:32]
  wire  _GEN_27944 = _T_1530 ? _GEN_27936 : _GEN_27536; // @[sequencer-master.scala 168:32]
  wire  _GEN_27945 = _T_1530 ? _GEN_27937 : _GEN_27537; // @[sequencer-master.scala 168:32]
  wire  _GEN_27946 = _GEN_36426 | _GEN_27554; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27947 = _GEN_36427 | _GEN_27555; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27948 = _GEN_36428 | _GEN_27556; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27949 = _GEN_36429 | _GEN_27557; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27950 = _GEN_36430 | _GEN_27558; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27951 = _GEN_36431 | _GEN_27559; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27952 = _GEN_36432 | _GEN_27560; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27953 = _GEN_36433 | _GEN_27561; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27954 = _T_1552 ? _GEN_27946 : _GEN_27554; // @[sequencer-master.scala 168:32]
  wire  _GEN_27955 = _T_1552 ? _GEN_27947 : _GEN_27555; // @[sequencer-master.scala 168:32]
  wire  _GEN_27956 = _T_1552 ? _GEN_27948 : _GEN_27556; // @[sequencer-master.scala 168:32]
  wire  _GEN_27957 = _T_1552 ? _GEN_27949 : _GEN_27557; // @[sequencer-master.scala 168:32]
  wire  _GEN_27958 = _T_1552 ? _GEN_27950 : _GEN_27558; // @[sequencer-master.scala 168:32]
  wire  _GEN_27959 = _T_1552 ? _GEN_27951 : _GEN_27559; // @[sequencer-master.scala 168:32]
  wire  _GEN_27960 = _T_1552 ? _GEN_27952 : _GEN_27560; // @[sequencer-master.scala 168:32]
  wire  _GEN_27961 = _T_1552 ? _GEN_27953 : _GEN_27561; // @[sequencer-master.scala 168:32]
  wire  _GEN_27962 = _GEN_36426 | _GEN_27578; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27963 = _GEN_36427 | _GEN_27579; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27964 = _GEN_36428 | _GEN_27580; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27965 = _GEN_36429 | _GEN_27581; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27966 = _GEN_36430 | _GEN_27582; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27967 = _GEN_36431 | _GEN_27583; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27968 = _GEN_36432 | _GEN_27584; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27969 = _GEN_36433 | _GEN_27585; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27970 = _T_1574 ? _GEN_27962 : _GEN_27578; // @[sequencer-master.scala 168:32]
  wire  _GEN_27971 = _T_1574 ? _GEN_27963 : _GEN_27579; // @[sequencer-master.scala 168:32]
  wire  _GEN_27972 = _T_1574 ? _GEN_27964 : _GEN_27580; // @[sequencer-master.scala 168:32]
  wire  _GEN_27973 = _T_1574 ? _GEN_27965 : _GEN_27581; // @[sequencer-master.scala 168:32]
  wire  _GEN_27974 = _T_1574 ? _GEN_27966 : _GEN_27582; // @[sequencer-master.scala 168:32]
  wire  _GEN_27975 = _T_1574 ? _GEN_27967 : _GEN_27583; // @[sequencer-master.scala 168:32]
  wire  _GEN_27976 = _T_1574 ? _GEN_27968 : _GEN_27584; // @[sequencer-master.scala 168:32]
  wire  _GEN_27977 = _T_1574 ? _GEN_27969 : _GEN_27585; // @[sequencer-master.scala 168:32]
  wire  _GEN_27978 = _GEN_36426 | _GEN_27602; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27979 = _GEN_36427 | _GEN_27603; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27980 = _GEN_36428 | _GEN_27604; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27981 = _GEN_36429 | _GEN_27605; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27982 = _GEN_36430 | _GEN_27606; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27983 = _GEN_36431 | _GEN_27607; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27984 = _GEN_36432 | _GEN_27608; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27985 = _GEN_36433 | _GEN_27609; // @[sequencer-master.scala 133:52 sequencer-master.scala 133:52]
  wire  _GEN_27986 = _T_1596 ? _GEN_27978 : _GEN_27602; // @[sequencer-master.scala 168:32]
  wire  _GEN_27987 = _T_1596 ? _GEN_27979 : _GEN_27603; // @[sequencer-master.scala 168:32]
  wire  _GEN_27988 = _T_1596 ? _GEN_27980 : _GEN_27604; // @[sequencer-master.scala 168:32]
  wire  _GEN_27989 = _T_1596 ? _GEN_27981 : _GEN_27605; // @[sequencer-master.scala 168:32]
  wire  _GEN_27990 = _T_1596 ? _GEN_27982 : _GEN_27606; // @[sequencer-master.scala 168:32]
  wire  _GEN_27991 = _T_1596 ? _GEN_27983 : _GEN_27607; // @[sequencer-master.scala 168:32]
  wire  _GEN_27992 = _T_1596 ? _GEN_27984 : _GEN_27608; // @[sequencer-master.scala 168:32]
  wire  _GEN_27993 = _T_1596 ? _GEN_27985 : _GEN_27609; // @[sequencer-master.scala 168:32]
  wire [1:0] _GEN_27994 = 3'h0 == _T_1647 ? 2'h0 : _GEN_27074; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27995 = 3'h1 == _T_1647 ? 2'h0 : _GEN_27075; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27996 = 3'h2 == _T_1647 ? 2'h0 : _GEN_27076; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27997 = 3'h3 == _T_1647 ? 2'h0 : _GEN_27077; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27998 = 3'h4 == _T_1647 ? 2'h0 : _GEN_27078; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_27999 = 3'h5 == _T_1647 ? 2'h0 : _GEN_27079; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28000 = 3'h6 == _T_1647 ? 2'h0 : _GEN_27080; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28001 = 3'h7 == _T_1647 ? 2'h0 : _GEN_27081; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_28002 = 3'h0 == _T_1647 ? 4'h0 : _GEN_27082; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28003 = 3'h1 == _T_1647 ? 4'h0 : _GEN_27083; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28004 = 3'h2 == _T_1647 ? 4'h0 : _GEN_27084; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28005 = 3'h3 == _T_1647 ? 4'h0 : _GEN_27085; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28006 = 3'h4 == _T_1647 ? 4'h0 : _GEN_27086; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28007 = 3'h5 == _T_1647 ? 4'h0 : _GEN_27087; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28008 = 3'h6 == _T_1647 ? 4'h0 : _GEN_27088; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28009 = 3'h7 == _T_1647 ? 4'h0 : _GEN_27089; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_28010 = 3'h0 == _T_1647 ? 3'h0 : _GEN_27090; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28011 = 3'h1 == _T_1647 ? 3'h0 : _GEN_27091; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28012 = 3'h2 == _T_1647 ? 3'h0 : _GEN_27092; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28013 = 3'h3 == _T_1647 ? 3'h0 : _GEN_27093; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28014 = 3'h4 == _T_1647 ? 3'h0 : _GEN_27094; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28015 = 3'h5 == _T_1647 ? 3'h0 : _GEN_27095; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28016 = 3'h6 == _T_1647 ? 3'h0 : _GEN_27096; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28017 = 3'h7 == _T_1647 ? 3'h0 : _GEN_27097; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_28018 = io_op_bits_active_vld ? _GEN_27354 : _GEN_25856; // @[sequencer-master.scala 653:38]
  wire  _GEN_28019 = io_op_bits_active_vld ? _GEN_27355 : _GEN_25857; // @[sequencer-master.scala 653:38]
  wire  _GEN_28020 = io_op_bits_active_vld ? _GEN_27356 : _GEN_25858; // @[sequencer-master.scala 653:38]
  wire  _GEN_28021 = io_op_bits_active_vld ? _GEN_27357 : _GEN_25859; // @[sequencer-master.scala 653:38]
  wire  _GEN_28022 = io_op_bits_active_vld ? _GEN_27358 : _GEN_25860; // @[sequencer-master.scala 653:38]
  wire  _GEN_28023 = io_op_bits_active_vld ? _GEN_27359 : _GEN_25861; // @[sequencer-master.scala 653:38]
  wire  _GEN_28024 = io_op_bits_active_vld ? _GEN_27360 : _GEN_25862; // @[sequencer-master.scala 653:38]
  wire  _GEN_28025 = io_op_bits_active_vld ? _GEN_27361 : _GEN_25863; // @[sequencer-master.scala 653:38]
  wire  _GEN_28034 = io_op_bits_active_vld ? _GEN_27370 : _GEN_25872; // @[sequencer-master.scala 653:38]
  wire  _GEN_28035 = io_op_bits_active_vld ? _GEN_27371 : _GEN_25873; // @[sequencer-master.scala 653:38]
  wire  _GEN_28036 = io_op_bits_active_vld ? _GEN_27372 : _GEN_25874; // @[sequencer-master.scala 653:38]
  wire  _GEN_28037 = io_op_bits_active_vld ? _GEN_27373 : _GEN_25875; // @[sequencer-master.scala 653:38]
  wire  _GEN_28038 = io_op_bits_active_vld ? _GEN_27374 : _GEN_25876; // @[sequencer-master.scala 653:38]
  wire  _GEN_28039 = io_op_bits_active_vld ? _GEN_27375 : _GEN_25877; // @[sequencer-master.scala 653:38]
  wire  _GEN_28040 = io_op_bits_active_vld ? _GEN_27376 : _GEN_25878; // @[sequencer-master.scala 653:38]
  wire  _GEN_28041 = io_op_bits_active_vld ? _GEN_27377 : _GEN_25879; // @[sequencer-master.scala 653:38]
  wire  _GEN_28042 = io_op_bits_active_vld ? _GEN_27378 : _GEN_25880; // @[sequencer-master.scala 653:38]
  wire  _GEN_28043 = io_op_bits_active_vld ? _GEN_27379 : _GEN_25881; // @[sequencer-master.scala 653:38]
  wire  _GEN_28044 = io_op_bits_active_vld ? _GEN_27380 : _GEN_25882; // @[sequencer-master.scala 653:38]
  wire  _GEN_28045 = io_op_bits_active_vld ? _GEN_27381 : _GEN_25883; // @[sequencer-master.scala 653:38]
  wire  _GEN_28046 = io_op_bits_active_vld ? _GEN_27382 : _GEN_25884; // @[sequencer-master.scala 653:38]
  wire  _GEN_28047 = io_op_bits_active_vld ? _GEN_27383 : _GEN_25885; // @[sequencer-master.scala 653:38]
  wire  _GEN_28048 = io_op_bits_active_vld ? _GEN_27384 : _GEN_25886; // @[sequencer-master.scala 653:38]
  wire  _GEN_28049 = io_op_bits_active_vld ? _GEN_27385 : _GEN_25887; // @[sequencer-master.scala 653:38]
  wire  _GEN_28050 = io_op_bits_active_vld ? _GEN_27386 : _GEN_25888; // @[sequencer-master.scala 653:38]
  wire  _GEN_28051 = io_op_bits_active_vld ? _GEN_27387 : _GEN_25889; // @[sequencer-master.scala 653:38]
  wire  _GEN_28052 = io_op_bits_active_vld ? _GEN_27388 : _GEN_25890; // @[sequencer-master.scala 653:38]
  wire  _GEN_28053 = io_op_bits_active_vld ? _GEN_27389 : _GEN_25891; // @[sequencer-master.scala 653:38]
  wire  _GEN_28054 = io_op_bits_active_vld ? _GEN_27390 : _GEN_25892; // @[sequencer-master.scala 653:38]
  wire  _GEN_28055 = io_op_bits_active_vld ? _GEN_27391 : _GEN_25893; // @[sequencer-master.scala 653:38]
  wire  _GEN_28056 = io_op_bits_active_vld ? _GEN_27392 : _GEN_25894; // @[sequencer-master.scala 653:38]
  wire  _GEN_28057 = io_op_bits_active_vld ? _GEN_27393 : _GEN_25895; // @[sequencer-master.scala 653:38]
  wire  _GEN_28058 = io_op_bits_active_vld ? _GEN_27394 : _GEN_25896; // @[sequencer-master.scala 653:38]
  wire  _GEN_28059 = io_op_bits_active_vld ? _GEN_27395 : _GEN_25897; // @[sequencer-master.scala 653:38]
  wire  _GEN_28060 = io_op_bits_active_vld ? _GEN_27396 : _GEN_25898; // @[sequencer-master.scala 653:38]
  wire  _GEN_28061 = io_op_bits_active_vld ? _GEN_27397 : _GEN_25899; // @[sequencer-master.scala 653:38]
  wire  _GEN_28062 = io_op_bits_active_vld ? _GEN_27398 : _GEN_25900; // @[sequencer-master.scala 653:38]
  wire  _GEN_28063 = io_op_bits_active_vld ? _GEN_27399 : _GEN_25901; // @[sequencer-master.scala 653:38]
  wire  _GEN_28064 = io_op_bits_active_vld ? _GEN_27400 : _GEN_25902; // @[sequencer-master.scala 653:38]
  wire  _GEN_28065 = io_op_bits_active_vld ? _GEN_27401 : _GEN_25903; // @[sequencer-master.scala 653:38]
  wire  _GEN_28066 = io_op_bits_active_vld ? _GEN_27698 : _GEN_25904; // @[sequencer-master.scala 653:38]
  wire  _GEN_28067 = io_op_bits_active_vld ? _GEN_27699 : _GEN_25905; // @[sequencer-master.scala 653:38]
  wire  _GEN_28068 = io_op_bits_active_vld ? _GEN_27700 : _GEN_25906; // @[sequencer-master.scala 653:38]
  wire  _GEN_28069 = io_op_bits_active_vld ? _GEN_27701 : _GEN_25907; // @[sequencer-master.scala 653:38]
  wire  _GEN_28070 = io_op_bits_active_vld ? _GEN_27702 : _GEN_25908; // @[sequencer-master.scala 653:38]
  wire  _GEN_28071 = io_op_bits_active_vld ? _GEN_27703 : _GEN_25909; // @[sequencer-master.scala 653:38]
  wire  _GEN_28072 = io_op_bits_active_vld ? _GEN_27704 : _GEN_25910; // @[sequencer-master.scala 653:38]
  wire  _GEN_28073 = io_op_bits_active_vld ? _GEN_27705 : _GEN_25911; // @[sequencer-master.scala 653:38]
  wire  _GEN_28074 = io_op_bits_active_vld ? _GEN_27410 : _GEN_25912; // @[sequencer-master.scala 653:38]
  wire  _GEN_28075 = io_op_bits_active_vld ? _GEN_27411 : _GEN_25913; // @[sequencer-master.scala 653:38]
  wire  _GEN_28076 = io_op_bits_active_vld ? _GEN_27412 : _GEN_25914; // @[sequencer-master.scala 653:38]
  wire  _GEN_28077 = io_op_bits_active_vld ? _GEN_27413 : _GEN_25915; // @[sequencer-master.scala 653:38]
  wire  _GEN_28078 = io_op_bits_active_vld ? _GEN_27414 : _GEN_25916; // @[sequencer-master.scala 653:38]
  wire  _GEN_28079 = io_op_bits_active_vld ? _GEN_27415 : _GEN_25917; // @[sequencer-master.scala 653:38]
  wire  _GEN_28080 = io_op_bits_active_vld ? _GEN_27416 : _GEN_25918; // @[sequencer-master.scala 653:38]
  wire  _GEN_28081 = io_op_bits_active_vld ? _GEN_27417 : _GEN_25919; // @[sequencer-master.scala 653:38]
  wire  _GEN_28082 = io_op_bits_active_vld ? _GEN_27418 : _GEN_25920; // @[sequencer-master.scala 653:38]
  wire  _GEN_28083 = io_op_bits_active_vld ? _GEN_27419 : _GEN_25921; // @[sequencer-master.scala 653:38]
  wire  _GEN_28084 = io_op_bits_active_vld ? _GEN_27420 : _GEN_25922; // @[sequencer-master.scala 653:38]
  wire  _GEN_28085 = io_op_bits_active_vld ? _GEN_27421 : _GEN_25923; // @[sequencer-master.scala 653:38]
  wire  _GEN_28086 = io_op_bits_active_vld ? _GEN_27422 : _GEN_25924; // @[sequencer-master.scala 653:38]
  wire  _GEN_28087 = io_op_bits_active_vld ? _GEN_27423 : _GEN_25925; // @[sequencer-master.scala 653:38]
  wire  _GEN_28088 = io_op_bits_active_vld ? _GEN_27424 : _GEN_25926; // @[sequencer-master.scala 653:38]
  wire  _GEN_28089 = io_op_bits_active_vld ? _GEN_27425 : _GEN_25927; // @[sequencer-master.scala 653:38]
  wire  _GEN_28090 = io_op_bits_active_vld ? _GEN_27746 : _GEN_25928; // @[sequencer-master.scala 653:38]
  wire  _GEN_28091 = io_op_bits_active_vld ? _GEN_27747 : _GEN_25929; // @[sequencer-master.scala 653:38]
  wire  _GEN_28092 = io_op_bits_active_vld ? _GEN_27748 : _GEN_25930; // @[sequencer-master.scala 653:38]
  wire  _GEN_28093 = io_op_bits_active_vld ? _GEN_27749 : _GEN_25931; // @[sequencer-master.scala 653:38]
  wire  _GEN_28094 = io_op_bits_active_vld ? _GEN_27750 : _GEN_25932; // @[sequencer-master.scala 653:38]
  wire  _GEN_28095 = io_op_bits_active_vld ? _GEN_27751 : _GEN_25933; // @[sequencer-master.scala 653:38]
  wire  _GEN_28096 = io_op_bits_active_vld ? _GEN_27752 : _GEN_25934; // @[sequencer-master.scala 653:38]
  wire  _GEN_28097 = io_op_bits_active_vld ? _GEN_27753 : _GEN_25935; // @[sequencer-master.scala 653:38]
  wire  _GEN_28098 = io_op_bits_active_vld ? _GEN_27874 : _GEN_25936; // @[sequencer-master.scala 653:38]
  wire  _GEN_28099 = io_op_bits_active_vld ? _GEN_27875 : _GEN_25937; // @[sequencer-master.scala 653:38]
  wire  _GEN_28100 = io_op_bits_active_vld ? _GEN_27876 : _GEN_25938; // @[sequencer-master.scala 653:38]
  wire  _GEN_28101 = io_op_bits_active_vld ? _GEN_27877 : _GEN_25939; // @[sequencer-master.scala 653:38]
  wire  _GEN_28102 = io_op_bits_active_vld ? _GEN_27878 : _GEN_25940; // @[sequencer-master.scala 653:38]
  wire  _GEN_28103 = io_op_bits_active_vld ? _GEN_27879 : _GEN_25941; // @[sequencer-master.scala 653:38]
  wire  _GEN_28104 = io_op_bits_active_vld ? _GEN_27880 : _GEN_25942; // @[sequencer-master.scala 653:38]
  wire  _GEN_28105 = io_op_bits_active_vld ? _GEN_27881 : _GEN_25943; // @[sequencer-master.scala 653:38]
  wire  _GEN_28106 = io_op_bits_active_vld ? _GEN_27442 : _GEN_25944; // @[sequencer-master.scala 653:38]
  wire  _GEN_28107 = io_op_bits_active_vld ? _GEN_27443 : _GEN_25945; // @[sequencer-master.scala 653:38]
  wire  _GEN_28108 = io_op_bits_active_vld ? _GEN_27444 : _GEN_25946; // @[sequencer-master.scala 653:38]
  wire  _GEN_28109 = io_op_bits_active_vld ? _GEN_27445 : _GEN_25947; // @[sequencer-master.scala 653:38]
  wire  _GEN_28110 = io_op_bits_active_vld ? _GEN_27446 : _GEN_25948; // @[sequencer-master.scala 653:38]
  wire  _GEN_28111 = io_op_bits_active_vld ? _GEN_27447 : _GEN_25949; // @[sequencer-master.scala 653:38]
  wire  _GEN_28112 = io_op_bits_active_vld ? _GEN_27448 : _GEN_25950; // @[sequencer-master.scala 653:38]
  wire  _GEN_28113 = io_op_bits_active_vld ? _GEN_27449 : _GEN_25951; // @[sequencer-master.scala 653:38]
  wire  _GEN_28114 = io_op_bits_active_vld ? _GEN_27762 : _GEN_25952; // @[sequencer-master.scala 653:38]
  wire  _GEN_28115 = io_op_bits_active_vld ? _GEN_27763 : _GEN_25953; // @[sequencer-master.scala 653:38]
  wire  _GEN_28116 = io_op_bits_active_vld ? _GEN_27764 : _GEN_25954; // @[sequencer-master.scala 653:38]
  wire  _GEN_28117 = io_op_bits_active_vld ? _GEN_27765 : _GEN_25955; // @[sequencer-master.scala 653:38]
  wire  _GEN_28118 = io_op_bits_active_vld ? _GEN_27766 : _GEN_25956; // @[sequencer-master.scala 653:38]
  wire  _GEN_28119 = io_op_bits_active_vld ? _GEN_27767 : _GEN_25957; // @[sequencer-master.scala 653:38]
  wire  _GEN_28120 = io_op_bits_active_vld ? _GEN_27768 : _GEN_25958; // @[sequencer-master.scala 653:38]
  wire  _GEN_28121 = io_op_bits_active_vld ? _GEN_27769 : _GEN_25959; // @[sequencer-master.scala 653:38]
  wire  _GEN_28122 = io_op_bits_active_vld ? _GEN_27890 : _GEN_25960; // @[sequencer-master.scala 653:38]
  wire  _GEN_28123 = io_op_bits_active_vld ? _GEN_27891 : _GEN_25961; // @[sequencer-master.scala 653:38]
  wire  _GEN_28124 = io_op_bits_active_vld ? _GEN_27892 : _GEN_25962; // @[sequencer-master.scala 653:38]
  wire  _GEN_28125 = io_op_bits_active_vld ? _GEN_27893 : _GEN_25963; // @[sequencer-master.scala 653:38]
  wire  _GEN_28126 = io_op_bits_active_vld ? _GEN_27894 : _GEN_25964; // @[sequencer-master.scala 653:38]
  wire  _GEN_28127 = io_op_bits_active_vld ? _GEN_27895 : _GEN_25965; // @[sequencer-master.scala 653:38]
  wire  _GEN_28128 = io_op_bits_active_vld ? _GEN_27896 : _GEN_25966; // @[sequencer-master.scala 653:38]
  wire  _GEN_28129 = io_op_bits_active_vld ? _GEN_27897 : _GEN_25967; // @[sequencer-master.scala 653:38]
  wire  _GEN_28130 = io_op_bits_active_vld ? _GEN_27466 : _GEN_25968; // @[sequencer-master.scala 653:38]
  wire  _GEN_28131 = io_op_bits_active_vld ? _GEN_27467 : _GEN_25969; // @[sequencer-master.scala 653:38]
  wire  _GEN_28132 = io_op_bits_active_vld ? _GEN_27468 : _GEN_25970; // @[sequencer-master.scala 653:38]
  wire  _GEN_28133 = io_op_bits_active_vld ? _GEN_27469 : _GEN_25971; // @[sequencer-master.scala 653:38]
  wire  _GEN_28134 = io_op_bits_active_vld ? _GEN_27470 : _GEN_25972; // @[sequencer-master.scala 653:38]
  wire  _GEN_28135 = io_op_bits_active_vld ? _GEN_27471 : _GEN_25973; // @[sequencer-master.scala 653:38]
  wire  _GEN_28136 = io_op_bits_active_vld ? _GEN_27472 : _GEN_25974; // @[sequencer-master.scala 653:38]
  wire  _GEN_28137 = io_op_bits_active_vld ? _GEN_27473 : _GEN_25975; // @[sequencer-master.scala 653:38]
  wire  _GEN_28138 = io_op_bits_active_vld ? _GEN_27778 : _GEN_25976; // @[sequencer-master.scala 653:38]
  wire  _GEN_28139 = io_op_bits_active_vld ? _GEN_27779 : _GEN_25977; // @[sequencer-master.scala 653:38]
  wire  _GEN_28140 = io_op_bits_active_vld ? _GEN_27780 : _GEN_25978; // @[sequencer-master.scala 653:38]
  wire  _GEN_28141 = io_op_bits_active_vld ? _GEN_27781 : _GEN_25979; // @[sequencer-master.scala 653:38]
  wire  _GEN_28142 = io_op_bits_active_vld ? _GEN_27782 : _GEN_25980; // @[sequencer-master.scala 653:38]
  wire  _GEN_28143 = io_op_bits_active_vld ? _GEN_27783 : _GEN_25981; // @[sequencer-master.scala 653:38]
  wire  _GEN_28144 = io_op_bits_active_vld ? _GEN_27784 : _GEN_25982; // @[sequencer-master.scala 653:38]
  wire  _GEN_28145 = io_op_bits_active_vld ? _GEN_27785 : _GEN_25983; // @[sequencer-master.scala 653:38]
  wire  _GEN_28146 = io_op_bits_active_vld ? _GEN_27906 : _GEN_25984; // @[sequencer-master.scala 653:38]
  wire  _GEN_28147 = io_op_bits_active_vld ? _GEN_27907 : _GEN_25985; // @[sequencer-master.scala 653:38]
  wire  _GEN_28148 = io_op_bits_active_vld ? _GEN_27908 : _GEN_25986; // @[sequencer-master.scala 653:38]
  wire  _GEN_28149 = io_op_bits_active_vld ? _GEN_27909 : _GEN_25987; // @[sequencer-master.scala 653:38]
  wire  _GEN_28150 = io_op_bits_active_vld ? _GEN_27910 : _GEN_25988; // @[sequencer-master.scala 653:38]
  wire  _GEN_28151 = io_op_bits_active_vld ? _GEN_27911 : _GEN_25989; // @[sequencer-master.scala 653:38]
  wire  _GEN_28152 = io_op_bits_active_vld ? _GEN_27912 : _GEN_25990; // @[sequencer-master.scala 653:38]
  wire  _GEN_28153 = io_op_bits_active_vld ? _GEN_27913 : _GEN_25991; // @[sequencer-master.scala 653:38]
  wire  _GEN_28154 = io_op_bits_active_vld ? _GEN_27490 : _GEN_25992; // @[sequencer-master.scala 653:38]
  wire  _GEN_28155 = io_op_bits_active_vld ? _GEN_27491 : _GEN_25993; // @[sequencer-master.scala 653:38]
  wire  _GEN_28156 = io_op_bits_active_vld ? _GEN_27492 : _GEN_25994; // @[sequencer-master.scala 653:38]
  wire  _GEN_28157 = io_op_bits_active_vld ? _GEN_27493 : _GEN_25995; // @[sequencer-master.scala 653:38]
  wire  _GEN_28158 = io_op_bits_active_vld ? _GEN_27494 : _GEN_25996; // @[sequencer-master.scala 653:38]
  wire  _GEN_28159 = io_op_bits_active_vld ? _GEN_27495 : _GEN_25997; // @[sequencer-master.scala 653:38]
  wire  _GEN_28160 = io_op_bits_active_vld ? _GEN_27496 : _GEN_25998; // @[sequencer-master.scala 653:38]
  wire  _GEN_28161 = io_op_bits_active_vld ? _GEN_27497 : _GEN_25999; // @[sequencer-master.scala 653:38]
  wire  _GEN_28162 = io_op_bits_active_vld ? _GEN_27794 : _GEN_26000; // @[sequencer-master.scala 653:38]
  wire  _GEN_28163 = io_op_bits_active_vld ? _GEN_27795 : _GEN_26001; // @[sequencer-master.scala 653:38]
  wire  _GEN_28164 = io_op_bits_active_vld ? _GEN_27796 : _GEN_26002; // @[sequencer-master.scala 653:38]
  wire  _GEN_28165 = io_op_bits_active_vld ? _GEN_27797 : _GEN_26003; // @[sequencer-master.scala 653:38]
  wire  _GEN_28166 = io_op_bits_active_vld ? _GEN_27798 : _GEN_26004; // @[sequencer-master.scala 653:38]
  wire  _GEN_28167 = io_op_bits_active_vld ? _GEN_27799 : _GEN_26005; // @[sequencer-master.scala 653:38]
  wire  _GEN_28168 = io_op_bits_active_vld ? _GEN_27800 : _GEN_26006; // @[sequencer-master.scala 653:38]
  wire  _GEN_28169 = io_op_bits_active_vld ? _GEN_27801 : _GEN_26007; // @[sequencer-master.scala 653:38]
  wire  _GEN_28170 = io_op_bits_active_vld ? _GEN_27922 : _GEN_26008; // @[sequencer-master.scala 653:38]
  wire  _GEN_28171 = io_op_bits_active_vld ? _GEN_27923 : _GEN_26009; // @[sequencer-master.scala 653:38]
  wire  _GEN_28172 = io_op_bits_active_vld ? _GEN_27924 : _GEN_26010; // @[sequencer-master.scala 653:38]
  wire  _GEN_28173 = io_op_bits_active_vld ? _GEN_27925 : _GEN_26011; // @[sequencer-master.scala 653:38]
  wire  _GEN_28174 = io_op_bits_active_vld ? _GEN_27926 : _GEN_26012; // @[sequencer-master.scala 653:38]
  wire  _GEN_28175 = io_op_bits_active_vld ? _GEN_27927 : _GEN_26013; // @[sequencer-master.scala 653:38]
  wire  _GEN_28176 = io_op_bits_active_vld ? _GEN_27928 : _GEN_26014; // @[sequencer-master.scala 653:38]
  wire  _GEN_28177 = io_op_bits_active_vld ? _GEN_27929 : _GEN_26015; // @[sequencer-master.scala 653:38]
  wire  _GEN_28178 = io_op_bits_active_vld ? _GEN_27514 : _GEN_26016; // @[sequencer-master.scala 653:38]
  wire  _GEN_28179 = io_op_bits_active_vld ? _GEN_27515 : _GEN_26017; // @[sequencer-master.scala 653:38]
  wire  _GEN_28180 = io_op_bits_active_vld ? _GEN_27516 : _GEN_26018; // @[sequencer-master.scala 653:38]
  wire  _GEN_28181 = io_op_bits_active_vld ? _GEN_27517 : _GEN_26019; // @[sequencer-master.scala 653:38]
  wire  _GEN_28182 = io_op_bits_active_vld ? _GEN_27518 : _GEN_26020; // @[sequencer-master.scala 653:38]
  wire  _GEN_28183 = io_op_bits_active_vld ? _GEN_27519 : _GEN_26021; // @[sequencer-master.scala 653:38]
  wire  _GEN_28184 = io_op_bits_active_vld ? _GEN_27520 : _GEN_26022; // @[sequencer-master.scala 653:38]
  wire  _GEN_28185 = io_op_bits_active_vld ? _GEN_27521 : _GEN_26023; // @[sequencer-master.scala 653:38]
  wire  _GEN_28186 = io_op_bits_active_vld ? _GEN_27810 : _GEN_26024; // @[sequencer-master.scala 653:38]
  wire  _GEN_28187 = io_op_bits_active_vld ? _GEN_27811 : _GEN_26025; // @[sequencer-master.scala 653:38]
  wire  _GEN_28188 = io_op_bits_active_vld ? _GEN_27812 : _GEN_26026; // @[sequencer-master.scala 653:38]
  wire  _GEN_28189 = io_op_bits_active_vld ? _GEN_27813 : _GEN_26027; // @[sequencer-master.scala 653:38]
  wire  _GEN_28190 = io_op_bits_active_vld ? _GEN_27814 : _GEN_26028; // @[sequencer-master.scala 653:38]
  wire  _GEN_28191 = io_op_bits_active_vld ? _GEN_27815 : _GEN_26029; // @[sequencer-master.scala 653:38]
  wire  _GEN_28192 = io_op_bits_active_vld ? _GEN_27816 : _GEN_26030; // @[sequencer-master.scala 653:38]
  wire  _GEN_28193 = io_op_bits_active_vld ? _GEN_27817 : _GEN_26031; // @[sequencer-master.scala 653:38]
  wire  _GEN_28194 = io_op_bits_active_vld ? _GEN_27938 : _GEN_26032; // @[sequencer-master.scala 653:38]
  wire  _GEN_28195 = io_op_bits_active_vld ? _GEN_27939 : _GEN_26033; // @[sequencer-master.scala 653:38]
  wire  _GEN_28196 = io_op_bits_active_vld ? _GEN_27940 : _GEN_26034; // @[sequencer-master.scala 653:38]
  wire  _GEN_28197 = io_op_bits_active_vld ? _GEN_27941 : _GEN_26035; // @[sequencer-master.scala 653:38]
  wire  _GEN_28198 = io_op_bits_active_vld ? _GEN_27942 : _GEN_26036; // @[sequencer-master.scala 653:38]
  wire  _GEN_28199 = io_op_bits_active_vld ? _GEN_27943 : _GEN_26037; // @[sequencer-master.scala 653:38]
  wire  _GEN_28200 = io_op_bits_active_vld ? _GEN_27944 : _GEN_26038; // @[sequencer-master.scala 653:38]
  wire  _GEN_28201 = io_op_bits_active_vld ? _GEN_27945 : _GEN_26039; // @[sequencer-master.scala 653:38]
  wire  _GEN_28202 = io_op_bits_active_vld ? _GEN_27538 : _GEN_26040; // @[sequencer-master.scala 653:38]
  wire  _GEN_28203 = io_op_bits_active_vld ? _GEN_27539 : _GEN_26041; // @[sequencer-master.scala 653:38]
  wire  _GEN_28204 = io_op_bits_active_vld ? _GEN_27540 : _GEN_26042; // @[sequencer-master.scala 653:38]
  wire  _GEN_28205 = io_op_bits_active_vld ? _GEN_27541 : _GEN_26043; // @[sequencer-master.scala 653:38]
  wire  _GEN_28206 = io_op_bits_active_vld ? _GEN_27542 : _GEN_26044; // @[sequencer-master.scala 653:38]
  wire  _GEN_28207 = io_op_bits_active_vld ? _GEN_27543 : _GEN_26045; // @[sequencer-master.scala 653:38]
  wire  _GEN_28208 = io_op_bits_active_vld ? _GEN_27544 : _GEN_26046; // @[sequencer-master.scala 653:38]
  wire  _GEN_28209 = io_op_bits_active_vld ? _GEN_27545 : _GEN_26047; // @[sequencer-master.scala 653:38]
  wire  _GEN_28210 = io_op_bits_active_vld ? _GEN_27826 : _GEN_26048; // @[sequencer-master.scala 653:38]
  wire  _GEN_28211 = io_op_bits_active_vld ? _GEN_27827 : _GEN_26049; // @[sequencer-master.scala 653:38]
  wire  _GEN_28212 = io_op_bits_active_vld ? _GEN_27828 : _GEN_26050; // @[sequencer-master.scala 653:38]
  wire  _GEN_28213 = io_op_bits_active_vld ? _GEN_27829 : _GEN_26051; // @[sequencer-master.scala 653:38]
  wire  _GEN_28214 = io_op_bits_active_vld ? _GEN_27830 : _GEN_26052; // @[sequencer-master.scala 653:38]
  wire  _GEN_28215 = io_op_bits_active_vld ? _GEN_27831 : _GEN_26053; // @[sequencer-master.scala 653:38]
  wire  _GEN_28216 = io_op_bits_active_vld ? _GEN_27832 : _GEN_26054; // @[sequencer-master.scala 653:38]
  wire  _GEN_28217 = io_op_bits_active_vld ? _GEN_27833 : _GEN_26055; // @[sequencer-master.scala 653:38]
  wire  _GEN_28218 = io_op_bits_active_vld ? _GEN_27954 : _GEN_26056; // @[sequencer-master.scala 653:38]
  wire  _GEN_28219 = io_op_bits_active_vld ? _GEN_27955 : _GEN_26057; // @[sequencer-master.scala 653:38]
  wire  _GEN_28220 = io_op_bits_active_vld ? _GEN_27956 : _GEN_26058; // @[sequencer-master.scala 653:38]
  wire  _GEN_28221 = io_op_bits_active_vld ? _GEN_27957 : _GEN_26059; // @[sequencer-master.scala 653:38]
  wire  _GEN_28222 = io_op_bits_active_vld ? _GEN_27958 : _GEN_26060; // @[sequencer-master.scala 653:38]
  wire  _GEN_28223 = io_op_bits_active_vld ? _GEN_27959 : _GEN_26061; // @[sequencer-master.scala 653:38]
  wire  _GEN_28224 = io_op_bits_active_vld ? _GEN_27960 : _GEN_26062; // @[sequencer-master.scala 653:38]
  wire  _GEN_28225 = io_op_bits_active_vld ? _GEN_27961 : _GEN_26063; // @[sequencer-master.scala 653:38]
  wire  _GEN_28226 = io_op_bits_active_vld ? _GEN_27562 : _GEN_26064; // @[sequencer-master.scala 653:38]
  wire  _GEN_28227 = io_op_bits_active_vld ? _GEN_27563 : _GEN_26065; // @[sequencer-master.scala 653:38]
  wire  _GEN_28228 = io_op_bits_active_vld ? _GEN_27564 : _GEN_26066; // @[sequencer-master.scala 653:38]
  wire  _GEN_28229 = io_op_bits_active_vld ? _GEN_27565 : _GEN_26067; // @[sequencer-master.scala 653:38]
  wire  _GEN_28230 = io_op_bits_active_vld ? _GEN_27566 : _GEN_26068; // @[sequencer-master.scala 653:38]
  wire  _GEN_28231 = io_op_bits_active_vld ? _GEN_27567 : _GEN_26069; // @[sequencer-master.scala 653:38]
  wire  _GEN_28232 = io_op_bits_active_vld ? _GEN_27568 : _GEN_26070; // @[sequencer-master.scala 653:38]
  wire  _GEN_28233 = io_op_bits_active_vld ? _GEN_27569 : _GEN_26071; // @[sequencer-master.scala 653:38]
  wire  _GEN_28234 = io_op_bits_active_vld ? _GEN_27842 : _GEN_26072; // @[sequencer-master.scala 653:38]
  wire  _GEN_28235 = io_op_bits_active_vld ? _GEN_27843 : _GEN_26073; // @[sequencer-master.scala 653:38]
  wire  _GEN_28236 = io_op_bits_active_vld ? _GEN_27844 : _GEN_26074; // @[sequencer-master.scala 653:38]
  wire  _GEN_28237 = io_op_bits_active_vld ? _GEN_27845 : _GEN_26075; // @[sequencer-master.scala 653:38]
  wire  _GEN_28238 = io_op_bits_active_vld ? _GEN_27846 : _GEN_26076; // @[sequencer-master.scala 653:38]
  wire  _GEN_28239 = io_op_bits_active_vld ? _GEN_27847 : _GEN_26077; // @[sequencer-master.scala 653:38]
  wire  _GEN_28240 = io_op_bits_active_vld ? _GEN_27848 : _GEN_26078; // @[sequencer-master.scala 653:38]
  wire  _GEN_28241 = io_op_bits_active_vld ? _GEN_27849 : _GEN_26079; // @[sequencer-master.scala 653:38]
  wire  _GEN_28242 = io_op_bits_active_vld ? _GEN_27970 : _GEN_26080; // @[sequencer-master.scala 653:38]
  wire  _GEN_28243 = io_op_bits_active_vld ? _GEN_27971 : _GEN_26081; // @[sequencer-master.scala 653:38]
  wire  _GEN_28244 = io_op_bits_active_vld ? _GEN_27972 : _GEN_26082; // @[sequencer-master.scala 653:38]
  wire  _GEN_28245 = io_op_bits_active_vld ? _GEN_27973 : _GEN_26083; // @[sequencer-master.scala 653:38]
  wire  _GEN_28246 = io_op_bits_active_vld ? _GEN_27974 : _GEN_26084; // @[sequencer-master.scala 653:38]
  wire  _GEN_28247 = io_op_bits_active_vld ? _GEN_27975 : _GEN_26085; // @[sequencer-master.scala 653:38]
  wire  _GEN_28248 = io_op_bits_active_vld ? _GEN_27976 : _GEN_26086; // @[sequencer-master.scala 653:38]
  wire  _GEN_28249 = io_op_bits_active_vld ? _GEN_27977 : _GEN_26087; // @[sequencer-master.scala 653:38]
  wire  _GEN_28250 = io_op_bits_active_vld ? _GEN_27586 : _GEN_26088; // @[sequencer-master.scala 653:38]
  wire  _GEN_28251 = io_op_bits_active_vld ? _GEN_27587 : _GEN_26089; // @[sequencer-master.scala 653:38]
  wire  _GEN_28252 = io_op_bits_active_vld ? _GEN_27588 : _GEN_26090; // @[sequencer-master.scala 653:38]
  wire  _GEN_28253 = io_op_bits_active_vld ? _GEN_27589 : _GEN_26091; // @[sequencer-master.scala 653:38]
  wire  _GEN_28254 = io_op_bits_active_vld ? _GEN_27590 : _GEN_26092; // @[sequencer-master.scala 653:38]
  wire  _GEN_28255 = io_op_bits_active_vld ? _GEN_27591 : _GEN_26093; // @[sequencer-master.scala 653:38]
  wire  _GEN_28256 = io_op_bits_active_vld ? _GEN_27592 : _GEN_26094; // @[sequencer-master.scala 653:38]
  wire  _GEN_28257 = io_op_bits_active_vld ? _GEN_27593 : _GEN_26095; // @[sequencer-master.scala 653:38]
  wire  _GEN_28258 = io_op_bits_active_vld ? _GEN_27858 : _GEN_26096; // @[sequencer-master.scala 653:38]
  wire  _GEN_28259 = io_op_bits_active_vld ? _GEN_27859 : _GEN_26097; // @[sequencer-master.scala 653:38]
  wire  _GEN_28260 = io_op_bits_active_vld ? _GEN_27860 : _GEN_26098; // @[sequencer-master.scala 653:38]
  wire  _GEN_28261 = io_op_bits_active_vld ? _GEN_27861 : _GEN_26099; // @[sequencer-master.scala 653:38]
  wire  _GEN_28262 = io_op_bits_active_vld ? _GEN_27862 : _GEN_26100; // @[sequencer-master.scala 653:38]
  wire  _GEN_28263 = io_op_bits_active_vld ? _GEN_27863 : _GEN_26101; // @[sequencer-master.scala 653:38]
  wire  _GEN_28264 = io_op_bits_active_vld ? _GEN_27864 : _GEN_26102; // @[sequencer-master.scala 653:38]
  wire  _GEN_28265 = io_op_bits_active_vld ? _GEN_27865 : _GEN_26103; // @[sequencer-master.scala 653:38]
  wire  _GEN_28266 = io_op_bits_active_vld ? _GEN_27986 : _GEN_26104; // @[sequencer-master.scala 653:38]
  wire  _GEN_28267 = io_op_bits_active_vld ? _GEN_27987 : _GEN_26105; // @[sequencer-master.scala 653:38]
  wire  _GEN_28268 = io_op_bits_active_vld ? _GEN_27988 : _GEN_26106; // @[sequencer-master.scala 653:38]
  wire  _GEN_28269 = io_op_bits_active_vld ? _GEN_27989 : _GEN_26107; // @[sequencer-master.scala 653:38]
  wire  _GEN_28270 = io_op_bits_active_vld ? _GEN_27990 : _GEN_26108; // @[sequencer-master.scala 653:38]
  wire  _GEN_28271 = io_op_bits_active_vld ? _GEN_27991 : _GEN_26109; // @[sequencer-master.scala 653:38]
  wire  _GEN_28272 = io_op_bits_active_vld ? _GEN_27992 : _GEN_26110; // @[sequencer-master.scala 653:38]
  wire  _GEN_28273 = io_op_bits_active_vld ? _GEN_27993 : _GEN_26111; // @[sequencer-master.scala 653:38]
  wire  _GEN_28274 = io_op_bits_active_vld ? _GEN_27610 : _GEN_26112; // @[sequencer-master.scala 653:38]
  wire  _GEN_28275 = io_op_bits_active_vld ? _GEN_27611 : _GEN_26113; // @[sequencer-master.scala 653:38]
  wire  _GEN_28276 = io_op_bits_active_vld ? _GEN_27612 : _GEN_26114; // @[sequencer-master.scala 653:38]
  wire  _GEN_28277 = io_op_bits_active_vld ? _GEN_27613 : _GEN_26115; // @[sequencer-master.scala 653:38]
  wire  _GEN_28278 = io_op_bits_active_vld ? _GEN_27614 : _GEN_26116; // @[sequencer-master.scala 653:38]
  wire  _GEN_28279 = io_op_bits_active_vld ? _GEN_27615 : _GEN_26117; // @[sequencer-master.scala 653:38]
  wire  _GEN_28280 = io_op_bits_active_vld ? _GEN_27616 : _GEN_26118; // @[sequencer-master.scala 653:38]
  wire  _GEN_28281 = io_op_bits_active_vld ? _GEN_27617 : _GEN_26119; // @[sequencer-master.scala 653:38]
  wire  _GEN_28290 = io_op_bits_active_vld ? _GEN_26538 : e_0_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28291 = io_op_bits_active_vld ? _GEN_26539 : e_1_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28292 = io_op_bits_active_vld ? _GEN_26540 : e_2_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28293 = io_op_bits_active_vld ? _GEN_26541 : e_3_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28294 = io_op_bits_active_vld ? _GEN_26542 : e_4_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28295 = io_op_bits_active_vld ? _GEN_26543 : e_5_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28296 = io_op_bits_active_vld ? _GEN_26544 : e_6_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire  _GEN_28297 = io_op_bits_active_vld ? _GEN_26545 : e_7_active_vpu; // @[sequencer-master.scala 653:38 sequencer-master.scala 109:14]
  wire [9:0] _GEN_28298 = io_op_bits_active_vld ? _GEN_27634 : _GEN_26136; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28299 = io_op_bits_active_vld ? _GEN_27635 : _GEN_26137; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28300 = io_op_bits_active_vld ? _GEN_27636 : _GEN_26138; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28301 = io_op_bits_active_vld ? _GEN_27637 : _GEN_26139; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28302 = io_op_bits_active_vld ? _GEN_27638 : _GEN_26140; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28303 = io_op_bits_active_vld ? _GEN_27639 : _GEN_26141; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28304 = io_op_bits_active_vld ? _GEN_27640 : _GEN_26142; // @[sequencer-master.scala 653:38]
  wire [9:0] _GEN_28305 = io_op_bits_active_vld ? _GEN_27641 : _GEN_26143; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28306 = io_op_bits_active_vld ? _GEN_26594 : _GEN_26144; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28307 = io_op_bits_active_vld ? _GEN_26595 : _GEN_26145; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28308 = io_op_bits_active_vld ? _GEN_26596 : _GEN_26146; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28309 = io_op_bits_active_vld ? _GEN_26597 : _GEN_26147; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28310 = io_op_bits_active_vld ? _GEN_26598 : _GEN_26148; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28311 = io_op_bits_active_vld ? _GEN_26599 : _GEN_26149; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28312 = io_op_bits_active_vld ? _GEN_26600 : _GEN_26150; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28313 = io_op_bits_active_vld ? _GEN_26601 : _GEN_26151; // @[sequencer-master.scala 653:38]
  wire  _GEN_28314 = io_op_bits_active_vld ? _GEN_26610 : _GEN_26152; // @[sequencer-master.scala 653:38]
  wire  _GEN_28315 = io_op_bits_active_vld ? _GEN_26611 : _GEN_26153; // @[sequencer-master.scala 653:38]
  wire  _GEN_28316 = io_op_bits_active_vld ? _GEN_26612 : _GEN_26154; // @[sequencer-master.scala 653:38]
  wire  _GEN_28317 = io_op_bits_active_vld ? _GEN_26613 : _GEN_26155; // @[sequencer-master.scala 653:38]
  wire  _GEN_28318 = io_op_bits_active_vld ? _GEN_26614 : _GEN_26156; // @[sequencer-master.scala 653:38]
  wire  _GEN_28319 = io_op_bits_active_vld ? _GEN_26615 : _GEN_26157; // @[sequencer-master.scala 653:38]
  wire  _GEN_28320 = io_op_bits_active_vld ? _GEN_26616 : _GEN_26158; // @[sequencer-master.scala 653:38]
  wire  _GEN_28321 = io_op_bits_active_vld ? _GEN_26617 : _GEN_26159; // @[sequencer-master.scala 653:38]
  wire  _GEN_28322 = io_op_bits_active_vld ? _GEN_26618 : _GEN_26160; // @[sequencer-master.scala 653:38]
  wire  _GEN_28323 = io_op_bits_active_vld ? _GEN_26619 : _GEN_26161; // @[sequencer-master.scala 653:38]
  wire  _GEN_28324 = io_op_bits_active_vld ? _GEN_26620 : _GEN_26162; // @[sequencer-master.scala 653:38]
  wire  _GEN_28325 = io_op_bits_active_vld ? _GEN_26621 : _GEN_26163; // @[sequencer-master.scala 653:38]
  wire  _GEN_28326 = io_op_bits_active_vld ? _GEN_26622 : _GEN_26164; // @[sequencer-master.scala 653:38]
  wire  _GEN_28327 = io_op_bits_active_vld ? _GEN_26623 : _GEN_26165; // @[sequencer-master.scala 653:38]
  wire  _GEN_28328 = io_op_bits_active_vld ? _GEN_26624 : _GEN_26166; // @[sequencer-master.scala 653:38]
  wire  _GEN_28329 = io_op_bits_active_vld ? _GEN_26625 : _GEN_26167; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28330 = io_op_bits_active_vld ? _GEN_26626 : _GEN_26168; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28331 = io_op_bits_active_vld ? _GEN_26627 : _GEN_26169; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28332 = io_op_bits_active_vld ? _GEN_26628 : _GEN_26170; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28333 = io_op_bits_active_vld ? _GEN_26629 : _GEN_26171; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28334 = io_op_bits_active_vld ? _GEN_26630 : _GEN_26172; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28335 = io_op_bits_active_vld ? _GEN_26631 : _GEN_26173; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28336 = io_op_bits_active_vld ? _GEN_26632 : _GEN_26174; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28337 = io_op_bits_active_vld ? _GEN_26633 : _GEN_26175; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28338 = io_op_bits_active_vld ? _GEN_27994 : _GEN_26224; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28339 = io_op_bits_active_vld ? _GEN_27995 : _GEN_26225; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28340 = io_op_bits_active_vld ? _GEN_27996 : _GEN_26226; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28341 = io_op_bits_active_vld ? _GEN_27997 : _GEN_26227; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28342 = io_op_bits_active_vld ? _GEN_27998 : _GEN_26228; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28343 = io_op_bits_active_vld ? _GEN_27999 : _GEN_26229; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28344 = io_op_bits_active_vld ? _GEN_28000 : _GEN_26230; // @[sequencer-master.scala 653:38]
  wire [1:0] _GEN_28345 = io_op_bits_active_vld ? _GEN_28001 : _GEN_26231; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28346 = io_op_bits_active_vld ? _GEN_28002 : _GEN_26232; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28347 = io_op_bits_active_vld ? _GEN_28003 : _GEN_26233; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28348 = io_op_bits_active_vld ? _GEN_28004 : _GEN_26234; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28349 = io_op_bits_active_vld ? _GEN_28005 : _GEN_26235; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28350 = io_op_bits_active_vld ? _GEN_28006 : _GEN_26236; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28351 = io_op_bits_active_vld ? _GEN_28007 : _GEN_26237; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28352 = io_op_bits_active_vld ? _GEN_28008 : _GEN_26238; // @[sequencer-master.scala 653:38]
  wire [3:0] _GEN_28353 = io_op_bits_active_vld ? _GEN_28009 : _GEN_26239; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28354 = io_op_bits_active_vld ? _GEN_28010 : _GEN_26240; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28355 = io_op_bits_active_vld ? _GEN_28011 : _GEN_26241; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28356 = io_op_bits_active_vld ? _GEN_28012 : _GEN_26242; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28357 = io_op_bits_active_vld ? _GEN_28013 : _GEN_26243; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28358 = io_op_bits_active_vld ? _GEN_28014 : _GEN_26244; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28359 = io_op_bits_active_vld ? _GEN_28015 : _GEN_26245; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28360 = io_op_bits_active_vld ? _GEN_28016 : _GEN_26246; // @[sequencer-master.scala 653:38]
  wire [2:0] _GEN_28361 = io_op_bits_active_vld ? _GEN_28017 : _GEN_26247; // @[sequencer-master.scala 653:38]
  wire  _GEN_28362 = io_op_bits_active_vld ? _GEN_27058 : _GEN_26248; // @[sequencer-master.scala 653:38]
  wire  _GEN_28363 = io_op_bits_active_vld ? _GEN_27059 : _GEN_26249; // @[sequencer-master.scala 653:38]
  wire  _GEN_28364 = io_op_bits_active_vld ? _GEN_27060 : _GEN_26250; // @[sequencer-master.scala 653:38]
  wire  _GEN_28365 = io_op_bits_active_vld ? _GEN_27061 : _GEN_26251; // @[sequencer-master.scala 653:38]
  wire  _GEN_28366 = io_op_bits_active_vld ? _GEN_27062 : _GEN_26252; // @[sequencer-master.scala 653:38]
  wire  _GEN_28367 = io_op_bits_active_vld ? _GEN_27063 : _GEN_26253; // @[sequencer-master.scala 653:38]
  wire  _GEN_28368 = io_op_bits_active_vld ? _GEN_27064 : _GEN_26254; // @[sequencer-master.scala 653:38]
  wire  _GEN_28369 = io_op_bits_active_vld ? _GEN_27065 : _GEN_26255; // @[sequencer-master.scala 653:38]
  wire  _GEN_28370 = io_op_bits_active_vld ? _GEN_27626 : _GEN_23918; // @[sequencer-master.scala 653:38]
  wire  _GEN_28371 = io_op_bits_active_vld ? _GEN_27627 : _GEN_23919; // @[sequencer-master.scala 653:38]
  wire  _GEN_28372 = io_op_bits_active_vld ? _GEN_27628 : _GEN_23920; // @[sequencer-master.scala 653:38]
  wire  _GEN_28373 = io_op_bits_active_vld ? _GEN_27629 : _GEN_23921; // @[sequencer-master.scala 653:38]
  wire  _GEN_28374 = io_op_bits_active_vld ? _GEN_27630 : _GEN_23922; // @[sequencer-master.scala 653:38]
  wire  _GEN_28375 = io_op_bits_active_vld ? _GEN_27631 : _GEN_23923; // @[sequencer-master.scala 653:38]
  wire  _GEN_28376 = io_op_bits_active_vld ? _GEN_27632 : _GEN_23924; // @[sequencer-master.scala 653:38]
  wire  _GEN_28377 = io_op_bits_active_vld ? _GEN_27633 : _GEN_23925; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28410 = io_op_bits_active_vld ? _GEN_27730 : _GEN_23958; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28411 = io_op_bits_active_vld ? _GEN_27731 : _GEN_23959; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28412 = io_op_bits_active_vld ? _GEN_27732 : _GEN_23960; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28413 = io_op_bits_active_vld ? _GEN_27733 : _GEN_23961; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28414 = io_op_bits_active_vld ? _GEN_27734 : _GEN_23962; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28415 = io_op_bits_active_vld ? _GEN_27735 : _GEN_23963; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28416 = io_op_bits_active_vld ? _GEN_27736 : _GEN_23964; // @[sequencer-master.scala 653:38]
  wire [7:0] _GEN_28417 = io_op_bits_active_vld ? _GEN_27737 : _GEN_23965; // @[sequencer-master.scala 653:38]
  wire  _GEN_28418 = io_op_bits_active_vld | _GEN_26264; // @[sequencer-master.scala 653:38 sequencer-master.scala 265:41]
  wire [2:0] _GEN_28419 = io_op_bits_active_vld ? _T_1649 : _GEN_26265; // @[sequencer-master.scala 653:38 sequencer-master.scala 265:66]
  wire  _GEN_28436 = 3'h0 == tail ? 1'h0 : _GEN_28034; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28437 = 3'h1 == tail ? 1'h0 : _GEN_28035; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28438 = 3'h2 == tail ? 1'h0 : _GEN_28036; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28439 = 3'h3 == tail ? 1'h0 : _GEN_28037; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28440 = 3'h4 == tail ? 1'h0 : _GEN_28038; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28441 = 3'h5 == tail ? 1'h0 : _GEN_28039; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28442 = 3'h6 == tail ? 1'h0 : _GEN_28040; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28443 = 3'h7 == tail ? 1'h0 : _GEN_28041; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28444 = 3'h0 == tail ? 1'h0 : _GEN_28042; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28445 = 3'h1 == tail ? 1'h0 : _GEN_28043; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28446 = 3'h2 == tail ? 1'h0 : _GEN_28044; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28447 = 3'h3 == tail ? 1'h0 : _GEN_28045; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28448 = 3'h4 == tail ? 1'h0 : _GEN_28046; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28449 = 3'h5 == tail ? 1'h0 : _GEN_28047; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28450 = 3'h6 == tail ? 1'h0 : _GEN_28048; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28451 = 3'h7 == tail ? 1'h0 : _GEN_28049; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28452 = 3'h0 == tail ? 1'h0 : _GEN_28050; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28453 = 3'h1 == tail ? 1'h0 : _GEN_28051; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28454 = 3'h2 == tail ? 1'h0 : _GEN_28052; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28455 = 3'h3 == tail ? 1'h0 : _GEN_28053; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28456 = 3'h4 == tail ? 1'h0 : _GEN_28054; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28457 = 3'h5 == tail ? 1'h0 : _GEN_28055; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28458 = 3'h6 == tail ? 1'h0 : _GEN_28056; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28459 = 3'h7 == tail ? 1'h0 : _GEN_28057; // @[sequencer-master.scala 274:29 sequencer-master.scala 274:29]
  wire  _GEN_28460 = 3'h0 == tail ? 1'h0 : _GEN_28058; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28461 = 3'h1 == tail ? 1'h0 : _GEN_28059; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28462 = 3'h2 == tail ? 1'h0 : _GEN_28060; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28463 = 3'h3 == tail ? 1'h0 : _GEN_28061; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28464 = 3'h4 == tail ? 1'h0 : _GEN_28062; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28465 = 3'h5 == tail ? 1'h0 : _GEN_28063; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28466 = 3'h6 == tail ? 1'h0 : _GEN_28064; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28467 = 3'h7 == tail ? 1'h0 : _GEN_28065; // @[sequencer-master.scala 275:29 sequencer-master.scala 275:29]
  wire  _GEN_28468 = 3'h0 == tail ? 1'h0 : _GEN_28066; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28469 = 3'h1 == tail ? 1'h0 : _GEN_28067; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28470 = 3'h2 == tail ? 1'h0 : _GEN_28068; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28471 = 3'h3 == tail ? 1'h0 : _GEN_28069; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28472 = 3'h4 == tail ? 1'h0 : _GEN_28070; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28473 = 3'h5 == tail ? 1'h0 : _GEN_28071; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28474 = 3'h6 == tail ? 1'h0 : _GEN_28072; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28475 = 3'h7 == tail ? 1'h0 : _GEN_28073; // @[sequencer-master.scala 276:28 sequencer-master.scala 276:28]
  wire  _GEN_28484 = 3'h0 == tail ? 1'h0 : _GEN_28082; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28485 = 3'h1 == tail ? 1'h0 : _GEN_28083; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28486 = 3'h2 == tail ? 1'h0 : _GEN_28084; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28487 = 3'h3 == tail ? 1'h0 : _GEN_28085; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28488 = 3'h4 == tail ? 1'h0 : _GEN_28086; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28489 = 3'h5 == tail ? 1'h0 : _GEN_28087; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28490 = 3'h6 == tail ? 1'h0 : _GEN_28088; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28491 = 3'h7 == tail ? 1'h0 : _GEN_28089; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28492 = 3'h0 == tail ? 1'h0 : _GEN_28090; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28493 = 3'h1 == tail ? 1'h0 : _GEN_28091; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28494 = 3'h2 == tail ? 1'h0 : _GEN_28092; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28495 = 3'h3 == tail ? 1'h0 : _GEN_28093; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28496 = 3'h4 == tail ? 1'h0 : _GEN_28094; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28497 = 3'h5 == tail ? 1'h0 : _GEN_28095; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28498 = 3'h6 == tail ? 1'h0 : _GEN_28096; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28499 = 3'h7 == tail ? 1'h0 : _GEN_28097; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28500 = 3'h0 == tail ? 1'h0 : _GEN_28098; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28501 = 3'h1 == tail ? 1'h0 : _GEN_28099; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28502 = 3'h2 == tail ? 1'h0 : _GEN_28100; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28503 = 3'h3 == tail ? 1'h0 : _GEN_28101; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28504 = 3'h4 == tail ? 1'h0 : _GEN_28102; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28505 = 3'h5 == tail ? 1'h0 : _GEN_28103; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28506 = 3'h6 == tail ? 1'h0 : _GEN_28104; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28507 = 3'h7 == tail ? 1'h0 : _GEN_28105; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28508 = 3'h0 == tail ? 1'h0 : _GEN_28106; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28509 = 3'h1 == tail ? 1'h0 : _GEN_28107; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28510 = 3'h2 == tail ? 1'h0 : _GEN_28108; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28511 = 3'h3 == tail ? 1'h0 : _GEN_28109; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28512 = 3'h4 == tail ? 1'h0 : _GEN_28110; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28513 = 3'h5 == tail ? 1'h0 : _GEN_28111; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28514 = 3'h6 == tail ? 1'h0 : _GEN_28112; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28515 = 3'h7 == tail ? 1'h0 : _GEN_28113; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28516 = 3'h0 == tail ? 1'h0 : _GEN_28114; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28517 = 3'h1 == tail ? 1'h0 : _GEN_28115; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28518 = 3'h2 == tail ? 1'h0 : _GEN_28116; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28519 = 3'h3 == tail ? 1'h0 : _GEN_28117; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28520 = 3'h4 == tail ? 1'h0 : _GEN_28118; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28521 = 3'h5 == tail ? 1'h0 : _GEN_28119; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28522 = 3'h6 == tail ? 1'h0 : _GEN_28120; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28523 = 3'h7 == tail ? 1'h0 : _GEN_28121; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28524 = 3'h0 == tail ? 1'h0 : _GEN_28122; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28525 = 3'h1 == tail ? 1'h0 : _GEN_28123; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28526 = 3'h2 == tail ? 1'h0 : _GEN_28124; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28527 = 3'h3 == tail ? 1'h0 : _GEN_28125; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28528 = 3'h4 == tail ? 1'h0 : _GEN_28126; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28529 = 3'h5 == tail ? 1'h0 : _GEN_28127; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28530 = 3'h6 == tail ? 1'h0 : _GEN_28128; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28531 = 3'h7 == tail ? 1'h0 : _GEN_28129; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28532 = 3'h0 == tail ? 1'h0 : _GEN_28130; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28533 = 3'h1 == tail ? 1'h0 : _GEN_28131; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28534 = 3'h2 == tail ? 1'h0 : _GEN_28132; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28535 = 3'h3 == tail ? 1'h0 : _GEN_28133; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28536 = 3'h4 == tail ? 1'h0 : _GEN_28134; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28537 = 3'h5 == tail ? 1'h0 : _GEN_28135; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28538 = 3'h6 == tail ? 1'h0 : _GEN_28136; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28539 = 3'h7 == tail ? 1'h0 : _GEN_28137; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28540 = 3'h0 == tail ? 1'h0 : _GEN_28138; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28541 = 3'h1 == tail ? 1'h0 : _GEN_28139; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28542 = 3'h2 == tail ? 1'h0 : _GEN_28140; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28543 = 3'h3 == tail ? 1'h0 : _GEN_28141; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28544 = 3'h4 == tail ? 1'h0 : _GEN_28142; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28545 = 3'h5 == tail ? 1'h0 : _GEN_28143; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28546 = 3'h6 == tail ? 1'h0 : _GEN_28144; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28547 = 3'h7 == tail ? 1'h0 : _GEN_28145; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28548 = 3'h0 == tail ? 1'h0 : _GEN_28146; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28549 = 3'h1 == tail ? 1'h0 : _GEN_28147; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28550 = 3'h2 == tail ? 1'h0 : _GEN_28148; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28551 = 3'h3 == tail ? 1'h0 : _GEN_28149; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28552 = 3'h4 == tail ? 1'h0 : _GEN_28150; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28553 = 3'h5 == tail ? 1'h0 : _GEN_28151; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28554 = 3'h6 == tail ? 1'h0 : _GEN_28152; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28555 = 3'h7 == tail ? 1'h0 : _GEN_28153; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28556 = 3'h0 == tail ? 1'h0 : _GEN_28154; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28557 = 3'h1 == tail ? 1'h0 : _GEN_28155; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28558 = 3'h2 == tail ? 1'h0 : _GEN_28156; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28559 = 3'h3 == tail ? 1'h0 : _GEN_28157; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28560 = 3'h4 == tail ? 1'h0 : _GEN_28158; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28561 = 3'h5 == tail ? 1'h0 : _GEN_28159; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28562 = 3'h6 == tail ? 1'h0 : _GEN_28160; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28563 = 3'h7 == tail ? 1'h0 : _GEN_28161; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28564 = 3'h0 == tail ? 1'h0 : _GEN_28162; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28565 = 3'h1 == tail ? 1'h0 : _GEN_28163; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28566 = 3'h2 == tail ? 1'h0 : _GEN_28164; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28567 = 3'h3 == tail ? 1'h0 : _GEN_28165; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28568 = 3'h4 == tail ? 1'h0 : _GEN_28166; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28569 = 3'h5 == tail ? 1'h0 : _GEN_28167; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28570 = 3'h6 == tail ? 1'h0 : _GEN_28168; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28571 = 3'h7 == tail ? 1'h0 : _GEN_28169; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28572 = 3'h0 == tail ? 1'h0 : _GEN_28170; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28573 = 3'h1 == tail ? 1'h0 : _GEN_28171; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28574 = 3'h2 == tail ? 1'h0 : _GEN_28172; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28575 = 3'h3 == tail ? 1'h0 : _GEN_28173; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28576 = 3'h4 == tail ? 1'h0 : _GEN_28174; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28577 = 3'h5 == tail ? 1'h0 : _GEN_28175; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28578 = 3'h6 == tail ? 1'h0 : _GEN_28176; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28579 = 3'h7 == tail ? 1'h0 : _GEN_28177; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28580 = 3'h0 == tail ? 1'h0 : _GEN_28178; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28581 = 3'h1 == tail ? 1'h0 : _GEN_28179; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28582 = 3'h2 == tail ? 1'h0 : _GEN_28180; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28583 = 3'h3 == tail ? 1'h0 : _GEN_28181; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28584 = 3'h4 == tail ? 1'h0 : _GEN_28182; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28585 = 3'h5 == tail ? 1'h0 : _GEN_28183; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28586 = 3'h6 == tail ? 1'h0 : _GEN_28184; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28587 = 3'h7 == tail ? 1'h0 : _GEN_28185; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28588 = 3'h0 == tail ? 1'h0 : _GEN_28186; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28589 = 3'h1 == tail ? 1'h0 : _GEN_28187; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28590 = 3'h2 == tail ? 1'h0 : _GEN_28188; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28591 = 3'h3 == tail ? 1'h0 : _GEN_28189; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28592 = 3'h4 == tail ? 1'h0 : _GEN_28190; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28593 = 3'h5 == tail ? 1'h0 : _GEN_28191; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28594 = 3'h6 == tail ? 1'h0 : _GEN_28192; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28595 = 3'h7 == tail ? 1'h0 : _GEN_28193; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28596 = 3'h0 == tail ? 1'h0 : _GEN_28194; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28597 = 3'h1 == tail ? 1'h0 : _GEN_28195; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28598 = 3'h2 == tail ? 1'h0 : _GEN_28196; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28599 = 3'h3 == tail ? 1'h0 : _GEN_28197; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28600 = 3'h4 == tail ? 1'h0 : _GEN_28198; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28601 = 3'h5 == tail ? 1'h0 : _GEN_28199; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28602 = 3'h6 == tail ? 1'h0 : _GEN_28200; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28603 = 3'h7 == tail ? 1'h0 : _GEN_28201; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28604 = 3'h0 == tail ? 1'h0 : _GEN_28202; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28605 = 3'h1 == tail ? 1'h0 : _GEN_28203; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28606 = 3'h2 == tail ? 1'h0 : _GEN_28204; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28607 = 3'h3 == tail ? 1'h0 : _GEN_28205; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28608 = 3'h4 == tail ? 1'h0 : _GEN_28206; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28609 = 3'h5 == tail ? 1'h0 : _GEN_28207; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28610 = 3'h6 == tail ? 1'h0 : _GEN_28208; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28611 = 3'h7 == tail ? 1'h0 : _GEN_28209; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28612 = 3'h0 == tail ? 1'h0 : _GEN_28210; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28613 = 3'h1 == tail ? 1'h0 : _GEN_28211; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28614 = 3'h2 == tail ? 1'h0 : _GEN_28212; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28615 = 3'h3 == tail ? 1'h0 : _GEN_28213; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28616 = 3'h4 == tail ? 1'h0 : _GEN_28214; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28617 = 3'h5 == tail ? 1'h0 : _GEN_28215; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28618 = 3'h6 == tail ? 1'h0 : _GEN_28216; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28619 = 3'h7 == tail ? 1'h0 : _GEN_28217; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28620 = 3'h0 == tail ? 1'h0 : _GEN_28218; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28621 = 3'h1 == tail ? 1'h0 : _GEN_28219; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28622 = 3'h2 == tail ? 1'h0 : _GEN_28220; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28623 = 3'h3 == tail ? 1'h0 : _GEN_28221; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28624 = 3'h4 == tail ? 1'h0 : _GEN_28222; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28625 = 3'h5 == tail ? 1'h0 : _GEN_28223; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28626 = 3'h6 == tail ? 1'h0 : _GEN_28224; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28627 = 3'h7 == tail ? 1'h0 : _GEN_28225; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28628 = 3'h0 == tail ? 1'h0 : _GEN_28226; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28629 = 3'h1 == tail ? 1'h0 : _GEN_28227; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28630 = 3'h2 == tail ? 1'h0 : _GEN_28228; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28631 = 3'h3 == tail ? 1'h0 : _GEN_28229; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28632 = 3'h4 == tail ? 1'h0 : _GEN_28230; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28633 = 3'h5 == tail ? 1'h0 : _GEN_28231; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28634 = 3'h6 == tail ? 1'h0 : _GEN_28232; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28635 = 3'h7 == tail ? 1'h0 : _GEN_28233; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28636 = 3'h0 == tail ? 1'h0 : _GEN_28234; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28637 = 3'h1 == tail ? 1'h0 : _GEN_28235; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28638 = 3'h2 == tail ? 1'h0 : _GEN_28236; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28639 = 3'h3 == tail ? 1'h0 : _GEN_28237; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28640 = 3'h4 == tail ? 1'h0 : _GEN_28238; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28641 = 3'h5 == tail ? 1'h0 : _GEN_28239; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28642 = 3'h6 == tail ? 1'h0 : _GEN_28240; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28643 = 3'h7 == tail ? 1'h0 : _GEN_28241; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28644 = 3'h0 == tail ? 1'h0 : _GEN_28242; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28645 = 3'h1 == tail ? 1'h0 : _GEN_28243; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28646 = 3'h2 == tail ? 1'h0 : _GEN_28244; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28647 = 3'h3 == tail ? 1'h0 : _GEN_28245; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28648 = 3'h4 == tail ? 1'h0 : _GEN_28246; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28649 = 3'h5 == tail ? 1'h0 : _GEN_28247; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28650 = 3'h6 == tail ? 1'h0 : _GEN_28248; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28651 = 3'h7 == tail ? 1'h0 : _GEN_28249; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28652 = 3'h0 == tail ? 1'h0 : _GEN_28250; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28653 = 3'h1 == tail ? 1'h0 : _GEN_28251; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28654 = 3'h2 == tail ? 1'h0 : _GEN_28252; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28655 = 3'h3 == tail ? 1'h0 : _GEN_28253; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28656 = 3'h4 == tail ? 1'h0 : _GEN_28254; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28657 = 3'h5 == tail ? 1'h0 : _GEN_28255; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28658 = 3'h6 == tail ? 1'h0 : _GEN_28256; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28659 = 3'h7 == tail ? 1'h0 : _GEN_28257; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_28660 = 3'h0 == tail ? 1'h0 : _GEN_28258; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28661 = 3'h1 == tail ? 1'h0 : _GEN_28259; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28662 = 3'h2 == tail ? 1'h0 : _GEN_28260; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28663 = 3'h3 == tail ? 1'h0 : _GEN_28261; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28664 = 3'h4 == tail ? 1'h0 : _GEN_28262; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28665 = 3'h5 == tail ? 1'h0 : _GEN_28263; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28666 = 3'h6 == tail ? 1'h0 : _GEN_28264; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28667 = 3'h7 == tail ? 1'h0 : _GEN_28265; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_28668 = 3'h0 == tail ? 1'h0 : _GEN_28266; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28669 = 3'h1 == tail ? 1'h0 : _GEN_28267; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28670 = 3'h2 == tail ? 1'h0 : _GEN_28268; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28671 = 3'h3 == tail ? 1'h0 : _GEN_28269; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28672 = 3'h4 == tail ? 1'h0 : _GEN_28270; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28673 = 3'h5 == tail ? 1'h0 : _GEN_28271; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28674 = 3'h6 == tail ? 1'h0 : _GEN_28272; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28675 = 3'h7 == tail ? 1'h0 : _GEN_28273; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_28676 = 3'h0 == tail ? 1'h0 : _GEN_28274; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28677 = 3'h1 == tail ? 1'h0 : _GEN_28275; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28678 = 3'h2 == tail ? 1'h0 : _GEN_28276; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28679 = 3'h3 == tail ? 1'h0 : _GEN_28277; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28680 = 3'h4 == tail ? 1'h0 : _GEN_28278; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28681 = 3'h5 == tail ? 1'h0 : _GEN_28279; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28682 = 3'h6 == tail ? 1'h0 : _GEN_28280; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28683 = 3'h7 == tail ? 1'h0 : _GEN_28281; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_28692 = _GEN_32729 | _GEN_28290; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28693 = _GEN_32730 | _GEN_28291; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28694 = _GEN_32731 | _GEN_28292; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28695 = _GEN_32732 | _GEN_28293; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28696 = _GEN_32733 | _GEN_28294; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28697 = _GEN_32734 | _GEN_28295; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28698 = _GEN_32735 | _GEN_28296; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_28699 = _GEN_32736 | _GEN_28297; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [9:0] _GEN_28700 = 3'h0 == tail ? io_op_bits_fn_union : _GEN_28298; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28701 = 3'h1 == tail ? io_op_bits_fn_union : _GEN_28299; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28702 = 3'h2 == tail ? io_op_bits_fn_union : _GEN_28300; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28703 = 3'h3 == tail ? io_op_bits_fn_union : _GEN_28301; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28704 = 3'h4 == tail ? io_op_bits_fn_union : _GEN_28302; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28705 = 3'h5 == tail ? io_op_bits_fn_union : _GEN_28303; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28706 = 3'h6 == tail ? io_op_bits_fn_union : _GEN_28304; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [9:0] _GEN_28707 = 3'h7 == tail ? io_op_bits_fn_union : _GEN_28305; // @[sequencer-master.scala 289:23 sequencer-master.scala 289:23]
  wire [3:0] _GEN_28708 = 3'h0 == tail ? io_op_bits_base_vp_id : _GEN_28306; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28709 = 3'h1 == tail ? io_op_bits_base_vp_id : _GEN_28307; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28710 = 3'h2 == tail ? io_op_bits_base_vp_id : _GEN_28308; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28711 = 3'h3 == tail ? io_op_bits_base_vp_id : _GEN_28309; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28712 = 3'h4 == tail ? io_op_bits_base_vp_id : _GEN_28310; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28713 = 3'h5 == tail ? io_op_bits_base_vp_id : _GEN_28311; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28714 = 3'h6 == tail ? io_op_bits_base_vp_id : _GEN_28312; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [3:0] _GEN_28715 = 3'h7 == tail ? io_op_bits_base_vp_id : _GEN_28313; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28716 = 3'h0 == tail ? io_op_bits_base_vp_valid : _GEN_28436; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28717 = 3'h1 == tail ? io_op_bits_base_vp_valid : _GEN_28437; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28718 = 3'h2 == tail ? io_op_bits_base_vp_valid : _GEN_28438; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28719 = 3'h3 == tail ? io_op_bits_base_vp_valid : _GEN_28439; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28720 = 3'h4 == tail ? io_op_bits_base_vp_valid : _GEN_28440; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28721 = 3'h5 == tail ? io_op_bits_base_vp_valid : _GEN_28441; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28722 = 3'h6 == tail ? io_op_bits_base_vp_valid : _GEN_28442; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28723 = 3'h7 == tail ? io_op_bits_base_vp_valid : _GEN_28443; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28724 = 3'h0 == tail ? io_op_bits_base_vp_scalar : _GEN_28314; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28725 = 3'h1 == tail ? io_op_bits_base_vp_scalar : _GEN_28315; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28726 = 3'h2 == tail ? io_op_bits_base_vp_scalar : _GEN_28316; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28727 = 3'h3 == tail ? io_op_bits_base_vp_scalar : _GEN_28317; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28728 = 3'h4 == tail ? io_op_bits_base_vp_scalar : _GEN_28318; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28729 = 3'h5 == tail ? io_op_bits_base_vp_scalar : _GEN_28319; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28730 = 3'h6 == tail ? io_op_bits_base_vp_scalar : _GEN_28320; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28731 = 3'h7 == tail ? io_op_bits_base_vp_scalar : _GEN_28321; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28732 = 3'h0 == tail ? io_op_bits_base_vp_pred : _GEN_28322; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28733 = 3'h1 == tail ? io_op_bits_base_vp_pred : _GEN_28323; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28734 = 3'h2 == tail ? io_op_bits_base_vp_pred : _GEN_28324; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28735 = 3'h3 == tail ? io_op_bits_base_vp_pred : _GEN_28325; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28736 = 3'h4 == tail ? io_op_bits_base_vp_pred : _GEN_28326; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28737 = 3'h5 == tail ? io_op_bits_base_vp_pred : _GEN_28327; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28738 = 3'h6 == tail ? io_op_bits_base_vp_pred : _GEN_28328; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire  _GEN_28739 = 3'h7 == tail ? io_op_bits_base_vp_pred : _GEN_28329; // @[sequencer-master.scala 321:24 sequencer-master.scala 321:24]
  wire [7:0] _GEN_28740 = 3'h0 == tail ? io_op_bits_reg_vp_id : _GEN_28330; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28741 = 3'h1 == tail ? io_op_bits_reg_vp_id : _GEN_28331; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28742 = 3'h2 == tail ? io_op_bits_reg_vp_id : _GEN_28332; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28743 = 3'h3 == tail ? io_op_bits_reg_vp_id : _GEN_28333; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28744 = 3'h4 == tail ? io_op_bits_reg_vp_id : _GEN_28334; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28745 = 3'h5 == tail ? io_op_bits_reg_vp_id : _GEN_28335; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28746 = 3'h6 == tail ? io_op_bits_reg_vp_id : _GEN_28336; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_28747 = 3'h7 == tail ? io_op_bits_reg_vp_id : _GEN_28337; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [3:0] _GEN_28748 = io_op_bits_base_vp_valid ? _GEN_28708 : _GEN_28306; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28749 = io_op_bits_base_vp_valid ? _GEN_28709 : _GEN_28307; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28750 = io_op_bits_base_vp_valid ? _GEN_28710 : _GEN_28308; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28751 = io_op_bits_base_vp_valid ? _GEN_28711 : _GEN_28309; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28752 = io_op_bits_base_vp_valid ? _GEN_28712 : _GEN_28310; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28753 = io_op_bits_base_vp_valid ? _GEN_28713 : _GEN_28311; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28754 = io_op_bits_base_vp_valid ? _GEN_28714 : _GEN_28312; // @[sequencer-master.scala 320:41]
  wire [3:0] _GEN_28755 = io_op_bits_base_vp_valid ? _GEN_28715 : _GEN_28313; // @[sequencer-master.scala 320:41]
  wire  _GEN_28756 = io_op_bits_base_vp_valid ? _GEN_28716 : _GEN_28436; // @[sequencer-master.scala 320:41]
  wire  _GEN_28757 = io_op_bits_base_vp_valid ? _GEN_28717 : _GEN_28437; // @[sequencer-master.scala 320:41]
  wire  _GEN_28758 = io_op_bits_base_vp_valid ? _GEN_28718 : _GEN_28438; // @[sequencer-master.scala 320:41]
  wire  _GEN_28759 = io_op_bits_base_vp_valid ? _GEN_28719 : _GEN_28439; // @[sequencer-master.scala 320:41]
  wire  _GEN_28760 = io_op_bits_base_vp_valid ? _GEN_28720 : _GEN_28440; // @[sequencer-master.scala 320:41]
  wire  _GEN_28761 = io_op_bits_base_vp_valid ? _GEN_28721 : _GEN_28441; // @[sequencer-master.scala 320:41]
  wire  _GEN_28762 = io_op_bits_base_vp_valid ? _GEN_28722 : _GEN_28442; // @[sequencer-master.scala 320:41]
  wire  _GEN_28763 = io_op_bits_base_vp_valid ? _GEN_28723 : _GEN_28443; // @[sequencer-master.scala 320:41]
  wire  _GEN_28764 = io_op_bits_base_vp_valid ? _GEN_28724 : _GEN_28314; // @[sequencer-master.scala 320:41]
  wire  _GEN_28765 = io_op_bits_base_vp_valid ? _GEN_28725 : _GEN_28315; // @[sequencer-master.scala 320:41]
  wire  _GEN_28766 = io_op_bits_base_vp_valid ? _GEN_28726 : _GEN_28316; // @[sequencer-master.scala 320:41]
  wire  _GEN_28767 = io_op_bits_base_vp_valid ? _GEN_28727 : _GEN_28317; // @[sequencer-master.scala 320:41]
  wire  _GEN_28768 = io_op_bits_base_vp_valid ? _GEN_28728 : _GEN_28318; // @[sequencer-master.scala 320:41]
  wire  _GEN_28769 = io_op_bits_base_vp_valid ? _GEN_28729 : _GEN_28319; // @[sequencer-master.scala 320:41]
  wire  _GEN_28770 = io_op_bits_base_vp_valid ? _GEN_28730 : _GEN_28320; // @[sequencer-master.scala 320:41]
  wire  _GEN_28771 = io_op_bits_base_vp_valid ? _GEN_28731 : _GEN_28321; // @[sequencer-master.scala 320:41]
  wire  _GEN_28772 = io_op_bits_base_vp_valid ? _GEN_28732 : _GEN_28322; // @[sequencer-master.scala 320:41]
  wire  _GEN_28773 = io_op_bits_base_vp_valid ? _GEN_28733 : _GEN_28323; // @[sequencer-master.scala 320:41]
  wire  _GEN_28774 = io_op_bits_base_vp_valid ? _GEN_28734 : _GEN_28324; // @[sequencer-master.scala 320:41]
  wire  _GEN_28775 = io_op_bits_base_vp_valid ? _GEN_28735 : _GEN_28325; // @[sequencer-master.scala 320:41]
  wire  _GEN_28776 = io_op_bits_base_vp_valid ? _GEN_28736 : _GEN_28326; // @[sequencer-master.scala 320:41]
  wire  _GEN_28777 = io_op_bits_base_vp_valid ? _GEN_28737 : _GEN_28327; // @[sequencer-master.scala 320:41]
  wire  _GEN_28778 = io_op_bits_base_vp_valid ? _GEN_28738 : _GEN_28328; // @[sequencer-master.scala 320:41]
  wire  _GEN_28779 = io_op_bits_base_vp_valid ? _GEN_28739 : _GEN_28329; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28780 = io_op_bits_base_vp_valid ? _GEN_28740 : _GEN_28330; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28781 = io_op_bits_base_vp_valid ? _GEN_28741 : _GEN_28331; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28782 = io_op_bits_base_vp_valid ? _GEN_28742 : _GEN_28332; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28783 = io_op_bits_base_vp_valid ? _GEN_28743 : _GEN_28333; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28784 = io_op_bits_base_vp_valid ? _GEN_28744 : _GEN_28334; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28785 = io_op_bits_base_vp_valid ? _GEN_28745 : _GEN_28335; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28786 = io_op_bits_base_vp_valid ? _GEN_28746 : _GEN_28336; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_28787 = io_op_bits_base_vp_valid ? _GEN_28747 : _GEN_28337; // @[sequencer-master.scala 320:41]
  wire  _GEN_28788 = _GEN_32729 | _GEN_28484; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28789 = _GEN_32730 | _GEN_28485; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28790 = _GEN_32731 | _GEN_28486; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28791 = _GEN_32732 | _GEN_28487; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28792 = _GEN_32733 | _GEN_28488; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28793 = _GEN_32734 | _GEN_28489; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28794 = _GEN_32735 | _GEN_28490; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28795 = _GEN_32736 | _GEN_28491; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28796 = _T_26 ? _GEN_28788 : _GEN_28484; // @[sequencer-master.scala 154:24]
  wire  _GEN_28797 = _T_26 ? _GEN_28789 : _GEN_28485; // @[sequencer-master.scala 154:24]
  wire  _GEN_28798 = _T_26 ? _GEN_28790 : _GEN_28486; // @[sequencer-master.scala 154:24]
  wire  _GEN_28799 = _T_26 ? _GEN_28791 : _GEN_28487; // @[sequencer-master.scala 154:24]
  wire  _GEN_28800 = _T_26 ? _GEN_28792 : _GEN_28488; // @[sequencer-master.scala 154:24]
  wire  _GEN_28801 = _T_26 ? _GEN_28793 : _GEN_28489; // @[sequencer-master.scala 154:24]
  wire  _GEN_28802 = _T_26 ? _GEN_28794 : _GEN_28490; // @[sequencer-master.scala 154:24]
  wire  _GEN_28803 = _T_26 ? _GEN_28795 : _GEN_28491; // @[sequencer-master.scala 154:24]
  wire  _GEN_28804 = _GEN_32729 | _GEN_28508; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28805 = _GEN_32730 | _GEN_28509; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28806 = _GEN_32731 | _GEN_28510; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28807 = _GEN_32732 | _GEN_28511; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28808 = _GEN_32733 | _GEN_28512; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28809 = _GEN_32734 | _GEN_28513; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28810 = _GEN_32735 | _GEN_28514; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28811 = _GEN_32736 | _GEN_28515; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28812 = _T_48 ? _GEN_28804 : _GEN_28508; // @[sequencer-master.scala 154:24]
  wire  _GEN_28813 = _T_48 ? _GEN_28805 : _GEN_28509; // @[sequencer-master.scala 154:24]
  wire  _GEN_28814 = _T_48 ? _GEN_28806 : _GEN_28510; // @[sequencer-master.scala 154:24]
  wire  _GEN_28815 = _T_48 ? _GEN_28807 : _GEN_28511; // @[sequencer-master.scala 154:24]
  wire  _GEN_28816 = _T_48 ? _GEN_28808 : _GEN_28512; // @[sequencer-master.scala 154:24]
  wire  _GEN_28817 = _T_48 ? _GEN_28809 : _GEN_28513; // @[sequencer-master.scala 154:24]
  wire  _GEN_28818 = _T_48 ? _GEN_28810 : _GEN_28514; // @[sequencer-master.scala 154:24]
  wire  _GEN_28819 = _T_48 ? _GEN_28811 : _GEN_28515; // @[sequencer-master.scala 154:24]
  wire  _GEN_28820 = _GEN_32729 | _GEN_28532; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28821 = _GEN_32730 | _GEN_28533; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28822 = _GEN_32731 | _GEN_28534; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28823 = _GEN_32732 | _GEN_28535; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28824 = _GEN_32733 | _GEN_28536; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28825 = _GEN_32734 | _GEN_28537; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28826 = _GEN_32735 | _GEN_28538; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28827 = _GEN_32736 | _GEN_28539; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28828 = _T_70 ? _GEN_28820 : _GEN_28532; // @[sequencer-master.scala 154:24]
  wire  _GEN_28829 = _T_70 ? _GEN_28821 : _GEN_28533; // @[sequencer-master.scala 154:24]
  wire  _GEN_28830 = _T_70 ? _GEN_28822 : _GEN_28534; // @[sequencer-master.scala 154:24]
  wire  _GEN_28831 = _T_70 ? _GEN_28823 : _GEN_28535; // @[sequencer-master.scala 154:24]
  wire  _GEN_28832 = _T_70 ? _GEN_28824 : _GEN_28536; // @[sequencer-master.scala 154:24]
  wire  _GEN_28833 = _T_70 ? _GEN_28825 : _GEN_28537; // @[sequencer-master.scala 154:24]
  wire  _GEN_28834 = _T_70 ? _GEN_28826 : _GEN_28538; // @[sequencer-master.scala 154:24]
  wire  _GEN_28835 = _T_70 ? _GEN_28827 : _GEN_28539; // @[sequencer-master.scala 154:24]
  wire  _GEN_28836 = _GEN_32729 | _GEN_28556; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28837 = _GEN_32730 | _GEN_28557; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28838 = _GEN_32731 | _GEN_28558; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28839 = _GEN_32732 | _GEN_28559; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28840 = _GEN_32733 | _GEN_28560; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28841 = _GEN_32734 | _GEN_28561; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28842 = _GEN_32735 | _GEN_28562; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28843 = _GEN_32736 | _GEN_28563; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28844 = _T_92 ? _GEN_28836 : _GEN_28556; // @[sequencer-master.scala 154:24]
  wire  _GEN_28845 = _T_92 ? _GEN_28837 : _GEN_28557; // @[sequencer-master.scala 154:24]
  wire  _GEN_28846 = _T_92 ? _GEN_28838 : _GEN_28558; // @[sequencer-master.scala 154:24]
  wire  _GEN_28847 = _T_92 ? _GEN_28839 : _GEN_28559; // @[sequencer-master.scala 154:24]
  wire  _GEN_28848 = _T_92 ? _GEN_28840 : _GEN_28560; // @[sequencer-master.scala 154:24]
  wire  _GEN_28849 = _T_92 ? _GEN_28841 : _GEN_28561; // @[sequencer-master.scala 154:24]
  wire  _GEN_28850 = _T_92 ? _GEN_28842 : _GEN_28562; // @[sequencer-master.scala 154:24]
  wire  _GEN_28851 = _T_92 ? _GEN_28843 : _GEN_28563; // @[sequencer-master.scala 154:24]
  wire  _GEN_28852 = _GEN_32729 | _GEN_28580; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28853 = _GEN_32730 | _GEN_28581; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28854 = _GEN_32731 | _GEN_28582; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28855 = _GEN_32732 | _GEN_28583; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28856 = _GEN_32733 | _GEN_28584; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28857 = _GEN_32734 | _GEN_28585; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28858 = _GEN_32735 | _GEN_28586; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28859 = _GEN_32736 | _GEN_28587; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28860 = _T_114 ? _GEN_28852 : _GEN_28580; // @[sequencer-master.scala 154:24]
  wire  _GEN_28861 = _T_114 ? _GEN_28853 : _GEN_28581; // @[sequencer-master.scala 154:24]
  wire  _GEN_28862 = _T_114 ? _GEN_28854 : _GEN_28582; // @[sequencer-master.scala 154:24]
  wire  _GEN_28863 = _T_114 ? _GEN_28855 : _GEN_28583; // @[sequencer-master.scala 154:24]
  wire  _GEN_28864 = _T_114 ? _GEN_28856 : _GEN_28584; // @[sequencer-master.scala 154:24]
  wire  _GEN_28865 = _T_114 ? _GEN_28857 : _GEN_28585; // @[sequencer-master.scala 154:24]
  wire  _GEN_28866 = _T_114 ? _GEN_28858 : _GEN_28586; // @[sequencer-master.scala 154:24]
  wire  _GEN_28867 = _T_114 ? _GEN_28859 : _GEN_28587; // @[sequencer-master.scala 154:24]
  wire  _GEN_28868 = _GEN_32729 | _GEN_28604; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28869 = _GEN_32730 | _GEN_28605; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28870 = _GEN_32731 | _GEN_28606; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28871 = _GEN_32732 | _GEN_28607; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28872 = _GEN_32733 | _GEN_28608; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28873 = _GEN_32734 | _GEN_28609; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28874 = _GEN_32735 | _GEN_28610; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28875 = _GEN_32736 | _GEN_28611; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28876 = _T_136 ? _GEN_28868 : _GEN_28604; // @[sequencer-master.scala 154:24]
  wire  _GEN_28877 = _T_136 ? _GEN_28869 : _GEN_28605; // @[sequencer-master.scala 154:24]
  wire  _GEN_28878 = _T_136 ? _GEN_28870 : _GEN_28606; // @[sequencer-master.scala 154:24]
  wire  _GEN_28879 = _T_136 ? _GEN_28871 : _GEN_28607; // @[sequencer-master.scala 154:24]
  wire  _GEN_28880 = _T_136 ? _GEN_28872 : _GEN_28608; // @[sequencer-master.scala 154:24]
  wire  _GEN_28881 = _T_136 ? _GEN_28873 : _GEN_28609; // @[sequencer-master.scala 154:24]
  wire  _GEN_28882 = _T_136 ? _GEN_28874 : _GEN_28610; // @[sequencer-master.scala 154:24]
  wire  _GEN_28883 = _T_136 ? _GEN_28875 : _GEN_28611; // @[sequencer-master.scala 154:24]
  wire  _GEN_28884 = _GEN_32729 | _GEN_28628; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28885 = _GEN_32730 | _GEN_28629; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28886 = _GEN_32731 | _GEN_28630; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28887 = _GEN_32732 | _GEN_28631; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28888 = _GEN_32733 | _GEN_28632; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28889 = _GEN_32734 | _GEN_28633; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28890 = _GEN_32735 | _GEN_28634; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28891 = _GEN_32736 | _GEN_28635; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28892 = _T_158 ? _GEN_28884 : _GEN_28628; // @[sequencer-master.scala 154:24]
  wire  _GEN_28893 = _T_158 ? _GEN_28885 : _GEN_28629; // @[sequencer-master.scala 154:24]
  wire  _GEN_28894 = _T_158 ? _GEN_28886 : _GEN_28630; // @[sequencer-master.scala 154:24]
  wire  _GEN_28895 = _T_158 ? _GEN_28887 : _GEN_28631; // @[sequencer-master.scala 154:24]
  wire  _GEN_28896 = _T_158 ? _GEN_28888 : _GEN_28632; // @[sequencer-master.scala 154:24]
  wire  _GEN_28897 = _T_158 ? _GEN_28889 : _GEN_28633; // @[sequencer-master.scala 154:24]
  wire  _GEN_28898 = _T_158 ? _GEN_28890 : _GEN_28634; // @[sequencer-master.scala 154:24]
  wire  _GEN_28899 = _T_158 ? _GEN_28891 : _GEN_28635; // @[sequencer-master.scala 154:24]
  wire  _GEN_28900 = _GEN_32729 | _GEN_28652; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28901 = _GEN_32730 | _GEN_28653; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28902 = _GEN_32731 | _GEN_28654; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28903 = _GEN_32732 | _GEN_28655; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28904 = _GEN_32733 | _GEN_28656; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28905 = _GEN_32734 | _GEN_28657; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28906 = _GEN_32735 | _GEN_28658; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28907 = _GEN_32736 | _GEN_28659; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_28908 = _T_180 ? _GEN_28900 : _GEN_28652; // @[sequencer-master.scala 154:24]
  wire  _GEN_28909 = _T_180 ? _GEN_28901 : _GEN_28653; // @[sequencer-master.scala 154:24]
  wire  _GEN_28910 = _T_180 ? _GEN_28902 : _GEN_28654; // @[sequencer-master.scala 154:24]
  wire  _GEN_28911 = _T_180 ? _GEN_28903 : _GEN_28655; // @[sequencer-master.scala 154:24]
  wire  _GEN_28912 = _T_180 ? _GEN_28904 : _GEN_28656; // @[sequencer-master.scala 154:24]
  wire  _GEN_28913 = _T_180 ? _GEN_28905 : _GEN_28657; // @[sequencer-master.scala 154:24]
  wire  _GEN_28914 = _T_180 ? _GEN_28906 : _GEN_28658; // @[sequencer-master.scala 154:24]
  wire  _GEN_28915 = _T_180 ? _GEN_28907 : _GEN_28659; // @[sequencer-master.scala 154:24]
  wire [1:0] _GEN_28916 = 3'h0 == tail ? 2'h0 : _GEN_28338; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28917 = 3'h1 == tail ? 2'h0 : _GEN_28339; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28918 = 3'h2 == tail ? 2'h0 : _GEN_28340; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28919 = 3'h3 == tail ? 2'h0 : _GEN_28341; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28920 = 3'h4 == tail ? 2'h0 : _GEN_28342; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28921 = 3'h5 == tail ? 2'h0 : _GEN_28343; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28922 = 3'h6 == tail ? 2'h0 : _GEN_28344; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [1:0] _GEN_28923 = 3'h7 == tail ? 2'h0 : _GEN_28345; // @[sequencer-master.scala 230:21 sequencer-master.scala 230:21]
  wire [3:0] _GEN_28924 = 3'h0 == tail ? 4'h0 : _GEN_28346; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28925 = 3'h1 == tail ? 4'h0 : _GEN_28347; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28926 = 3'h2 == tail ? 4'h0 : _GEN_28348; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28927 = 3'h3 == tail ? 4'h0 : _GEN_28349; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28928 = 3'h4 == tail ? 4'h0 : _GEN_28350; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28929 = 3'h5 == tail ? 4'h0 : _GEN_28351; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28930 = 3'h6 == tail ? 4'h0 : _GEN_28352; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [3:0] _GEN_28931 = 3'h7 == tail ? 4'h0 : _GEN_28353; // @[sequencer-master.scala 231:25 sequencer-master.scala 231:25]
  wire [2:0] _GEN_28932 = 3'h0 == tail ? 3'h0 : _GEN_28354; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28933 = 3'h1 == tail ? 3'h0 : _GEN_28355; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28934 = 3'h2 == tail ? 3'h0 : _GEN_28356; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28935 = 3'h3 == tail ? 3'h0 : _GEN_28357; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28936 = 3'h4 == tail ? 3'h0 : _GEN_28358; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28937 = 3'h5 == tail ? 3'h0 : _GEN_28359; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28938 = 3'h6 == tail ? 3'h0 : _GEN_28360; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire [2:0] _GEN_28939 = 3'h7 == tail ? 3'h0 : _GEN_28361; // @[sequencer-master.scala 232:25 sequencer-master.scala 232:25]
  wire  _GEN_28956 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28756; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28957 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28757; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28958 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28758; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28959 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28759; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28960 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28760; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28961 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28761; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28962 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28762; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28963 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28763; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_28964 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28444; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28965 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28445; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28966 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28446; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28967 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28447; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28968 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28448; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28969 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28449; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28970 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28450; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_28971 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28451; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29004 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28796; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29005 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28797; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29006 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28798; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29007 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28799; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29008 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28800; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29009 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28801; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29010 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28802; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29011 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28803; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29012 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28492; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29013 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28493; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29014 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28494; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29015 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28495; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29016 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28496; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29017 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28497; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29018 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28498; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29019 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28499; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29020 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28500; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29021 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28501; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29022 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28502; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29023 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28503; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29024 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28504; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29025 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28505; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29026 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28506; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29027 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28507; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29028 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28812; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29029 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28813; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29030 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28814; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29031 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28815; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29032 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28816; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29033 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28817; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29034 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28818; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29035 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28819; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29036 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28516; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29037 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28517; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29038 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28518; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29039 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28519; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29040 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28520; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29041 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28521; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29042 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28522; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29043 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28523; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29044 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28524; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29045 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28525; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29046 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28526; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29047 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28527; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29048 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28528; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29049 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28529; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29050 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28530; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29051 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28531; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29052 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28828; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29053 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28829; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29054 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28830; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29055 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28831; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29056 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28832; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29057 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28833; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29058 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28834; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29059 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28835; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29060 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28540; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29061 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28541; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29062 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28542; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29063 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28543; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29064 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28544; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29065 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28545; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29066 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28546; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29067 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28547; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29068 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28548; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29069 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28549; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29070 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28550; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29071 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28551; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29072 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28552; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29073 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28553; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29074 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28554; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29075 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28555; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29076 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28844; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29077 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28845; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29078 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28846; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29079 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28847; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29080 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28848; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29081 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28849; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29082 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28850; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29083 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28851; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29084 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28564; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29085 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28565; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29086 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28566; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29087 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28567; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29088 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28568; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29089 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28569; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29090 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28570; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29091 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28571; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29092 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28572; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29093 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28573; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29094 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28574; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29095 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28575; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29096 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28576; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29097 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28577; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29098 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28578; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29099 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28579; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29100 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28860; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29101 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28861; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29102 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28862; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29103 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28863; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29104 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28864; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29105 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28865; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29106 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28866; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29107 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28867; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29108 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28588; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29109 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28589; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29110 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28590; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29111 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28591; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29112 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28592; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29113 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28593; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29114 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28594; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29115 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28595; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29116 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28596; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29117 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28597; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29118 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28598; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29119 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28599; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29120 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28600; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29121 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28601; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29122 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28602; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29123 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28603; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29124 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28876; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29125 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28877; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29126 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28878; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29127 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28879; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29128 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28880; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29129 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28881; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29130 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28882; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29131 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28883; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29132 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28612; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29133 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28613; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29134 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28614; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29135 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28615; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29136 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28616; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29137 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28617; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29138 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28618; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29139 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28619; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29140 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28620; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29141 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28621; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29142 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28622; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29143 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28623; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29144 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28624; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29145 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28625; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29146 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28626; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29147 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28627; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29148 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28892; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29149 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28893; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29150 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28894; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29151 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28895; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29152 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28896; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29153 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28897; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29154 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28898; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29155 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28899; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29156 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28636; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29157 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28637; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29158 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28638; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29159 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28639; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29160 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28640; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29161 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28641; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29162 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28642; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29163 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28643; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29164 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28644; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29165 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28645; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29166 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28646; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29167 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28647; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29168 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28648; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29169 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28649; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29170 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28650; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29171 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28651; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29172 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28908; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29173 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28909; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29174 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28910; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29175 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28911; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29176 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28912; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29177 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28913; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29178 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28914; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29179 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28915; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29180 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28660; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29181 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28661; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29182 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28662; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29183 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28663; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29184 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28664; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29185 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28665; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29186 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28666; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29187 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28667; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29188 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28668; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29189 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28669; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29190 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28670; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29191 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28671; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29192 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28672; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29193 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28673; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29194 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28674; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29195 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28675; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29196 = 3'h0 == _T_1645 ? 1'h0 : _GEN_28676; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29197 = 3'h1 == _T_1645 ? 1'h0 : _GEN_28677; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29198 = 3'h2 == _T_1645 ? 1'h0 : _GEN_28678; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29199 = 3'h3 == _T_1645 ? 1'h0 : _GEN_28679; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29200 = 3'h4 == _T_1645 ? 1'h0 : _GEN_28680; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29201 = 3'h5 == _T_1645 ? 1'h0 : _GEN_28681; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29202 = 3'h6 == _T_1645 ? 1'h0 : _GEN_28682; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29203 = 3'h7 == _T_1645 ? 1'h0 : _GEN_28683; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29212 = _GEN_34121 | _GEN_28362; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29213 = _GEN_34122 | _GEN_28363; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29214 = _GEN_34123 | _GEN_28364; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29215 = _GEN_34124 | _GEN_28365; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29216 = _GEN_34125 | _GEN_28366; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29217 = _GEN_34126 | _GEN_28367; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29218 = _GEN_34127 | _GEN_28368; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29219 = _GEN_34128 | _GEN_28369; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29252 = 3'h0 == _T_1647 | (3'h0 == _T_1645 | (_GEN_32729 | _GEN_28018)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29253 = 3'h1 == _T_1647 | (3'h1 == _T_1645 | (_GEN_32730 | _GEN_28019)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29254 = 3'h2 == _T_1647 | (3'h2 == _T_1645 | (_GEN_32731 | _GEN_28020)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29255 = 3'h3 == _T_1647 | (3'h3 == _T_1645 | (_GEN_32732 | _GEN_28021)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29256 = 3'h4 == _T_1647 | (3'h4 == _T_1645 | (_GEN_32733 | _GEN_28022)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29257 = 3'h5 == _T_1647 | (3'h5 == _T_1645 | (_GEN_32734 | _GEN_28023)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29258 = 3'h6 == _T_1647 | (3'h6 == _T_1645 | (_GEN_32735 | _GEN_28024)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29259 = 3'h7 == _T_1647 | (3'h7 == _T_1645 | (_GEN_32736 | _GEN_28025)); // @[sequencer-master.scala 267:35 sequencer-master.scala 267:35]
  wire  _GEN_29268 = 3'h0 == _T_1647 ? 1'h0 : _GEN_28956; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29269 = 3'h1 == _T_1647 ? 1'h0 : _GEN_28957; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29270 = 3'h2 == _T_1647 ? 1'h0 : _GEN_28958; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29271 = 3'h3 == _T_1647 ? 1'h0 : _GEN_28959; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29272 = 3'h4 == _T_1647 ? 1'h0 : _GEN_28960; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29273 = 3'h5 == _T_1647 ? 1'h0 : _GEN_28961; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29274 = 3'h6 == _T_1647 ? 1'h0 : _GEN_28962; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29275 = 3'h7 == _T_1647 ? 1'h0 : _GEN_28963; // @[sequencer-master.scala 272:28 sequencer-master.scala 272:28]
  wire  _GEN_29276 = 3'h0 == _T_1647 ? 1'h0 : _GEN_28964; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29277 = 3'h1 == _T_1647 ? 1'h0 : _GEN_28965; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29278 = 3'h2 == _T_1647 ? 1'h0 : _GEN_28966; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29279 = 3'h3 == _T_1647 ? 1'h0 : _GEN_28967; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29280 = 3'h4 == _T_1647 ? 1'h0 : _GEN_28968; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29281 = 3'h5 == _T_1647 ? 1'h0 : _GEN_28969; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29282 = 3'h6 == _T_1647 ? 1'h0 : _GEN_28970; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29283 = 3'h7 == _T_1647 ? 1'h0 : _GEN_28971; // @[sequencer-master.scala 273:29 sequencer-master.scala 273:29]
  wire  _GEN_29308 = _GEN_36426 | (_GEN_34121 | (_GEN_32729 | _GEN_28074)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29309 = _GEN_36427 | (_GEN_34122 | (_GEN_32730 | _GEN_28075)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29310 = _GEN_36428 | (_GEN_34123 | (_GEN_32731 | _GEN_28076)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29311 = _GEN_36429 | (_GEN_34124 | (_GEN_32732 | _GEN_28077)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29312 = _GEN_36430 | (_GEN_34125 | (_GEN_32733 | _GEN_28078)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29313 = _GEN_36431 | (_GEN_34126 | (_GEN_32734 | _GEN_28079)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29314 = _GEN_36432 | (_GEN_34127 | (_GEN_32735 | _GEN_28080)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29315 = _GEN_36433 | (_GEN_34128 | (_GEN_32736 | _GEN_28081)); // @[sequencer-master.scala 188:42 sequencer-master.scala 188:42]
  wire  _GEN_29316 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29004; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29317 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29005; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29318 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29006; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29319 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29007; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29320 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29008; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29321 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29009; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29322 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29010; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29323 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29011; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29324 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29012; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29325 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29013; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29326 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29014; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29327 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29015; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29328 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29016; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29329 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29017; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29330 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29018; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29331 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29019; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29332 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29020; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29333 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29021; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29334 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29022; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29335 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29023; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29336 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29024; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29337 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29025; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29338 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29026; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29339 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29027; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29340 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29028; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29341 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29029; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29342 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29030; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29343 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29031; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29344 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29032; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29345 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29033; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29346 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29034; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29347 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29035; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29348 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29036; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29349 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29037; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29350 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29038; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29351 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29039; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29352 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29040; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29353 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29041; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29354 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29042; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29355 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29043; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29356 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29044; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29357 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29045; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29358 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29046; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29359 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29047; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29360 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29048; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29361 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29049; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29362 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29050; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29363 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29051; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29364 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29052; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29365 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29053; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29366 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29054; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29367 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29055; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29368 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29056; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29369 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29057; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29370 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29058; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29371 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29059; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29372 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29060; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29373 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29061; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29374 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29062; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29375 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29063; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29376 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29064; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29377 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29065; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29378 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29066; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29379 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29067; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29380 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29068; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29381 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29069; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29382 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29070; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29383 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29071; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29384 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29072; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29385 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29073; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29386 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29074; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29387 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29075; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29388 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29076; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29389 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29077; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29390 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29078; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29391 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29079; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29392 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29080; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29393 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29081; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29394 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29082; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29395 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29083; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29396 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29084; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29397 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29085; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29398 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29086; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29399 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29087; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29400 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29088; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29401 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29089; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29402 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29090; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29403 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29091; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29404 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29092; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29405 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29093; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29406 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29094; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29407 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29095; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29408 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29096; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29409 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29097; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29410 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29098; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29411 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29099; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29412 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29100; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29413 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29101; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29414 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29102; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29415 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29103; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29416 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29104; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29417 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29105; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29418 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29106; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29419 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29107; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29420 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29108; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29421 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29109; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29422 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29110; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29423 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29111; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29424 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29112; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29425 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29113; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29426 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29114; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29427 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29115; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29428 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29116; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29429 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29117; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29430 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29118; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29431 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29119; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29432 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29120; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29433 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29121; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29434 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29122; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29435 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29123; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29436 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29124; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29437 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29125; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29438 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29126; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29439 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29127; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29440 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29128; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29441 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29129; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29442 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29130; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29443 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29131; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29444 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29132; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29445 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29133; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29446 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29134; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29447 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29135; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29448 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29136; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29449 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29137; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29450 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29138; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29451 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29139; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29452 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29140; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29453 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29141; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29454 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29142; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29455 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29143; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29456 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29144; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29457 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29145; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29458 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29146; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29459 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29147; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29460 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29148; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29461 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29149; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29462 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29150; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29463 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29151; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29464 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29152; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29465 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29153; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29466 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29154; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29467 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29155; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29468 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29156; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29469 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29157; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29470 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29158; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29471 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29159; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29472 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29160; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29473 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29161; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29474 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29162; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29475 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29163; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29476 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29164; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29477 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29165; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29478 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29166; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29479 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29167; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29480 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29168; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29481 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29169; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29482 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29170; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29483 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29171; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29484 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29172; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29485 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29173; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29486 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29174; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29487 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29175; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29488 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29176; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29489 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29177; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29490 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29178; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29491 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29179; // @[sequencer-master.scala 183:52 sequencer-master.scala 183:52]
  wire  _GEN_29492 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29180; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29493 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29181; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29494 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29182; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29495 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29183; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29496 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29184; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29497 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29185; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29498 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29186; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29499 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29187; // @[sequencer-master.scala 184:52 sequencer-master.scala 184:52]
  wire  _GEN_29500 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29188; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29501 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29189; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29502 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29190; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29503 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29191; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29504 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29192; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29505 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29193; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29506 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29194; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29507 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29195; // @[sequencer-master.scala 185:52 sequencer-master.scala 185:52]
  wire  _GEN_29508 = 3'h0 == _T_1647 ? 1'h0 : _GEN_29196; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29509 = 3'h1 == _T_1647 ? 1'h0 : _GEN_29197; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29510 = 3'h2 == _T_1647 ? 1'h0 : _GEN_29198; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29511 = 3'h3 == _T_1647 ? 1'h0 : _GEN_29199; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29512 = 3'h4 == _T_1647 ? 1'h0 : _GEN_29200; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29513 = 3'h5 == _T_1647 ? 1'h0 : _GEN_29201; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29514 = 3'h6 == _T_1647 ? 1'h0 : _GEN_29202; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29515 = 3'h7 == _T_1647 ? 1'h0 : _GEN_29203; // @[sequencer-master.scala 283:19 sequencer-master.scala 283:19]
  wire  _GEN_29524 = _GEN_36426 | _GEN_26256; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29525 = _GEN_36427 | _GEN_26257; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29526 = _GEN_36428 | _GEN_26258; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29527 = _GEN_36429 | _GEN_26259; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29528 = _GEN_36430 | _GEN_26260; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29529 = _GEN_36431 | _GEN_26261; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29530 = _GEN_36432 | _GEN_26262; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire  _GEN_29531 = _GEN_36433 | _GEN_26263; // @[sequencer-master.scala 288:26 sequencer-master.scala 288:26]
  wire [7:0] _GEN_29572 = 3'h0 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28780; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29573 = 3'h1 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28781; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29574 = 3'h2 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28782; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29575 = 3'h3 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28783; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29576 = 3'h4 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28784; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29577 = 3'h5 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28785; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29578 = 3'h6 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28786; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29579 = 3'h7 == _T_1647 ? io_op_bits_reg_vp_id : _GEN_28787; // @[sequencer-master.scala 322:41 sequencer-master.scala 322:41]
  wire [7:0] _GEN_29612 = io_op_bits_base_vp_valid ? _GEN_29572 : _GEN_28780; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29613 = io_op_bits_base_vp_valid ? _GEN_29573 : _GEN_28781; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29614 = io_op_bits_base_vp_valid ? _GEN_29574 : _GEN_28782; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29615 = io_op_bits_base_vp_valid ? _GEN_29575 : _GEN_28783; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29616 = io_op_bits_base_vp_valid ? _GEN_29576 : _GEN_28784; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29617 = io_op_bits_base_vp_valid ? _GEN_29577 : _GEN_28785; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29618 = io_op_bits_base_vp_valid ? _GEN_29578 : _GEN_28786; // @[sequencer-master.scala 320:41]
  wire [7:0] _GEN_29619 = io_op_bits_base_vp_valid ? _GEN_29579 : _GEN_28787; // @[sequencer-master.scala 320:41]
  wire  _GEN_29620 = _GEN_36426 | _GEN_29316; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29621 = _GEN_36427 | _GEN_29317; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29622 = _GEN_36428 | _GEN_29318; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29623 = _GEN_36429 | _GEN_29319; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29624 = _GEN_36430 | _GEN_29320; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29625 = _GEN_36431 | _GEN_29321; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29626 = _GEN_36432 | _GEN_29322; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29627 = _GEN_36433 | _GEN_29323; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29628 = _T_26 ? _GEN_29620 : _GEN_29316; // @[sequencer-master.scala 154:24]
  wire  _GEN_29629 = _T_26 ? _GEN_29621 : _GEN_29317; // @[sequencer-master.scala 154:24]
  wire  _GEN_29630 = _T_26 ? _GEN_29622 : _GEN_29318; // @[sequencer-master.scala 154:24]
  wire  _GEN_29631 = _T_26 ? _GEN_29623 : _GEN_29319; // @[sequencer-master.scala 154:24]
  wire  _GEN_29632 = _T_26 ? _GEN_29624 : _GEN_29320; // @[sequencer-master.scala 154:24]
  wire  _GEN_29633 = _T_26 ? _GEN_29625 : _GEN_29321; // @[sequencer-master.scala 154:24]
  wire  _GEN_29634 = _T_26 ? _GEN_29626 : _GEN_29322; // @[sequencer-master.scala 154:24]
  wire  _GEN_29635 = _T_26 ? _GEN_29627 : _GEN_29323; // @[sequencer-master.scala 154:24]
  wire  _GEN_29636 = _GEN_36426 | _GEN_29340; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29637 = _GEN_36427 | _GEN_29341; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29638 = _GEN_36428 | _GEN_29342; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29639 = _GEN_36429 | _GEN_29343; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29640 = _GEN_36430 | _GEN_29344; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29641 = _GEN_36431 | _GEN_29345; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29642 = _GEN_36432 | _GEN_29346; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29643 = _GEN_36433 | _GEN_29347; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29644 = _T_48 ? _GEN_29636 : _GEN_29340; // @[sequencer-master.scala 154:24]
  wire  _GEN_29645 = _T_48 ? _GEN_29637 : _GEN_29341; // @[sequencer-master.scala 154:24]
  wire  _GEN_29646 = _T_48 ? _GEN_29638 : _GEN_29342; // @[sequencer-master.scala 154:24]
  wire  _GEN_29647 = _T_48 ? _GEN_29639 : _GEN_29343; // @[sequencer-master.scala 154:24]
  wire  _GEN_29648 = _T_48 ? _GEN_29640 : _GEN_29344; // @[sequencer-master.scala 154:24]
  wire  _GEN_29649 = _T_48 ? _GEN_29641 : _GEN_29345; // @[sequencer-master.scala 154:24]
  wire  _GEN_29650 = _T_48 ? _GEN_29642 : _GEN_29346; // @[sequencer-master.scala 154:24]
  wire  _GEN_29651 = _T_48 ? _GEN_29643 : _GEN_29347; // @[sequencer-master.scala 154:24]
  wire  _GEN_29652 = _GEN_36426 | _GEN_29364; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29653 = _GEN_36427 | _GEN_29365; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29654 = _GEN_36428 | _GEN_29366; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29655 = _GEN_36429 | _GEN_29367; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29656 = _GEN_36430 | _GEN_29368; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29657 = _GEN_36431 | _GEN_29369; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29658 = _GEN_36432 | _GEN_29370; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29659 = _GEN_36433 | _GEN_29371; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29660 = _T_70 ? _GEN_29652 : _GEN_29364; // @[sequencer-master.scala 154:24]
  wire  _GEN_29661 = _T_70 ? _GEN_29653 : _GEN_29365; // @[sequencer-master.scala 154:24]
  wire  _GEN_29662 = _T_70 ? _GEN_29654 : _GEN_29366; // @[sequencer-master.scala 154:24]
  wire  _GEN_29663 = _T_70 ? _GEN_29655 : _GEN_29367; // @[sequencer-master.scala 154:24]
  wire  _GEN_29664 = _T_70 ? _GEN_29656 : _GEN_29368; // @[sequencer-master.scala 154:24]
  wire  _GEN_29665 = _T_70 ? _GEN_29657 : _GEN_29369; // @[sequencer-master.scala 154:24]
  wire  _GEN_29666 = _T_70 ? _GEN_29658 : _GEN_29370; // @[sequencer-master.scala 154:24]
  wire  _GEN_29667 = _T_70 ? _GEN_29659 : _GEN_29371; // @[sequencer-master.scala 154:24]
  wire  _GEN_29668 = _GEN_36426 | _GEN_29388; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29669 = _GEN_36427 | _GEN_29389; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29670 = _GEN_36428 | _GEN_29390; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29671 = _GEN_36429 | _GEN_29391; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29672 = _GEN_36430 | _GEN_29392; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29673 = _GEN_36431 | _GEN_29393; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29674 = _GEN_36432 | _GEN_29394; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29675 = _GEN_36433 | _GEN_29395; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29676 = _T_92 ? _GEN_29668 : _GEN_29388; // @[sequencer-master.scala 154:24]
  wire  _GEN_29677 = _T_92 ? _GEN_29669 : _GEN_29389; // @[sequencer-master.scala 154:24]
  wire  _GEN_29678 = _T_92 ? _GEN_29670 : _GEN_29390; // @[sequencer-master.scala 154:24]
  wire  _GEN_29679 = _T_92 ? _GEN_29671 : _GEN_29391; // @[sequencer-master.scala 154:24]
  wire  _GEN_29680 = _T_92 ? _GEN_29672 : _GEN_29392; // @[sequencer-master.scala 154:24]
  wire  _GEN_29681 = _T_92 ? _GEN_29673 : _GEN_29393; // @[sequencer-master.scala 154:24]
  wire  _GEN_29682 = _T_92 ? _GEN_29674 : _GEN_29394; // @[sequencer-master.scala 154:24]
  wire  _GEN_29683 = _T_92 ? _GEN_29675 : _GEN_29395; // @[sequencer-master.scala 154:24]
  wire  _GEN_29684 = _GEN_36426 | _GEN_29412; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29685 = _GEN_36427 | _GEN_29413; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29686 = _GEN_36428 | _GEN_29414; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29687 = _GEN_36429 | _GEN_29415; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29688 = _GEN_36430 | _GEN_29416; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29689 = _GEN_36431 | _GEN_29417; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29690 = _GEN_36432 | _GEN_29418; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29691 = _GEN_36433 | _GEN_29419; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29692 = _T_114 ? _GEN_29684 : _GEN_29412; // @[sequencer-master.scala 154:24]
  wire  _GEN_29693 = _T_114 ? _GEN_29685 : _GEN_29413; // @[sequencer-master.scala 154:24]
  wire  _GEN_29694 = _T_114 ? _GEN_29686 : _GEN_29414; // @[sequencer-master.scala 154:24]
  wire  _GEN_29695 = _T_114 ? _GEN_29687 : _GEN_29415; // @[sequencer-master.scala 154:24]
  wire  _GEN_29696 = _T_114 ? _GEN_29688 : _GEN_29416; // @[sequencer-master.scala 154:24]
  wire  _GEN_29697 = _T_114 ? _GEN_29689 : _GEN_29417; // @[sequencer-master.scala 154:24]
  wire  _GEN_29698 = _T_114 ? _GEN_29690 : _GEN_29418; // @[sequencer-master.scala 154:24]
  wire  _GEN_29699 = _T_114 ? _GEN_29691 : _GEN_29419; // @[sequencer-master.scala 154:24]
  wire  _GEN_29700 = _GEN_36426 | _GEN_29436; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29701 = _GEN_36427 | _GEN_29437; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29702 = _GEN_36428 | _GEN_29438; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29703 = _GEN_36429 | _GEN_29439; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29704 = _GEN_36430 | _GEN_29440; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29705 = _GEN_36431 | _GEN_29441; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29706 = _GEN_36432 | _GEN_29442; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29707 = _GEN_36433 | _GEN_29443; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29708 = _T_136 ? _GEN_29700 : _GEN_29436; // @[sequencer-master.scala 154:24]
  wire  _GEN_29709 = _T_136 ? _GEN_29701 : _GEN_29437; // @[sequencer-master.scala 154:24]
  wire  _GEN_29710 = _T_136 ? _GEN_29702 : _GEN_29438; // @[sequencer-master.scala 154:24]
  wire  _GEN_29711 = _T_136 ? _GEN_29703 : _GEN_29439; // @[sequencer-master.scala 154:24]
  wire  _GEN_29712 = _T_136 ? _GEN_29704 : _GEN_29440; // @[sequencer-master.scala 154:24]
  wire  _GEN_29713 = _T_136 ? _GEN_29705 : _GEN_29441; // @[sequencer-master.scala 154:24]
  wire  _GEN_29714 = _T_136 ? _GEN_29706 : _GEN_29442; // @[sequencer-master.scala 154:24]
  wire  _GEN_29715 = _T_136 ? _GEN_29707 : _GEN_29443; // @[sequencer-master.scala 154:24]
  wire  _GEN_29716 = _GEN_36426 | _GEN_29460; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29717 = _GEN_36427 | _GEN_29461; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29718 = _GEN_36428 | _GEN_29462; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29719 = _GEN_36429 | _GEN_29463; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29720 = _GEN_36430 | _GEN_29464; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29721 = _GEN_36431 | _GEN_29465; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29722 = _GEN_36432 | _GEN_29466; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29723 = _GEN_36433 | _GEN_29467; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29724 = _T_158 ? _GEN_29716 : _GEN_29460; // @[sequencer-master.scala 154:24]
  wire  _GEN_29725 = _T_158 ? _GEN_29717 : _GEN_29461; // @[sequencer-master.scala 154:24]
  wire  _GEN_29726 = _T_158 ? _GEN_29718 : _GEN_29462; // @[sequencer-master.scala 154:24]
  wire  _GEN_29727 = _T_158 ? _GEN_29719 : _GEN_29463; // @[sequencer-master.scala 154:24]
  wire  _GEN_29728 = _T_158 ? _GEN_29720 : _GEN_29464; // @[sequencer-master.scala 154:24]
  wire  _GEN_29729 = _T_158 ? _GEN_29721 : _GEN_29465; // @[sequencer-master.scala 154:24]
  wire  _GEN_29730 = _T_158 ? _GEN_29722 : _GEN_29466; // @[sequencer-master.scala 154:24]
  wire  _GEN_29731 = _T_158 ? _GEN_29723 : _GEN_29467; // @[sequencer-master.scala 154:24]
  wire  _GEN_29732 = _GEN_36426 | _GEN_29484; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29733 = _GEN_36427 | _GEN_29485; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29734 = _GEN_36428 | _GEN_29486; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29735 = _GEN_36429 | _GEN_29487; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29736 = _GEN_36430 | _GEN_29488; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29737 = _GEN_36431 | _GEN_29489; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29738 = _GEN_36432 | _GEN_29490; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29739 = _GEN_36433 | _GEN_29491; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29740 = _T_180 ? _GEN_29732 : _GEN_29484; // @[sequencer-master.scala 154:24]
  wire  _GEN_29741 = _T_180 ? _GEN_29733 : _GEN_29485; // @[sequencer-master.scala 154:24]
  wire  _GEN_29742 = _T_180 ? _GEN_29734 : _GEN_29486; // @[sequencer-master.scala 154:24]
  wire  _GEN_29743 = _T_180 ? _GEN_29735 : _GEN_29487; // @[sequencer-master.scala 154:24]
  wire  _GEN_29744 = _T_180 ? _GEN_29736 : _GEN_29488; // @[sequencer-master.scala 154:24]
  wire  _GEN_29745 = _T_180 ? _GEN_29737 : _GEN_29489; // @[sequencer-master.scala 154:24]
  wire  _GEN_29746 = _T_180 ? _GEN_29738 : _GEN_29490; // @[sequencer-master.scala 154:24]
  wire  _GEN_29747 = _T_180 ? _GEN_29739 : _GEN_29491; // @[sequencer-master.scala 154:24]
  wire [7:0] _GEN_29788 = 3'h0 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26208; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29789 = 3'h1 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26209; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29790 = 3'h2 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26210; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29791 = 3'h3 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26211; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29792 = 3'h4 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26212; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29793 = 3'h5 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26213; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29794 = 3'h6 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26214; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29795 = 3'h7 == _T_1647 ? io_op_bits_reg_vd_id : _GEN_26215; // @[sequencer-master.scala 356:42 sequencer-master.scala 356:42]
  wire [7:0] _GEN_29836 = io_op_bits_base_vd_valid ? _GEN_29788 : _GEN_26208; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29837 = io_op_bits_base_vd_valid ? _GEN_29789 : _GEN_26209; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29838 = io_op_bits_base_vd_valid ? _GEN_29790 : _GEN_26210; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29839 = io_op_bits_base_vd_valid ? _GEN_29791 : _GEN_26211; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29840 = io_op_bits_base_vd_valid ? _GEN_29792 : _GEN_26212; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29841 = io_op_bits_base_vd_valid ? _GEN_29793 : _GEN_26213; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29842 = io_op_bits_base_vd_valid ? _GEN_29794 : _GEN_26214; // @[sequencer-master.scala 354:41]
  wire [7:0] _GEN_29843 = io_op_bits_base_vd_valid ? _GEN_29795 : _GEN_26215; // @[sequencer-master.scala 354:41]
  wire  _GEN_29844 = _GEN_36426 | _GEN_29628; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29845 = _GEN_36427 | _GEN_29629; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29846 = _GEN_36428 | _GEN_29630; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29847 = _GEN_36429 | _GEN_29631; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29848 = _GEN_36430 | _GEN_29632; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29849 = _GEN_36431 | _GEN_29633; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29850 = _GEN_36432 | _GEN_29634; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29851 = _GEN_36433 | _GEN_29635; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29852 = _T_1442 ? _GEN_29844 : _GEN_29628; // @[sequencer-master.scala 154:24]
  wire  _GEN_29853 = _T_1442 ? _GEN_29845 : _GEN_29629; // @[sequencer-master.scala 154:24]
  wire  _GEN_29854 = _T_1442 ? _GEN_29846 : _GEN_29630; // @[sequencer-master.scala 154:24]
  wire  _GEN_29855 = _T_1442 ? _GEN_29847 : _GEN_29631; // @[sequencer-master.scala 154:24]
  wire  _GEN_29856 = _T_1442 ? _GEN_29848 : _GEN_29632; // @[sequencer-master.scala 154:24]
  wire  _GEN_29857 = _T_1442 ? _GEN_29849 : _GEN_29633; // @[sequencer-master.scala 154:24]
  wire  _GEN_29858 = _T_1442 ? _GEN_29850 : _GEN_29634; // @[sequencer-master.scala 154:24]
  wire  _GEN_29859 = _T_1442 ? _GEN_29851 : _GEN_29635; // @[sequencer-master.scala 154:24]
  wire  _GEN_29860 = _GEN_36426 | _GEN_29644; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29861 = _GEN_36427 | _GEN_29645; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29862 = _GEN_36428 | _GEN_29646; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29863 = _GEN_36429 | _GEN_29647; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29864 = _GEN_36430 | _GEN_29648; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29865 = _GEN_36431 | _GEN_29649; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29866 = _GEN_36432 | _GEN_29650; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29867 = _GEN_36433 | _GEN_29651; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29868 = _T_1464 ? _GEN_29860 : _GEN_29644; // @[sequencer-master.scala 154:24]
  wire  _GEN_29869 = _T_1464 ? _GEN_29861 : _GEN_29645; // @[sequencer-master.scala 154:24]
  wire  _GEN_29870 = _T_1464 ? _GEN_29862 : _GEN_29646; // @[sequencer-master.scala 154:24]
  wire  _GEN_29871 = _T_1464 ? _GEN_29863 : _GEN_29647; // @[sequencer-master.scala 154:24]
  wire  _GEN_29872 = _T_1464 ? _GEN_29864 : _GEN_29648; // @[sequencer-master.scala 154:24]
  wire  _GEN_29873 = _T_1464 ? _GEN_29865 : _GEN_29649; // @[sequencer-master.scala 154:24]
  wire  _GEN_29874 = _T_1464 ? _GEN_29866 : _GEN_29650; // @[sequencer-master.scala 154:24]
  wire  _GEN_29875 = _T_1464 ? _GEN_29867 : _GEN_29651; // @[sequencer-master.scala 154:24]
  wire  _GEN_29876 = _GEN_36426 | _GEN_29660; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29877 = _GEN_36427 | _GEN_29661; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29878 = _GEN_36428 | _GEN_29662; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29879 = _GEN_36429 | _GEN_29663; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29880 = _GEN_36430 | _GEN_29664; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29881 = _GEN_36431 | _GEN_29665; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29882 = _GEN_36432 | _GEN_29666; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29883 = _GEN_36433 | _GEN_29667; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29884 = _T_1486 ? _GEN_29876 : _GEN_29660; // @[sequencer-master.scala 154:24]
  wire  _GEN_29885 = _T_1486 ? _GEN_29877 : _GEN_29661; // @[sequencer-master.scala 154:24]
  wire  _GEN_29886 = _T_1486 ? _GEN_29878 : _GEN_29662; // @[sequencer-master.scala 154:24]
  wire  _GEN_29887 = _T_1486 ? _GEN_29879 : _GEN_29663; // @[sequencer-master.scala 154:24]
  wire  _GEN_29888 = _T_1486 ? _GEN_29880 : _GEN_29664; // @[sequencer-master.scala 154:24]
  wire  _GEN_29889 = _T_1486 ? _GEN_29881 : _GEN_29665; // @[sequencer-master.scala 154:24]
  wire  _GEN_29890 = _T_1486 ? _GEN_29882 : _GEN_29666; // @[sequencer-master.scala 154:24]
  wire  _GEN_29891 = _T_1486 ? _GEN_29883 : _GEN_29667; // @[sequencer-master.scala 154:24]
  wire  _GEN_29892 = _GEN_36426 | _GEN_29676; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29893 = _GEN_36427 | _GEN_29677; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29894 = _GEN_36428 | _GEN_29678; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29895 = _GEN_36429 | _GEN_29679; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29896 = _GEN_36430 | _GEN_29680; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29897 = _GEN_36431 | _GEN_29681; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29898 = _GEN_36432 | _GEN_29682; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29899 = _GEN_36433 | _GEN_29683; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29900 = _T_1508 ? _GEN_29892 : _GEN_29676; // @[sequencer-master.scala 154:24]
  wire  _GEN_29901 = _T_1508 ? _GEN_29893 : _GEN_29677; // @[sequencer-master.scala 154:24]
  wire  _GEN_29902 = _T_1508 ? _GEN_29894 : _GEN_29678; // @[sequencer-master.scala 154:24]
  wire  _GEN_29903 = _T_1508 ? _GEN_29895 : _GEN_29679; // @[sequencer-master.scala 154:24]
  wire  _GEN_29904 = _T_1508 ? _GEN_29896 : _GEN_29680; // @[sequencer-master.scala 154:24]
  wire  _GEN_29905 = _T_1508 ? _GEN_29897 : _GEN_29681; // @[sequencer-master.scala 154:24]
  wire  _GEN_29906 = _T_1508 ? _GEN_29898 : _GEN_29682; // @[sequencer-master.scala 154:24]
  wire  _GEN_29907 = _T_1508 ? _GEN_29899 : _GEN_29683; // @[sequencer-master.scala 154:24]
  wire  _GEN_29908 = _GEN_36426 | _GEN_29692; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29909 = _GEN_36427 | _GEN_29693; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29910 = _GEN_36428 | _GEN_29694; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29911 = _GEN_36429 | _GEN_29695; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29912 = _GEN_36430 | _GEN_29696; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29913 = _GEN_36431 | _GEN_29697; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29914 = _GEN_36432 | _GEN_29698; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29915 = _GEN_36433 | _GEN_29699; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29916 = _T_1530 ? _GEN_29908 : _GEN_29692; // @[sequencer-master.scala 154:24]
  wire  _GEN_29917 = _T_1530 ? _GEN_29909 : _GEN_29693; // @[sequencer-master.scala 154:24]
  wire  _GEN_29918 = _T_1530 ? _GEN_29910 : _GEN_29694; // @[sequencer-master.scala 154:24]
  wire  _GEN_29919 = _T_1530 ? _GEN_29911 : _GEN_29695; // @[sequencer-master.scala 154:24]
  wire  _GEN_29920 = _T_1530 ? _GEN_29912 : _GEN_29696; // @[sequencer-master.scala 154:24]
  wire  _GEN_29921 = _T_1530 ? _GEN_29913 : _GEN_29697; // @[sequencer-master.scala 154:24]
  wire  _GEN_29922 = _T_1530 ? _GEN_29914 : _GEN_29698; // @[sequencer-master.scala 154:24]
  wire  _GEN_29923 = _T_1530 ? _GEN_29915 : _GEN_29699; // @[sequencer-master.scala 154:24]
  wire  _GEN_29924 = _GEN_36426 | _GEN_29708; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29925 = _GEN_36427 | _GEN_29709; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29926 = _GEN_36428 | _GEN_29710; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29927 = _GEN_36429 | _GEN_29711; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29928 = _GEN_36430 | _GEN_29712; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29929 = _GEN_36431 | _GEN_29713; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29930 = _GEN_36432 | _GEN_29714; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29931 = _GEN_36433 | _GEN_29715; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29932 = _T_1552 ? _GEN_29924 : _GEN_29708; // @[sequencer-master.scala 154:24]
  wire  _GEN_29933 = _T_1552 ? _GEN_29925 : _GEN_29709; // @[sequencer-master.scala 154:24]
  wire  _GEN_29934 = _T_1552 ? _GEN_29926 : _GEN_29710; // @[sequencer-master.scala 154:24]
  wire  _GEN_29935 = _T_1552 ? _GEN_29927 : _GEN_29711; // @[sequencer-master.scala 154:24]
  wire  _GEN_29936 = _T_1552 ? _GEN_29928 : _GEN_29712; // @[sequencer-master.scala 154:24]
  wire  _GEN_29937 = _T_1552 ? _GEN_29929 : _GEN_29713; // @[sequencer-master.scala 154:24]
  wire  _GEN_29938 = _T_1552 ? _GEN_29930 : _GEN_29714; // @[sequencer-master.scala 154:24]
  wire  _GEN_29939 = _T_1552 ? _GEN_29931 : _GEN_29715; // @[sequencer-master.scala 154:24]
  wire  _GEN_29940 = _GEN_36426 | _GEN_29724; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29941 = _GEN_36427 | _GEN_29725; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29942 = _GEN_36428 | _GEN_29726; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29943 = _GEN_36429 | _GEN_29727; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29944 = _GEN_36430 | _GEN_29728; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29945 = _GEN_36431 | _GEN_29729; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29946 = _GEN_36432 | _GEN_29730; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29947 = _GEN_36433 | _GEN_29731; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29948 = _T_1574 ? _GEN_29940 : _GEN_29724; // @[sequencer-master.scala 154:24]
  wire  _GEN_29949 = _T_1574 ? _GEN_29941 : _GEN_29725; // @[sequencer-master.scala 154:24]
  wire  _GEN_29950 = _T_1574 ? _GEN_29942 : _GEN_29726; // @[sequencer-master.scala 154:24]
  wire  _GEN_29951 = _T_1574 ? _GEN_29943 : _GEN_29727; // @[sequencer-master.scala 154:24]
  wire  _GEN_29952 = _T_1574 ? _GEN_29944 : _GEN_29728; // @[sequencer-master.scala 154:24]
  wire  _GEN_29953 = _T_1574 ? _GEN_29945 : _GEN_29729; // @[sequencer-master.scala 154:24]
  wire  _GEN_29954 = _T_1574 ? _GEN_29946 : _GEN_29730; // @[sequencer-master.scala 154:24]
  wire  _GEN_29955 = _T_1574 ? _GEN_29947 : _GEN_29731; // @[sequencer-master.scala 154:24]
  wire  _GEN_29956 = _GEN_36426 | _GEN_29740; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29957 = _GEN_36427 | _GEN_29741; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29958 = _GEN_36428 | _GEN_29742; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29959 = _GEN_36429 | _GEN_29743; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29960 = _GEN_36430 | _GEN_29744; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29961 = _GEN_36431 | _GEN_29745; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29962 = _GEN_36432 | _GEN_29746; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29963 = _GEN_36433 | _GEN_29747; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29964 = _T_1596 ? _GEN_29956 : _GEN_29740; // @[sequencer-master.scala 154:24]
  wire  _GEN_29965 = _T_1596 ? _GEN_29957 : _GEN_29741; // @[sequencer-master.scala 154:24]
  wire  _GEN_29966 = _T_1596 ? _GEN_29958 : _GEN_29742; // @[sequencer-master.scala 154:24]
  wire  _GEN_29967 = _T_1596 ? _GEN_29959 : _GEN_29743; // @[sequencer-master.scala 154:24]
  wire  _GEN_29968 = _T_1596 ? _GEN_29960 : _GEN_29744; // @[sequencer-master.scala 154:24]
  wire  _GEN_29969 = _T_1596 ? _GEN_29961 : _GEN_29745; // @[sequencer-master.scala 154:24]
  wire  _GEN_29970 = _T_1596 ? _GEN_29962 : _GEN_29746; // @[sequencer-master.scala 154:24]
  wire  _GEN_29971 = _T_1596 ? _GEN_29963 : _GEN_29747; // @[sequencer-master.scala 154:24]
  wire  _GEN_29996 = _GEN_36426 & _GEN_34121 | _GEN_29852; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29997 = _GEN_36426 & _GEN_34122 | _GEN_29868; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29998 = _GEN_36426 & _GEN_34123 | _GEN_29884; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_29999 = _GEN_36426 & _GEN_34124 | _GEN_29900; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30000 = _GEN_36426 & _GEN_34125 | _GEN_29916; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30001 = _GEN_36426 & _GEN_34126 | _GEN_29932; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30002 = _GEN_36426 & _GEN_34127 | _GEN_29948; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30003 = _GEN_36426 & _GEN_34128 | _GEN_29964; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30004 = _GEN_36427 & _GEN_34121 | _GEN_29853; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30005 = _GEN_36427 & _GEN_34122 | _GEN_29869; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30006 = _GEN_36427 & _GEN_34123 | _GEN_29885; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30007 = _GEN_36427 & _GEN_34124 | _GEN_29901; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30008 = _GEN_36427 & _GEN_34125 | _GEN_29917; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30009 = _GEN_36427 & _GEN_34126 | _GEN_29933; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30010 = _GEN_36427 & _GEN_34127 | _GEN_29949; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30011 = _GEN_36427 & _GEN_34128 | _GEN_29965; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30012 = _GEN_36428 & _GEN_34121 | _GEN_29854; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30013 = _GEN_36428 & _GEN_34122 | _GEN_29870; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30014 = _GEN_36428 & _GEN_34123 | _GEN_29886; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30015 = _GEN_36428 & _GEN_34124 | _GEN_29902; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30016 = _GEN_36428 & _GEN_34125 | _GEN_29918; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30017 = _GEN_36428 & _GEN_34126 | _GEN_29934; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30018 = _GEN_36428 & _GEN_34127 | _GEN_29950; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30019 = _GEN_36428 & _GEN_34128 | _GEN_29966; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30020 = _GEN_36429 & _GEN_34121 | _GEN_29855; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30021 = _GEN_36429 & _GEN_34122 | _GEN_29871; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30022 = _GEN_36429 & _GEN_34123 | _GEN_29887; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30023 = _GEN_36429 & _GEN_34124 | _GEN_29903; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30024 = _GEN_36429 & _GEN_34125 | _GEN_29919; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30025 = _GEN_36429 & _GEN_34126 | _GEN_29935; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30026 = _GEN_36429 & _GEN_34127 | _GEN_29951; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30027 = _GEN_36429 & _GEN_34128 | _GEN_29967; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30028 = _GEN_36430 & _GEN_34121 | _GEN_29856; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30029 = _GEN_36430 & _GEN_34122 | _GEN_29872; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30030 = _GEN_36430 & _GEN_34123 | _GEN_29888; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30031 = _GEN_36430 & _GEN_34124 | _GEN_29904; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30032 = _GEN_36430 & _GEN_34125 | _GEN_29920; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30033 = _GEN_36430 & _GEN_34126 | _GEN_29936; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30034 = _GEN_36430 & _GEN_34127 | _GEN_29952; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30035 = _GEN_36430 & _GEN_34128 | _GEN_29968; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30036 = _GEN_36431 & _GEN_34121 | _GEN_29857; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30037 = _GEN_36431 & _GEN_34122 | _GEN_29873; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30038 = _GEN_36431 & _GEN_34123 | _GEN_29889; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30039 = _GEN_36431 & _GEN_34124 | _GEN_29905; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30040 = _GEN_36431 & _GEN_34125 | _GEN_29921; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30041 = _GEN_36431 & _GEN_34126 | _GEN_29937; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30042 = _GEN_36431 & _GEN_34127 | _GEN_29953; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30043 = _GEN_36431 & _GEN_34128 | _GEN_29969; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30044 = _GEN_36432 & _GEN_34121 | _GEN_29858; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30045 = _GEN_36432 & _GEN_34122 | _GEN_29874; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30046 = _GEN_36432 & _GEN_34123 | _GEN_29890; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30047 = _GEN_36432 & _GEN_34124 | _GEN_29906; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30048 = _GEN_36432 & _GEN_34125 | _GEN_29922; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30049 = _GEN_36432 & _GEN_34126 | _GEN_29938; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30050 = _GEN_36432 & _GEN_34127 | _GEN_29954; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30051 = _GEN_36432 & _GEN_34128 | _GEN_29970; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30052 = _GEN_36433 & _GEN_34121 | _GEN_29859; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30053 = _GEN_36433 & _GEN_34122 | _GEN_29875; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30054 = _GEN_36433 & _GEN_34123 | _GEN_29891; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30055 = _GEN_36433 & _GEN_34124 | _GEN_29907; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30056 = _GEN_36433 & _GEN_34125 | _GEN_29923; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30057 = _GEN_36433 & _GEN_34126 | _GEN_29939; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30058 = _GEN_36433 & _GEN_34127 | _GEN_29955; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30059 = _GEN_36433 & _GEN_34128 | _GEN_29971; // @[sequencer-master.scala 131:52 sequencer-master.scala 131:52]
  wire  _GEN_30060 = io_op_bits_active_vst ? _GEN_29252 : _GEN_28018; // @[sequencer-master.scala 654:38]
  wire  _GEN_30061 = io_op_bits_active_vst ? _GEN_29253 : _GEN_28019; // @[sequencer-master.scala 654:38]
  wire  _GEN_30062 = io_op_bits_active_vst ? _GEN_29254 : _GEN_28020; // @[sequencer-master.scala 654:38]
  wire  _GEN_30063 = io_op_bits_active_vst ? _GEN_29255 : _GEN_28021; // @[sequencer-master.scala 654:38]
  wire  _GEN_30064 = io_op_bits_active_vst ? _GEN_29256 : _GEN_28022; // @[sequencer-master.scala 654:38]
  wire  _GEN_30065 = io_op_bits_active_vst ? _GEN_29257 : _GEN_28023; // @[sequencer-master.scala 654:38]
  wire  _GEN_30066 = io_op_bits_active_vst ? _GEN_29258 : _GEN_28024; // @[sequencer-master.scala 654:38]
  wire  _GEN_30067 = io_op_bits_active_vst ? _GEN_29259 : _GEN_28025; // @[sequencer-master.scala 654:38]
  wire  _GEN_30116 = io_op_bits_active_vst ? _GEN_29308 : _GEN_28074; // @[sequencer-master.scala 654:38]
  wire  _GEN_30117 = io_op_bits_active_vst ? _GEN_29309 : _GEN_28075; // @[sequencer-master.scala 654:38]
  wire  _GEN_30118 = io_op_bits_active_vst ? _GEN_29310 : _GEN_28076; // @[sequencer-master.scala 654:38]
  wire  _GEN_30119 = io_op_bits_active_vst ? _GEN_29311 : _GEN_28077; // @[sequencer-master.scala 654:38]
  wire  _GEN_30120 = io_op_bits_active_vst ? _GEN_29312 : _GEN_28078; // @[sequencer-master.scala 654:38]
  wire  _GEN_30121 = io_op_bits_active_vst ? _GEN_29313 : _GEN_28079; // @[sequencer-master.scala 654:38]
  wire  _GEN_30122 = io_op_bits_active_vst ? _GEN_29314 : _GEN_28080; // @[sequencer-master.scala 654:38]
  wire  _GEN_30123 = io_op_bits_active_vst ? _GEN_29315 : _GEN_28081; // @[sequencer-master.scala 654:38]
  wire  _GEN_30124 = io_op_bits_active_vst ? _GEN_29996 : _GEN_28082; // @[sequencer-master.scala 654:38]
  wire  _GEN_30125 = io_op_bits_active_vst ? _GEN_30004 : _GEN_28083; // @[sequencer-master.scala 654:38]
  wire  _GEN_30126 = io_op_bits_active_vst ? _GEN_30012 : _GEN_28084; // @[sequencer-master.scala 654:38]
  wire  _GEN_30127 = io_op_bits_active_vst ? _GEN_30020 : _GEN_28085; // @[sequencer-master.scala 654:38]
  wire  _GEN_30128 = io_op_bits_active_vst ? _GEN_30028 : _GEN_28086; // @[sequencer-master.scala 654:38]
  wire  _GEN_30129 = io_op_bits_active_vst ? _GEN_30036 : _GEN_28087; // @[sequencer-master.scala 654:38]
  wire  _GEN_30130 = io_op_bits_active_vst ? _GEN_30044 : _GEN_28088; // @[sequencer-master.scala 654:38]
  wire  _GEN_30131 = io_op_bits_active_vst ? _GEN_30052 : _GEN_28089; // @[sequencer-master.scala 654:38]
  wire  _GEN_30132 = io_op_bits_active_vst ? _GEN_29324 : _GEN_28090; // @[sequencer-master.scala 654:38]
  wire  _GEN_30133 = io_op_bits_active_vst ? _GEN_29325 : _GEN_28091; // @[sequencer-master.scala 654:38]
  wire  _GEN_30134 = io_op_bits_active_vst ? _GEN_29326 : _GEN_28092; // @[sequencer-master.scala 654:38]
  wire  _GEN_30135 = io_op_bits_active_vst ? _GEN_29327 : _GEN_28093; // @[sequencer-master.scala 654:38]
  wire  _GEN_30136 = io_op_bits_active_vst ? _GEN_29328 : _GEN_28094; // @[sequencer-master.scala 654:38]
  wire  _GEN_30137 = io_op_bits_active_vst ? _GEN_29329 : _GEN_28095; // @[sequencer-master.scala 654:38]
  wire  _GEN_30138 = io_op_bits_active_vst ? _GEN_29330 : _GEN_28096; // @[sequencer-master.scala 654:38]
  wire  _GEN_30139 = io_op_bits_active_vst ? _GEN_29331 : _GEN_28097; // @[sequencer-master.scala 654:38]
  wire  _GEN_30140 = io_op_bits_active_vst ? _GEN_29332 : _GEN_28098; // @[sequencer-master.scala 654:38]
  wire  _GEN_30141 = io_op_bits_active_vst ? _GEN_29333 : _GEN_28099; // @[sequencer-master.scala 654:38]
  wire  _GEN_30142 = io_op_bits_active_vst ? _GEN_29334 : _GEN_28100; // @[sequencer-master.scala 654:38]
  wire  _GEN_30143 = io_op_bits_active_vst ? _GEN_29335 : _GEN_28101; // @[sequencer-master.scala 654:38]
  wire  _GEN_30144 = io_op_bits_active_vst ? _GEN_29336 : _GEN_28102; // @[sequencer-master.scala 654:38]
  wire  _GEN_30145 = io_op_bits_active_vst ? _GEN_29337 : _GEN_28103; // @[sequencer-master.scala 654:38]
  wire  _GEN_30146 = io_op_bits_active_vst ? _GEN_29338 : _GEN_28104; // @[sequencer-master.scala 654:38]
  wire  _GEN_30147 = io_op_bits_active_vst ? _GEN_29339 : _GEN_28105; // @[sequencer-master.scala 654:38]
  wire  _GEN_30148 = io_op_bits_active_vst ? _GEN_29997 : _GEN_28106; // @[sequencer-master.scala 654:38]
  wire  _GEN_30149 = io_op_bits_active_vst ? _GEN_30005 : _GEN_28107; // @[sequencer-master.scala 654:38]
  wire  _GEN_30150 = io_op_bits_active_vst ? _GEN_30013 : _GEN_28108; // @[sequencer-master.scala 654:38]
  wire  _GEN_30151 = io_op_bits_active_vst ? _GEN_30021 : _GEN_28109; // @[sequencer-master.scala 654:38]
  wire  _GEN_30152 = io_op_bits_active_vst ? _GEN_30029 : _GEN_28110; // @[sequencer-master.scala 654:38]
  wire  _GEN_30153 = io_op_bits_active_vst ? _GEN_30037 : _GEN_28111; // @[sequencer-master.scala 654:38]
  wire  _GEN_30154 = io_op_bits_active_vst ? _GEN_30045 : _GEN_28112; // @[sequencer-master.scala 654:38]
  wire  _GEN_30155 = io_op_bits_active_vst ? _GEN_30053 : _GEN_28113; // @[sequencer-master.scala 654:38]
  wire  _GEN_30156 = io_op_bits_active_vst ? _GEN_29348 : _GEN_28114; // @[sequencer-master.scala 654:38]
  wire  _GEN_30157 = io_op_bits_active_vst ? _GEN_29349 : _GEN_28115; // @[sequencer-master.scala 654:38]
  wire  _GEN_30158 = io_op_bits_active_vst ? _GEN_29350 : _GEN_28116; // @[sequencer-master.scala 654:38]
  wire  _GEN_30159 = io_op_bits_active_vst ? _GEN_29351 : _GEN_28117; // @[sequencer-master.scala 654:38]
  wire  _GEN_30160 = io_op_bits_active_vst ? _GEN_29352 : _GEN_28118; // @[sequencer-master.scala 654:38]
  wire  _GEN_30161 = io_op_bits_active_vst ? _GEN_29353 : _GEN_28119; // @[sequencer-master.scala 654:38]
  wire  _GEN_30162 = io_op_bits_active_vst ? _GEN_29354 : _GEN_28120; // @[sequencer-master.scala 654:38]
  wire  _GEN_30163 = io_op_bits_active_vst ? _GEN_29355 : _GEN_28121; // @[sequencer-master.scala 654:38]
  wire  _GEN_30164 = io_op_bits_active_vst ? _GEN_29356 : _GEN_28122; // @[sequencer-master.scala 654:38]
  wire  _GEN_30165 = io_op_bits_active_vst ? _GEN_29357 : _GEN_28123; // @[sequencer-master.scala 654:38]
  wire  _GEN_30166 = io_op_bits_active_vst ? _GEN_29358 : _GEN_28124; // @[sequencer-master.scala 654:38]
  wire  _GEN_30167 = io_op_bits_active_vst ? _GEN_29359 : _GEN_28125; // @[sequencer-master.scala 654:38]
  wire  _GEN_30168 = io_op_bits_active_vst ? _GEN_29360 : _GEN_28126; // @[sequencer-master.scala 654:38]
  wire  _GEN_30169 = io_op_bits_active_vst ? _GEN_29361 : _GEN_28127; // @[sequencer-master.scala 654:38]
  wire  _GEN_30170 = io_op_bits_active_vst ? _GEN_29362 : _GEN_28128; // @[sequencer-master.scala 654:38]
  wire  _GEN_30171 = io_op_bits_active_vst ? _GEN_29363 : _GEN_28129; // @[sequencer-master.scala 654:38]
  wire  _GEN_30172 = io_op_bits_active_vst ? _GEN_29998 : _GEN_28130; // @[sequencer-master.scala 654:38]
  wire  _GEN_30173 = io_op_bits_active_vst ? _GEN_30006 : _GEN_28131; // @[sequencer-master.scala 654:38]
  wire  _GEN_30174 = io_op_bits_active_vst ? _GEN_30014 : _GEN_28132; // @[sequencer-master.scala 654:38]
  wire  _GEN_30175 = io_op_bits_active_vst ? _GEN_30022 : _GEN_28133; // @[sequencer-master.scala 654:38]
  wire  _GEN_30176 = io_op_bits_active_vst ? _GEN_30030 : _GEN_28134; // @[sequencer-master.scala 654:38]
  wire  _GEN_30177 = io_op_bits_active_vst ? _GEN_30038 : _GEN_28135; // @[sequencer-master.scala 654:38]
  wire  _GEN_30178 = io_op_bits_active_vst ? _GEN_30046 : _GEN_28136; // @[sequencer-master.scala 654:38]
  wire  _GEN_30179 = io_op_bits_active_vst ? _GEN_30054 : _GEN_28137; // @[sequencer-master.scala 654:38]
  wire  _GEN_30180 = io_op_bits_active_vst ? _GEN_29372 : _GEN_28138; // @[sequencer-master.scala 654:38]
  wire  _GEN_30181 = io_op_bits_active_vst ? _GEN_29373 : _GEN_28139; // @[sequencer-master.scala 654:38]
  wire  _GEN_30182 = io_op_bits_active_vst ? _GEN_29374 : _GEN_28140; // @[sequencer-master.scala 654:38]
  wire  _GEN_30183 = io_op_bits_active_vst ? _GEN_29375 : _GEN_28141; // @[sequencer-master.scala 654:38]
  wire  _GEN_30184 = io_op_bits_active_vst ? _GEN_29376 : _GEN_28142; // @[sequencer-master.scala 654:38]
  wire  _GEN_30185 = io_op_bits_active_vst ? _GEN_29377 : _GEN_28143; // @[sequencer-master.scala 654:38]
  wire  _GEN_30186 = io_op_bits_active_vst ? _GEN_29378 : _GEN_28144; // @[sequencer-master.scala 654:38]
  wire  _GEN_30187 = io_op_bits_active_vst ? _GEN_29379 : _GEN_28145; // @[sequencer-master.scala 654:38]
  wire  _GEN_30188 = io_op_bits_active_vst ? _GEN_29380 : _GEN_28146; // @[sequencer-master.scala 654:38]
  wire  _GEN_30189 = io_op_bits_active_vst ? _GEN_29381 : _GEN_28147; // @[sequencer-master.scala 654:38]
  wire  _GEN_30190 = io_op_bits_active_vst ? _GEN_29382 : _GEN_28148; // @[sequencer-master.scala 654:38]
  wire  _GEN_30191 = io_op_bits_active_vst ? _GEN_29383 : _GEN_28149; // @[sequencer-master.scala 654:38]
  wire  _GEN_30192 = io_op_bits_active_vst ? _GEN_29384 : _GEN_28150; // @[sequencer-master.scala 654:38]
  wire  _GEN_30193 = io_op_bits_active_vst ? _GEN_29385 : _GEN_28151; // @[sequencer-master.scala 654:38]
  wire  _GEN_30194 = io_op_bits_active_vst ? _GEN_29386 : _GEN_28152; // @[sequencer-master.scala 654:38]
  wire  _GEN_30195 = io_op_bits_active_vst ? _GEN_29387 : _GEN_28153; // @[sequencer-master.scala 654:38]
  wire  _GEN_30196 = io_op_bits_active_vst ? _GEN_29999 : _GEN_28154; // @[sequencer-master.scala 654:38]
  wire  _GEN_30197 = io_op_bits_active_vst ? _GEN_30007 : _GEN_28155; // @[sequencer-master.scala 654:38]
  wire  _GEN_30198 = io_op_bits_active_vst ? _GEN_30015 : _GEN_28156; // @[sequencer-master.scala 654:38]
  wire  _GEN_30199 = io_op_bits_active_vst ? _GEN_30023 : _GEN_28157; // @[sequencer-master.scala 654:38]
  wire  _GEN_30200 = io_op_bits_active_vst ? _GEN_30031 : _GEN_28158; // @[sequencer-master.scala 654:38]
  wire  _GEN_30201 = io_op_bits_active_vst ? _GEN_30039 : _GEN_28159; // @[sequencer-master.scala 654:38]
  wire  _GEN_30202 = io_op_bits_active_vst ? _GEN_30047 : _GEN_28160; // @[sequencer-master.scala 654:38]
  wire  _GEN_30203 = io_op_bits_active_vst ? _GEN_30055 : _GEN_28161; // @[sequencer-master.scala 654:38]
  wire  _GEN_30204 = io_op_bits_active_vst ? _GEN_29396 : _GEN_28162; // @[sequencer-master.scala 654:38]
  wire  _GEN_30205 = io_op_bits_active_vst ? _GEN_29397 : _GEN_28163; // @[sequencer-master.scala 654:38]
  wire  _GEN_30206 = io_op_bits_active_vst ? _GEN_29398 : _GEN_28164; // @[sequencer-master.scala 654:38]
  wire  _GEN_30207 = io_op_bits_active_vst ? _GEN_29399 : _GEN_28165; // @[sequencer-master.scala 654:38]
  wire  _GEN_30208 = io_op_bits_active_vst ? _GEN_29400 : _GEN_28166; // @[sequencer-master.scala 654:38]
  wire  _GEN_30209 = io_op_bits_active_vst ? _GEN_29401 : _GEN_28167; // @[sequencer-master.scala 654:38]
  wire  _GEN_30210 = io_op_bits_active_vst ? _GEN_29402 : _GEN_28168; // @[sequencer-master.scala 654:38]
  wire  _GEN_30211 = io_op_bits_active_vst ? _GEN_29403 : _GEN_28169; // @[sequencer-master.scala 654:38]
  wire  _GEN_30212 = io_op_bits_active_vst ? _GEN_29404 : _GEN_28170; // @[sequencer-master.scala 654:38]
  wire  _GEN_30213 = io_op_bits_active_vst ? _GEN_29405 : _GEN_28171; // @[sequencer-master.scala 654:38]
  wire  _GEN_30214 = io_op_bits_active_vst ? _GEN_29406 : _GEN_28172; // @[sequencer-master.scala 654:38]
  wire  _GEN_30215 = io_op_bits_active_vst ? _GEN_29407 : _GEN_28173; // @[sequencer-master.scala 654:38]
  wire  _GEN_30216 = io_op_bits_active_vst ? _GEN_29408 : _GEN_28174; // @[sequencer-master.scala 654:38]
  wire  _GEN_30217 = io_op_bits_active_vst ? _GEN_29409 : _GEN_28175; // @[sequencer-master.scala 654:38]
  wire  _GEN_30218 = io_op_bits_active_vst ? _GEN_29410 : _GEN_28176; // @[sequencer-master.scala 654:38]
  wire  _GEN_30219 = io_op_bits_active_vst ? _GEN_29411 : _GEN_28177; // @[sequencer-master.scala 654:38]
  wire  _GEN_30220 = io_op_bits_active_vst ? _GEN_30000 : _GEN_28178; // @[sequencer-master.scala 654:38]
  wire  _GEN_30221 = io_op_bits_active_vst ? _GEN_30008 : _GEN_28179; // @[sequencer-master.scala 654:38]
  wire  _GEN_30222 = io_op_bits_active_vst ? _GEN_30016 : _GEN_28180; // @[sequencer-master.scala 654:38]
  wire  _GEN_30223 = io_op_bits_active_vst ? _GEN_30024 : _GEN_28181; // @[sequencer-master.scala 654:38]
  wire  _GEN_30224 = io_op_bits_active_vst ? _GEN_30032 : _GEN_28182; // @[sequencer-master.scala 654:38]
  wire  _GEN_30225 = io_op_bits_active_vst ? _GEN_30040 : _GEN_28183; // @[sequencer-master.scala 654:38]
  wire  _GEN_30226 = io_op_bits_active_vst ? _GEN_30048 : _GEN_28184; // @[sequencer-master.scala 654:38]
  wire  _GEN_30227 = io_op_bits_active_vst ? _GEN_30056 : _GEN_28185; // @[sequencer-master.scala 654:38]
  wire  _GEN_30228 = io_op_bits_active_vst ? _GEN_29420 : _GEN_28186; // @[sequencer-master.scala 654:38]
  wire  _GEN_30229 = io_op_bits_active_vst ? _GEN_29421 : _GEN_28187; // @[sequencer-master.scala 654:38]
  wire  _GEN_30230 = io_op_bits_active_vst ? _GEN_29422 : _GEN_28188; // @[sequencer-master.scala 654:38]
  wire  _GEN_30231 = io_op_bits_active_vst ? _GEN_29423 : _GEN_28189; // @[sequencer-master.scala 654:38]
  wire  _GEN_30232 = io_op_bits_active_vst ? _GEN_29424 : _GEN_28190; // @[sequencer-master.scala 654:38]
  wire  _GEN_30233 = io_op_bits_active_vst ? _GEN_29425 : _GEN_28191; // @[sequencer-master.scala 654:38]
  wire  _GEN_30234 = io_op_bits_active_vst ? _GEN_29426 : _GEN_28192; // @[sequencer-master.scala 654:38]
  wire  _GEN_30235 = io_op_bits_active_vst ? _GEN_29427 : _GEN_28193; // @[sequencer-master.scala 654:38]
  wire  _GEN_30236 = io_op_bits_active_vst ? _GEN_29428 : _GEN_28194; // @[sequencer-master.scala 654:38]
  wire  _GEN_30237 = io_op_bits_active_vst ? _GEN_29429 : _GEN_28195; // @[sequencer-master.scala 654:38]
  wire  _GEN_30238 = io_op_bits_active_vst ? _GEN_29430 : _GEN_28196; // @[sequencer-master.scala 654:38]
  wire  _GEN_30239 = io_op_bits_active_vst ? _GEN_29431 : _GEN_28197; // @[sequencer-master.scala 654:38]
  wire  _GEN_30240 = io_op_bits_active_vst ? _GEN_29432 : _GEN_28198; // @[sequencer-master.scala 654:38]
  wire  _GEN_30241 = io_op_bits_active_vst ? _GEN_29433 : _GEN_28199; // @[sequencer-master.scala 654:38]
  wire  _GEN_30242 = io_op_bits_active_vst ? _GEN_29434 : _GEN_28200; // @[sequencer-master.scala 654:38]
  wire  _GEN_30243 = io_op_bits_active_vst ? _GEN_29435 : _GEN_28201; // @[sequencer-master.scala 654:38]
  wire  _GEN_30244 = io_op_bits_active_vst ? _GEN_30001 : _GEN_28202; // @[sequencer-master.scala 654:38]
  wire  _GEN_30245 = io_op_bits_active_vst ? _GEN_30009 : _GEN_28203; // @[sequencer-master.scala 654:38]
  wire  _GEN_30246 = io_op_bits_active_vst ? _GEN_30017 : _GEN_28204; // @[sequencer-master.scala 654:38]
  wire  _GEN_30247 = io_op_bits_active_vst ? _GEN_30025 : _GEN_28205; // @[sequencer-master.scala 654:38]
  wire  _GEN_30248 = io_op_bits_active_vst ? _GEN_30033 : _GEN_28206; // @[sequencer-master.scala 654:38]
  wire  _GEN_30249 = io_op_bits_active_vst ? _GEN_30041 : _GEN_28207; // @[sequencer-master.scala 654:38]
  wire  _GEN_30250 = io_op_bits_active_vst ? _GEN_30049 : _GEN_28208; // @[sequencer-master.scala 654:38]
  wire  _GEN_30251 = io_op_bits_active_vst ? _GEN_30057 : _GEN_28209; // @[sequencer-master.scala 654:38]
  wire  _GEN_30252 = io_op_bits_active_vst ? _GEN_29444 : _GEN_28210; // @[sequencer-master.scala 654:38]
  wire  _GEN_30253 = io_op_bits_active_vst ? _GEN_29445 : _GEN_28211; // @[sequencer-master.scala 654:38]
  wire  _GEN_30254 = io_op_bits_active_vst ? _GEN_29446 : _GEN_28212; // @[sequencer-master.scala 654:38]
  wire  _GEN_30255 = io_op_bits_active_vst ? _GEN_29447 : _GEN_28213; // @[sequencer-master.scala 654:38]
  wire  _GEN_30256 = io_op_bits_active_vst ? _GEN_29448 : _GEN_28214; // @[sequencer-master.scala 654:38]
  wire  _GEN_30257 = io_op_bits_active_vst ? _GEN_29449 : _GEN_28215; // @[sequencer-master.scala 654:38]
  wire  _GEN_30258 = io_op_bits_active_vst ? _GEN_29450 : _GEN_28216; // @[sequencer-master.scala 654:38]
  wire  _GEN_30259 = io_op_bits_active_vst ? _GEN_29451 : _GEN_28217; // @[sequencer-master.scala 654:38]
  wire  _GEN_30260 = io_op_bits_active_vst ? _GEN_29452 : _GEN_28218; // @[sequencer-master.scala 654:38]
  wire  _GEN_30261 = io_op_bits_active_vst ? _GEN_29453 : _GEN_28219; // @[sequencer-master.scala 654:38]
  wire  _GEN_30262 = io_op_bits_active_vst ? _GEN_29454 : _GEN_28220; // @[sequencer-master.scala 654:38]
  wire  _GEN_30263 = io_op_bits_active_vst ? _GEN_29455 : _GEN_28221; // @[sequencer-master.scala 654:38]
  wire  _GEN_30264 = io_op_bits_active_vst ? _GEN_29456 : _GEN_28222; // @[sequencer-master.scala 654:38]
  wire  _GEN_30265 = io_op_bits_active_vst ? _GEN_29457 : _GEN_28223; // @[sequencer-master.scala 654:38]
  wire  _GEN_30266 = io_op_bits_active_vst ? _GEN_29458 : _GEN_28224; // @[sequencer-master.scala 654:38]
  wire  _GEN_30267 = io_op_bits_active_vst ? _GEN_29459 : _GEN_28225; // @[sequencer-master.scala 654:38]
  wire  _GEN_30268 = io_op_bits_active_vst ? _GEN_30002 : _GEN_28226; // @[sequencer-master.scala 654:38]
  wire  _GEN_30269 = io_op_bits_active_vst ? _GEN_30010 : _GEN_28227; // @[sequencer-master.scala 654:38]
  wire  _GEN_30270 = io_op_bits_active_vst ? _GEN_30018 : _GEN_28228; // @[sequencer-master.scala 654:38]
  wire  _GEN_30271 = io_op_bits_active_vst ? _GEN_30026 : _GEN_28229; // @[sequencer-master.scala 654:38]
  wire  _GEN_30272 = io_op_bits_active_vst ? _GEN_30034 : _GEN_28230; // @[sequencer-master.scala 654:38]
  wire  _GEN_30273 = io_op_bits_active_vst ? _GEN_30042 : _GEN_28231; // @[sequencer-master.scala 654:38]
  wire  _GEN_30274 = io_op_bits_active_vst ? _GEN_30050 : _GEN_28232; // @[sequencer-master.scala 654:38]
  wire  _GEN_30275 = io_op_bits_active_vst ? _GEN_30058 : _GEN_28233; // @[sequencer-master.scala 654:38]
  wire  _GEN_30276 = io_op_bits_active_vst ? _GEN_29468 : _GEN_28234; // @[sequencer-master.scala 654:38]
  wire  _GEN_30277 = io_op_bits_active_vst ? _GEN_29469 : _GEN_28235; // @[sequencer-master.scala 654:38]
  wire  _GEN_30278 = io_op_bits_active_vst ? _GEN_29470 : _GEN_28236; // @[sequencer-master.scala 654:38]
  wire  _GEN_30279 = io_op_bits_active_vst ? _GEN_29471 : _GEN_28237; // @[sequencer-master.scala 654:38]
  wire  _GEN_30280 = io_op_bits_active_vst ? _GEN_29472 : _GEN_28238; // @[sequencer-master.scala 654:38]
  wire  _GEN_30281 = io_op_bits_active_vst ? _GEN_29473 : _GEN_28239; // @[sequencer-master.scala 654:38]
  wire  _GEN_30282 = io_op_bits_active_vst ? _GEN_29474 : _GEN_28240; // @[sequencer-master.scala 654:38]
  wire  _GEN_30283 = io_op_bits_active_vst ? _GEN_29475 : _GEN_28241; // @[sequencer-master.scala 654:38]
  wire  _GEN_30284 = io_op_bits_active_vst ? _GEN_29476 : _GEN_28242; // @[sequencer-master.scala 654:38]
  wire  _GEN_30285 = io_op_bits_active_vst ? _GEN_29477 : _GEN_28243; // @[sequencer-master.scala 654:38]
  wire  _GEN_30286 = io_op_bits_active_vst ? _GEN_29478 : _GEN_28244; // @[sequencer-master.scala 654:38]
  wire  _GEN_30287 = io_op_bits_active_vst ? _GEN_29479 : _GEN_28245; // @[sequencer-master.scala 654:38]
  wire  _GEN_30288 = io_op_bits_active_vst ? _GEN_29480 : _GEN_28246; // @[sequencer-master.scala 654:38]
  wire  _GEN_30289 = io_op_bits_active_vst ? _GEN_29481 : _GEN_28247; // @[sequencer-master.scala 654:38]
  wire  _GEN_30290 = io_op_bits_active_vst ? _GEN_29482 : _GEN_28248; // @[sequencer-master.scala 654:38]
  wire  _GEN_30291 = io_op_bits_active_vst ? _GEN_29483 : _GEN_28249; // @[sequencer-master.scala 654:38]
  wire  _GEN_30292 = io_op_bits_active_vst ? _GEN_30003 : _GEN_28250; // @[sequencer-master.scala 654:38]
  wire  _GEN_30293 = io_op_bits_active_vst ? _GEN_30011 : _GEN_28251; // @[sequencer-master.scala 654:38]
  wire  _GEN_30294 = io_op_bits_active_vst ? _GEN_30019 : _GEN_28252; // @[sequencer-master.scala 654:38]
  wire  _GEN_30295 = io_op_bits_active_vst ? _GEN_30027 : _GEN_28253; // @[sequencer-master.scala 654:38]
  wire  _GEN_30296 = io_op_bits_active_vst ? _GEN_30035 : _GEN_28254; // @[sequencer-master.scala 654:38]
  wire  _GEN_30297 = io_op_bits_active_vst ? _GEN_30043 : _GEN_28255; // @[sequencer-master.scala 654:38]
  wire  _GEN_30298 = io_op_bits_active_vst ? _GEN_30051 : _GEN_28256; // @[sequencer-master.scala 654:38]
  wire  _GEN_30299 = io_op_bits_active_vst ? _GEN_30059 : _GEN_28257; // @[sequencer-master.scala 654:38]
  wire  _GEN_30300 = io_op_bits_active_vst ? _GEN_29492 : _GEN_28258; // @[sequencer-master.scala 654:38]
  wire  _GEN_30301 = io_op_bits_active_vst ? _GEN_29493 : _GEN_28259; // @[sequencer-master.scala 654:38]
  wire  _GEN_30302 = io_op_bits_active_vst ? _GEN_29494 : _GEN_28260; // @[sequencer-master.scala 654:38]
  wire  _GEN_30303 = io_op_bits_active_vst ? _GEN_29495 : _GEN_28261; // @[sequencer-master.scala 654:38]
  wire  _GEN_30304 = io_op_bits_active_vst ? _GEN_29496 : _GEN_28262; // @[sequencer-master.scala 654:38]
  wire  _GEN_30305 = io_op_bits_active_vst ? _GEN_29497 : _GEN_28263; // @[sequencer-master.scala 654:38]
  wire  _GEN_30306 = io_op_bits_active_vst ? _GEN_29498 : _GEN_28264; // @[sequencer-master.scala 654:38]
  wire  _GEN_30307 = io_op_bits_active_vst ? _GEN_29499 : _GEN_28265; // @[sequencer-master.scala 654:38]
  wire  _GEN_30308 = io_op_bits_active_vst ? _GEN_29500 : _GEN_28266; // @[sequencer-master.scala 654:38]
  wire  _GEN_30309 = io_op_bits_active_vst ? _GEN_29501 : _GEN_28267; // @[sequencer-master.scala 654:38]
  wire  _GEN_30310 = io_op_bits_active_vst ? _GEN_29502 : _GEN_28268; // @[sequencer-master.scala 654:38]
  wire  _GEN_30311 = io_op_bits_active_vst ? _GEN_29503 : _GEN_28269; // @[sequencer-master.scala 654:38]
  wire  _GEN_30312 = io_op_bits_active_vst ? _GEN_29504 : _GEN_28270; // @[sequencer-master.scala 654:38]
  wire  _GEN_30313 = io_op_bits_active_vst ? _GEN_29505 : _GEN_28271; // @[sequencer-master.scala 654:38]
  wire  _GEN_30314 = io_op_bits_active_vst ? _GEN_29506 : _GEN_28272; // @[sequencer-master.scala 654:38]
  wire  _GEN_30315 = io_op_bits_active_vst ? _GEN_29507 : _GEN_28273; // @[sequencer-master.scala 654:38]
  wire  _GEN_30316 = io_op_bits_active_vst ? _GEN_29508 : _GEN_28274; // @[sequencer-master.scala 654:38]
  wire  _GEN_30317 = io_op_bits_active_vst ? _GEN_29509 : _GEN_28275; // @[sequencer-master.scala 654:38]
  wire  _GEN_30318 = io_op_bits_active_vst ? _GEN_29510 : _GEN_28276; // @[sequencer-master.scala 654:38]
  wire  _GEN_30319 = io_op_bits_active_vst ? _GEN_29511 : _GEN_28277; // @[sequencer-master.scala 654:38]
  wire  _GEN_30320 = io_op_bits_active_vst ? _GEN_29512 : _GEN_28278; // @[sequencer-master.scala 654:38]
  wire  _GEN_30321 = io_op_bits_active_vst ? _GEN_29513 : _GEN_28279; // @[sequencer-master.scala 654:38]
  wire  _GEN_30322 = io_op_bits_active_vst ? _GEN_29514 : _GEN_28280; // @[sequencer-master.scala 654:38]
  wire  _GEN_30323 = io_op_bits_active_vst ? _GEN_29515 : _GEN_28281; // @[sequencer-master.scala 654:38]
  wire  _GEN_30332 = io_op_bits_active_vst ? _GEN_28692 : _GEN_28290; // @[sequencer-master.scala 654:38]
  wire  _GEN_30333 = io_op_bits_active_vst ? _GEN_28693 : _GEN_28291; // @[sequencer-master.scala 654:38]
  wire  _GEN_30334 = io_op_bits_active_vst ? _GEN_28694 : _GEN_28292; // @[sequencer-master.scala 654:38]
  wire  _GEN_30335 = io_op_bits_active_vst ? _GEN_28695 : _GEN_28293; // @[sequencer-master.scala 654:38]
  wire  _GEN_30336 = io_op_bits_active_vst ? _GEN_28696 : _GEN_28294; // @[sequencer-master.scala 654:38]
  wire  _GEN_30337 = io_op_bits_active_vst ? _GEN_28697 : _GEN_28295; // @[sequencer-master.scala 654:38]
  wire  _GEN_30338 = io_op_bits_active_vst ? _GEN_28698 : _GEN_28296; // @[sequencer-master.scala 654:38]
  wire  _GEN_30339 = io_op_bits_active_vst ? _GEN_28699 : _GEN_28297; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30372 = io_op_bits_active_vst ? _GEN_29612 : _GEN_28330; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30373 = io_op_bits_active_vst ? _GEN_29613 : _GEN_28331; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30374 = io_op_bits_active_vst ? _GEN_29614 : _GEN_28332; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30375 = io_op_bits_active_vst ? _GEN_29615 : _GEN_28333; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30376 = io_op_bits_active_vst ? _GEN_29616 : _GEN_28334; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30377 = io_op_bits_active_vst ? _GEN_29617 : _GEN_28335; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30378 = io_op_bits_active_vst ? _GEN_29618 : _GEN_28336; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30379 = io_op_bits_active_vst ? _GEN_29619 : _GEN_28337; // @[sequencer-master.scala 654:38]
  wire  _GEN_30404 = io_op_bits_active_vst ? _GEN_29212 : _GEN_28362; // @[sequencer-master.scala 654:38]
  wire  _GEN_30405 = io_op_bits_active_vst ? _GEN_29213 : _GEN_28363; // @[sequencer-master.scala 654:38]
  wire  _GEN_30406 = io_op_bits_active_vst ? _GEN_29214 : _GEN_28364; // @[sequencer-master.scala 654:38]
  wire  _GEN_30407 = io_op_bits_active_vst ? _GEN_29215 : _GEN_28365; // @[sequencer-master.scala 654:38]
  wire  _GEN_30408 = io_op_bits_active_vst ? _GEN_29216 : _GEN_28366; // @[sequencer-master.scala 654:38]
  wire  _GEN_30409 = io_op_bits_active_vst ? _GEN_29217 : _GEN_28367; // @[sequencer-master.scala 654:38]
  wire  _GEN_30410 = io_op_bits_active_vst ? _GEN_29218 : _GEN_28368; // @[sequencer-master.scala 654:38]
  wire  _GEN_30411 = io_op_bits_active_vst ? _GEN_29219 : _GEN_28369; // @[sequencer-master.scala 654:38]
  wire  _GEN_30412 = io_op_bits_active_vst ? _GEN_29524 : _GEN_26256; // @[sequencer-master.scala 654:38]
  wire  _GEN_30413 = io_op_bits_active_vst ? _GEN_29525 : _GEN_26257; // @[sequencer-master.scala 654:38]
  wire  _GEN_30414 = io_op_bits_active_vst ? _GEN_29526 : _GEN_26258; // @[sequencer-master.scala 654:38]
  wire  _GEN_30415 = io_op_bits_active_vst ? _GEN_29527 : _GEN_26259; // @[sequencer-master.scala 654:38]
  wire  _GEN_30416 = io_op_bits_active_vst ? _GEN_29528 : _GEN_26260; // @[sequencer-master.scala 654:38]
  wire  _GEN_30417 = io_op_bits_active_vst ? _GEN_29529 : _GEN_26261; // @[sequencer-master.scala 654:38]
  wire  _GEN_30418 = io_op_bits_active_vst ? _GEN_29530 : _GEN_26262; // @[sequencer-master.scala 654:38]
  wire  _GEN_30419 = io_op_bits_active_vst ? _GEN_29531 : _GEN_26263; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30452 = io_op_bits_active_vst ? _GEN_29836 : _GEN_26208; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30453 = io_op_bits_active_vst ? _GEN_29837 : _GEN_26209; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30454 = io_op_bits_active_vst ? _GEN_29838 : _GEN_26210; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30455 = io_op_bits_active_vst ? _GEN_29839 : _GEN_26211; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30456 = io_op_bits_active_vst ? _GEN_29840 : _GEN_26212; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30457 = io_op_bits_active_vst ? _GEN_29841 : _GEN_26213; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30458 = io_op_bits_active_vst ? _GEN_29842 : _GEN_26214; // @[sequencer-master.scala 654:38]
  wire [7:0] _GEN_30459 = io_op_bits_active_vst ? _GEN_29843 : _GEN_26215; // @[sequencer-master.scala 654:38]
  wire  _GEN_30460 = io_op_bits_active_vst | _GEN_28418; // @[sequencer-master.scala 654:38 sequencer-master.scala 265:41]
  wire  _GEN_30462 = _T_1752 ? _GEN_30060 : v_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30463 = _T_1752 ? _GEN_30061 : v_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30464 = _T_1752 ? _GEN_30062 : v_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30465 = _T_1752 ? _GEN_30063 : v_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30466 = _T_1752 ? _GEN_30064 : v_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30467 = _T_1752 ? _GEN_30065 : v_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30468 = _T_1752 ? _GEN_30066 : v_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30469 = _T_1752 ? _GEN_30067 : v_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 107:14]
  wire  _GEN_30518 = _T_1752 & _GEN_30116; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30519 = _T_1752 & _GEN_30117; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30520 = _T_1752 & _GEN_30118; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30521 = _T_1752 & _GEN_30119; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30522 = _T_1752 & _GEN_30120; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30523 = _T_1752 & _GEN_30121; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30524 = _T_1752 & _GEN_30122; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30525 = _T_1752 & _GEN_30123; // @[sequencer-master.scala 639:27 sequencer-master.scala 192:24]
  wire  _GEN_30526 = _T_1752 ? _GEN_30124 : e_0_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30527 = _T_1752 ? _GEN_30125 : e_1_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30528 = _T_1752 ? _GEN_30126 : e_2_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30529 = _T_1752 ? _GEN_30127 : e_3_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30530 = _T_1752 ? _GEN_30128 : e_4_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30531 = _T_1752 ? _GEN_30129 : e_5_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30532 = _T_1752 ? _GEN_30130 : e_6_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30533 = _T_1752 ? _GEN_30131 : e_7_raw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30534 = _T_1752 ? _GEN_30132 : e_0_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30535 = _T_1752 ? _GEN_30133 : e_1_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30536 = _T_1752 ? _GEN_30134 : e_2_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30537 = _T_1752 ? _GEN_30135 : e_3_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30538 = _T_1752 ? _GEN_30136 : e_4_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30539 = _T_1752 ? _GEN_30137 : e_5_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30540 = _T_1752 ? _GEN_30138 : e_6_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30541 = _T_1752 ? _GEN_30139 : e_7_war_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30542 = _T_1752 ? _GEN_30140 : e_0_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30543 = _T_1752 ? _GEN_30141 : e_1_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30544 = _T_1752 ? _GEN_30142 : e_2_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30545 = _T_1752 ? _GEN_30143 : e_3_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30546 = _T_1752 ? _GEN_30144 : e_4_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30547 = _T_1752 ? _GEN_30145 : e_5_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30548 = _T_1752 ? _GEN_30146 : e_6_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30549 = _T_1752 ? _GEN_30147 : e_7_waw_0; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30550 = _T_1752 ? _GEN_30148 : e_0_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30551 = _T_1752 ? _GEN_30149 : e_1_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30552 = _T_1752 ? _GEN_30150 : e_2_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30553 = _T_1752 ? _GEN_30151 : e_3_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30554 = _T_1752 ? _GEN_30152 : e_4_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30555 = _T_1752 ? _GEN_30153 : e_5_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30556 = _T_1752 ? _GEN_30154 : e_6_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30557 = _T_1752 ? _GEN_30155 : e_7_raw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30558 = _T_1752 ? _GEN_30156 : e_0_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30559 = _T_1752 ? _GEN_30157 : e_1_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30560 = _T_1752 ? _GEN_30158 : e_2_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30561 = _T_1752 ? _GEN_30159 : e_3_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30562 = _T_1752 ? _GEN_30160 : e_4_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30563 = _T_1752 ? _GEN_30161 : e_5_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30564 = _T_1752 ? _GEN_30162 : e_6_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30565 = _T_1752 ? _GEN_30163 : e_7_war_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30566 = _T_1752 ? _GEN_30164 : e_0_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30567 = _T_1752 ? _GEN_30165 : e_1_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30568 = _T_1752 ? _GEN_30166 : e_2_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30569 = _T_1752 ? _GEN_30167 : e_3_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30570 = _T_1752 ? _GEN_30168 : e_4_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30571 = _T_1752 ? _GEN_30169 : e_5_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30572 = _T_1752 ? _GEN_30170 : e_6_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30573 = _T_1752 ? _GEN_30171 : e_7_waw_1; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30574 = _T_1752 ? _GEN_30172 : e_0_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30575 = _T_1752 ? _GEN_30173 : e_1_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30576 = _T_1752 ? _GEN_30174 : e_2_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30577 = _T_1752 ? _GEN_30175 : e_3_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30578 = _T_1752 ? _GEN_30176 : e_4_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30579 = _T_1752 ? _GEN_30177 : e_5_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30580 = _T_1752 ? _GEN_30178 : e_6_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30581 = _T_1752 ? _GEN_30179 : e_7_raw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30582 = _T_1752 ? _GEN_30180 : e_0_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30583 = _T_1752 ? _GEN_30181 : e_1_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30584 = _T_1752 ? _GEN_30182 : e_2_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30585 = _T_1752 ? _GEN_30183 : e_3_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30586 = _T_1752 ? _GEN_30184 : e_4_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30587 = _T_1752 ? _GEN_30185 : e_5_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30588 = _T_1752 ? _GEN_30186 : e_6_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30589 = _T_1752 ? _GEN_30187 : e_7_war_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30590 = _T_1752 ? _GEN_30188 : e_0_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30591 = _T_1752 ? _GEN_30189 : e_1_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30592 = _T_1752 ? _GEN_30190 : e_2_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30593 = _T_1752 ? _GEN_30191 : e_3_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30594 = _T_1752 ? _GEN_30192 : e_4_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30595 = _T_1752 ? _GEN_30193 : e_5_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30596 = _T_1752 ? _GEN_30194 : e_6_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30597 = _T_1752 ? _GEN_30195 : e_7_waw_2; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30598 = _T_1752 ? _GEN_30196 : e_0_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30599 = _T_1752 ? _GEN_30197 : e_1_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30600 = _T_1752 ? _GEN_30198 : e_2_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30601 = _T_1752 ? _GEN_30199 : e_3_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30602 = _T_1752 ? _GEN_30200 : e_4_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30603 = _T_1752 ? _GEN_30201 : e_5_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30604 = _T_1752 ? _GEN_30202 : e_6_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30605 = _T_1752 ? _GEN_30203 : e_7_raw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30606 = _T_1752 ? _GEN_30204 : e_0_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30607 = _T_1752 ? _GEN_30205 : e_1_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30608 = _T_1752 ? _GEN_30206 : e_2_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30609 = _T_1752 ? _GEN_30207 : e_3_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30610 = _T_1752 ? _GEN_30208 : e_4_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30611 = _T_1752 ? _GEN_30209 : e_5_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30612 = _T_1752 ? _GEN_30210 : e_6_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30613 = _T_1752 ? _GEN_30211 : e_7_war_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30614 = _T_1752 ? _GEN_30212 : e_0_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30615 = _T_1752 ? _GEN_30213 : e_1_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30616 = _T_1752 ? _GEN_30214 : e_2_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30617 = _T_1752 ? _GEN_30215 : e_3_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30618 = _T_1752 ? _GEN_30216 : e_4_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30619 = _T_1752 ? _GEN_30217 : e_5_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30620 = _T_1752 ? _GEN_30218 : e_6_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30621 = _T_1752 ? _GEN_30219 : e_7_waw_3; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30622 = _T_1752 ? _GEN_30220 : e_0_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30623 = _T_1752 ? _GEN_30221 : e_1_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30624 = _T_1752 ? _GEN_30222 : e_2_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30625 = _T_1752 ? _GEN_30223 : e_3_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30626 = _T_1752 ? _GEN_30224 : e_4_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30627 = _T_1752 ? _GEN_30225 : e_5_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30628 = _T_1752 ? _GEN_30226 : e_6_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30629 = _T_1752 ? _GEN_30227 : e_7_raw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30630 = _T_1752 ? _GEN_30228 : e_0_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30631 = _T_1752 ? _GEN_30229 : e_1_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30632 = _T_1752 ? _GEN_30230 : e_2_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30633 = _T_1752 ? _GEN_30231 : e_3_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30634 = _T_1752 ? _GEN_30232 : e_4_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30635 = _T_1752 ? _GEN_30233 : e_5_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30636 = _T_1752 ? _GEN_30234 : e_6_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30637 = _T_1752 ? _GEN_30235 : e_7_war_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30638 = _T_1752 ? _GEN_30236 : e_0_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30639 = _T_1752 ? _GEN_30237 : e_1_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30640 = _T_1752 ? _GEN_30238 : e_2_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30641 = _T_1752 ? _GEN_30239 : e_3_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30642 = _T_1752 ? _GEN_30240 : e_4_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30643 = _T_1752 ? _GEN_30241 : e_5_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30644 = _T_1752 ? _GEN_30242 : e_6_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30645 = _T_1752 ? _GEN_30243 : e_7_waw_4; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30646 = _T_1752 ? _GEN_30244 : e_0_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30647 = _T_1752 ? _GEN_30245 : e_1_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30648 = _T_1752 ? _GEN_30246 : e_2_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30649 = _T_1752 ? _GEN_30247 : e_3_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30650 = _T_1752 ? _GEN_30248 : e_4_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30651 = _T_1752 ? _GEN_30249 : e_5_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30652 = _T_1752 ? _GEN_30250 : e_6_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30653 = _T_1752 ? _GEN_30251 : e_7_raw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30654 = _T_1752 ? _GEN_30252 : e_0_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30655 = _T_1752 ? _GEN_30253 : e_1_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30656 = _T_1752 ? _GEN_30254 : e_2_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30657 = _T_1752 ? _GEN_30255 : e_3_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30658 = _T_1752 ? _GEN_30256 : e_4_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30659 = _T_1752 ? _GEN_30257 : e_5_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30660 = _T_1752 ? _GEN_30258 : e_6_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30661 = _T_1752 ? _GEN_30259 : e_7_war_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30662 = _T_1752 ? _GEN_30260 : e_0_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30663 = _T_1752 ? _GEN_30261 : e_1_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30664 = _T_1752 ? _GEN_30262 : e_2_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30665 = _T_1752 ? _GEN_30263 : e_3_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30666 = _T_1752 ? _GEN_30264 : e_4_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30667 = _T_1752 ? _GEN_30265 : e_5_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30668 = _T_1752 ? _GEN_30266 : e_6_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30669 = _T_1752 ? _GEN_30267 : e_7_waw_5; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30670 = _T_1752 ? _GEN_30268 : e_0_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30671 = _T_1752 ? _GEN_30269 : e_1_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30672 = _T_1752 ? _GEN_30270 : e_2_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30673 = _T_1752 ? _GEN_30271 : e_3_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30674 = _T_1752 ? _GEN_30272 : e_4_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30675 = _T_1752 ? _GEN_30273 : e_5_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30676 = _T_1752 ? _GEN_30274 : e_6_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30677 = _T_1752 ? _GEN_30275 : e_7_raw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30678 = _T_1752 ? _GEN_30276 : e_0_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30679 = _T_1752 ? _GEN_30277 : e_1_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30680 = _T_1752 ? _GEN_30278 : e_2_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30681 = _T_1752 ? _GEN_30279 : e_3_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30682 = _T_1752 ? _GEN_30280 : e_4_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30683 = _T_1752 ? _GEN_30281 : e_5_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30684 = _T_1752 ? _GEN_30282 : e_6_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30685 = _T_1752 ? _GEN_30283 : e_7_war_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30686 = _T_1752 ? _GEN_30284 : e_0_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30687 = _T_1752 ? _GEN_30285 : e_1_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30688 = _T_1752 ? _GEN_30286 : e_2_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30689 = _T_1752 ? _GEN_30287 : e_3_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30690 = _T_1752 ? _GEN_30288 : e_4_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30691 = _T_1752 ? _GEN_30289 : e_5_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30692 = _T_1752 ? _GEN_30290 : e_6_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30693 = _T_1752 ? _GEN_30291 : e_7_waw_6; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30694 = _T_1752 ? _GEN_30292 : e_0_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30695 = _T_1752 ? _GEN_30293 : e_1_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30696 = _T_1752 ? _GEN_30294 : e_2_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30697 = _T_1752 ? _GEN_30295 : e_3_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30698 = _T_1752 ? _GEN_30296 : e_4_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30699 = _T_1752 ? _GEN_30297 : e_5_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30700 = _T_1752 ? _GEN_30298 : e_6_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30701 = _T_1752 ? _GEN_30299 : e_7_raw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 194:26]
  wire  _GEN_30702 = _T_1752 ? _GEN_30300 : e_0_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30703 = _T_1752 ? _GEN_30301 : e_1_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30704 = _T_1752 ? _GEN_30302 : e_2_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30705 = _T_1752 ? _GEN_30303 : e_3_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30706 = _T_1752 ? _GEN_30304 : e_4_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30707 = _T_1752 ? _GEN_30305 : e_5_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30708 = _T_1752 ? _GEN_30306 : e_6_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30709 = _T_1752 ? _GEN_30307 : e_7_war_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 195:26]
  wire  _GEN_30710 = _T_1752 ? _GEN_30308 : e_0_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30711 = _T_1752 ? _GEN_30309 : e_1_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30712 = _T_1752 ? _GEN_30310 : e_2_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30713 = _T_1752 ? _GEN_30311 : e_3_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30714 = _T_1752 ? _GEN_30312 : e_4_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30715 = _T_1752 ? _GEN_30313 : e_5_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30716 = _T_1752 ? _GEN_30314 : e_6_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30717 = _T_1752 ? _GEN_30315 : e_7_waw_7; // @[sequencer-master.scala 639:27 sequencer-master.scala 196:26]
  wire  _GEN_30718 = _T_1752 ? _GEN_30316 : e_0_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30719 = _T_1752 ? _GEN_30317 : e_1_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30720 = _T_1752 ? _GEN_30318 : e_2_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30721 = _T_1752 ? _GEN_30319 : e_3_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30722 = _T_1752 ? _GEN_30320 : e_4_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30723 = _T_1752 ? _GEN_30321 : e_5_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30724 = _T_1752 ? _GEN_30322 : e_6_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30725 = _T_1752 ? _GEN_30323 : e_7_last; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30734 = _T_1752 ? _GEN_1672 : e_0_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30735 = _T_1752 ? _GEN_1673 : e_1_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30736 = _T_1752 ? _GEN_1674 : e_2_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30737 = _T_1752 ? _GEN_1675 : e_3_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30738 = _T_1752 ? _GEN_1676 : e_4_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30739 = _T_1752 ? _GEN_1677 : e_5_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30740 = _T_1752 ? _GEN_1678 : e_6_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30741 = _T_1752 ? _GEN_1679 : e_7_active_viu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30942 = _T_1752 & _GEN_30460; // @[sequencer-master.scala 639:27 sequencer-master.scala 405:19]
  wire  _GEN_30944 = _T_1752 ? _GEN_3594 : e_0_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30945 = _T_1752 ? _GEN_3595 : e_1_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30946 = _T_1752 ? _GEN_3596 : e_2_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30947 = _T_1752 ? _GEN_3597 : e_3_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30948 = _T_1752 ? _GEN_3598 : e_4_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30949 = _T_1752 ? _GEN_3599 : e_5_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30950 = _T_1752 ? _GEN_3600 : e_6_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_30951 = _T_1752 ? _GEN_3601 : e_7_active_vipu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31000 = _T_1752 ? _GEN_5492 : e_0_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31001 = _T_1752 ? _GEN_5493 : e_1_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31002 = _T_1752 ? _GEN_5494 : e_2_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31003 = _T_1752 ? _GEN_5495 : e_3_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31004 = _T_1752 ? _GEN_5496 : e_4_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31005 = _T_1752 ? _GEN_5497 : e_5_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31006 = _T_1752 ? _GEN_5498 : e_6_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31007 = _T_1752 ? _GEN_5499 : e_7_active_vimu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31008 = _T_1752 ? _GEN_18106 : e_0_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31009 = _T_1752 ? _GEN_18107 : e_1_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31010 = _T_1752 ? _GEN_18108 : e_2_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31011 = _T_1752 ? _GEN_18109 : e_3_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31012 = _T_1752 ? _GEN_18110 : e_4_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31013 = _T_1752 ? _GEN_18111 : e_5_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31014 = _T_1752 ? _GEN_18112 : e_6_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31015 = _T_1752 ? _GEN_18113 : e_7_active_vqu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31016 = _T_1752 ? _GEN_8078 : e_0_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31017 = _T_1752 ? _GEN_8079 : e_1_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31018 = _T_1752 ? _GEN_8080 : e_2_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31019 = _T_1752 ? _GEN_8081 : e_3_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31020 = _T_1752 ? _GEN_8082 : e_4_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31021 = _T_1752 ? _GEN_8083 : e_5_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31022 = _T_1752 ? _GEN_8084 : e_6_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31023 = _T_1752 ? _GEN_8085 : e_7_active_vidu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31024 = _T_1752 ? _GEN_10048 : e_0_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31025 = _T_1752 ? _GEN_10049 : e_1_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31026 = _T_1752 ? _GEN_10050 : e_2_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31027 = _T_1752 ? _GEN_10051 : e_3_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31028 = _T_1752 ? _GEN_10052 : e_4_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31029 = _T_1752 ? _GEN_10053 : e_5_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31030 = _T_1752 ? _GEN_10054 : e_6_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31031 = _T_1752 ? _GEN_10055 : e_7_active_vfmu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31032 = _T_1752 ? _GEN_12682 : e_0_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31033 = _T_1752 ? _GEN_12683 : e_1_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31034 = _T_1752 ? _GEN_12684 : e_2_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31035 = _T_1752 ? _GEN_12685 : e_3_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31036 = _T_1752 ? _GEN_12686 : e_4_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31037 = _T_1752 ? _GEN_12687 : e_5_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31038 = _T_1752 ? _GEN_12688 : e_6_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31039 = _T_1752 ? _GEN_12689 : e_7_active_vfdu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31040 = _T_1752 ? _GEN_14404 : e_0_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31041 = _T_1752 ? _GEN_14405 : e_1_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31042 = _T_1752 ? _GEN_14406 : e_2_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31043 = _T_1752 ? _GEN_14407 : e_3_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31044 = _T_1752 ? _GEN_14408 : e_4_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31045 = _T_1752 ? _GEN_14409 : e_5_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31046 = _T_1752 ? _GEN_14410 : e_6_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31047 = _T_1752 ? _GEN_14411 : e_7_active_vfcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31048 = _T_1752 ? _GEN_16038 : e_0_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31049 = _T_1752 ? _GEN_16039 : e_1_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31050 = _T_1752 ? _GEN_16040 : e_2_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31051 = _T_1752 ? _GEN_16041 : e_3_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31052 = _T_1752 ? _GEN_16042 : e_4_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31053 = _T_1752 ? _GEN_16043 : e_5_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31054 = _T_1752 ? _GEN_16044 : e_6_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31055 = _T_1752 ? _GEN_16045 : e_7_active_vfvu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31056 = _T_1752 ? _GEN_26128 : e_0_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31057 = _T_1752 ? _GEN_26129 : e_1_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31058 = _T_1752 ? _GEN_26130 : e_2_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31059 = _T_1752 ? _GEN_26131 : e_3_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31060 = _T_1752 ? _GEN_26132 : e_4_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31061 = _T_1752 ? _GEN_26133 : e_5_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31062 = _T_1752 ? _GEN_26134 : e_6_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31063 = _T_1752 ? _GEN_26135 : e_7_active_vgu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31064 = _T_1752 ? _GEN_30404 : e_0_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31065 = _T_1752 ? _GEN_30405 : e_1_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31066 = _T_1752 ? _GEN_30406 : e_2_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31067 = _T_1752 ? _GEN_30407 : e_3_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31068 = _T_1752 ? _GEN_30408 : e_4_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31069 = _T_1752 ? _GEN_30409 : e_5_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31070 = _T_1752 ? _GEN_30410 : e_6_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31071 = _T_1752 ? _GEN_30411 : e_7_active_vcu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31072 = _T_1752 ? _GEN_30412 : e_0_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31073 = _T_1752 ? _GEN_30413 : e_1_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31074 = _T_1752 ? _GEN_30414 : e_2_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31075 = _T_1752 ? _GEN_30415 : e_3_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31076 = _T_1752 ? _GEN_30416 : e_4_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31077 = _T_1752 ? _GEN_30417 : e_5_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31078 = _T_1752 ? _GEN_30418 : e_6_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31079 = _T_1752 ? _GEN_30419 : e_7_active_vsu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31080 = _T_1752 ? _GEN_28370 : e_0_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31081 = _T_1752 ? _GEN_28371 : e_1_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31082 = _T_1752 ? _GEN_28372 : e_2_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31083 = _T_1752 ? _GEN_28373 : e_3_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31084 = _T_1752 ? _GEN_28374 : e_4_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31085 = _T_1752 ? _GEN_28375 : e_5_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31086 = _T_1752 ? _GEN_28376 : e_6_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31087 = _T_1752 ? _GEN_28377 : e_7_active_vlu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31088 = _T_1752 ? _GEN_30332 : e_0_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31089 = _T_1752 ? _GEN_30333 : e_1_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31090 = _T_1752 ? _GEN_30334 : e_2_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31091 = _T_1752 ? _GEN_30335 : e_3_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31092 = _T_1752 ? _GEN_30336 : e_4_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31093 = _T_1752 ? _GEN_30337 : e_5_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31094 = _T_1752 ? _GEN_30338 : e_6_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _GEN_31095 = _T_1752 ? _GEN_30339 : e_7_active_vpu; // @[sequencer-master.scala 639:27 sequencer-master.scala 109:14]
  wire  _T_2411 = ~maybe_full & head == tail; // @[sequencer-master.scala 389:27]
  wire [2:0] _T_2413 = head - tail; // @[sequencer-master.scala 389:52]
  wire [3:0] _T_2414 = {_T_2411,_T_2413}; // @[Cat.scala 30:58]
  wire  _T_2426 = _T_2414 >= 4'h2 & _T_1884; // @[sequencer-master.scala 398:26]
  wire  _T_2427 = _T_2414 >= 4'h1 & (io_op_bits_active_vint | io_op_bits_active_vipred | io_op_bits_active_vimul |
    io_op_bits_active_vfma | io_op_bits_active_vfcmp | io_op_bits_active_vfconv | io_op_bits_active_vrpred |
    io_op_bits_active_vrfirst) | _T_2426; // @[sequencer-master.scala 397:119]
  wire  _T_2432 = _T_2414 >= 4'h3 & (io_op_bits_active_vld | io_op_bits_active_vst | io_op_bits_active_vldx |
    io_op_bits_active_vstx); // @[sequencer-master.scala 399:26]
  wire  _T_2433 = _T_2427 | _T_2432; // @[sequencer-master.scala 398:50]
  wire  _T_2435 = _T_2414 >= 4'h4 & io_op_bits_active_vamo; // @[sequencer-master.scala 400:26]
  wire  _GEN_31097 = _GEN_30942 | maybe_full; // @[sequencer-master.scala 418:26 sequencer-master.scala 420:20 sequencer-master.scala 111:23]
  wire  _GEN_31118 = 3'h1 == head ? v_1 : v_0; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31119 = 3'h2 == head ? v_2 : _GEN_31118; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31120 = 3'h3 == head ? v_3 : _GEN_31119; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31121 = 3'h4 == head ? v_4 : _GEN_31120; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31122 = 3'h5 == head ? v_5 : _GEN_31121; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31123 = 3'h6 == head ? v_6 : _GEN_31122; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31124 = 3'h7 == head ? v_7 : _GEN_31123; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31126 = 3'h1 == head ? io_master_clear_1 : io_master_clear_0; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31127 = 3'h2 == head ? io_master_clear_2 : _GEN_31126; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31128 = 3'h3 == head ? io_master_clear_3 : _GEN_31127; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31129 = 3'h4 == head ? io_master_clear_4 : _GEN_31128; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31130 = 3'h5 == head ? io_master_clear_5 : _GEN_31129; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31131 = 3'h6 == head ? io_master_clear_6 : _GEN_31130; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _GEN_31132 = 3'h7 == head ? io_master_clear_7 : _GEN_31131; // @[sequencer-master.scala 438:21 sequencer-master.scala 438:21]
  wire  _T_2443 = _GEN_31124 & _GEN_31132; // @[sequencer-master.scala 438:21]
  wire [2:0] _T_2440 = head + 3'h1; // @[util.scala 94:11]
  wire [2:0] _T_2438 = tail + 3'h7; // @[util.scala 94:11]
  wire  _GEN_31100 = 3'h0 == _T_2438 | _GEN_30718; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31101 = 3'h1 == _T_2438 | _GEN_30719; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31102 = 3'h2 == _T_2438 | _GEN_30720; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31103 = 3'h3 == _T_2438 | _GEN_30721; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31104 = 3'h4 == _T_2438 | _GEN_30722; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31105 = 3'h5 == _T_2438 | _GEN_30723; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31106 = 3'h6 == _T_2438 | _GEN_30724; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31107 = 3'h7 == _T_2438 | _GEN_30725; // @[sequencer-master.scala 293:19 sequencer-master.scala 293:19]
  wire  _GEN_31116 = io_vf_stop & ~io_pending_all; // @[sequencer-master.scala 433:25 sequencer-master.scala 435:17 sequencer-master.scala 432:15]
  wire  _GEN_31603 = 3'h1 == head ? e_1_last : e_0_last; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_31676 = 3'h2 == head ? e_2_last : _GEN_31603; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_31749 = 3'h3 == head ? e_3_last : _GEN_31676; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_31822 = 3'h4 == head ? e_4_last : _GEN_31749; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_31895 = 3'h5 == head ? e_5_last : _GEN_31822; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_31968 = 3'h6 == head ? e_6_last : _GEN_31895; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_32041 = 3'h7 == head ? e_7_last : _GEN_31968; // @[sequencer-master.scala 441:33 sequencer-master.scala 441:33]
  wire  _GEN_32181 = _GEN_31124 & _GEN_31132 | _GEN_30518; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32206 = _GEN_31124 & _GEN_31132 | _GEN_30519; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32231 = _GEN_31124 & _GEN_31132 | _GEN_30520; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32256 = _GEN_31124 & _GEN_31132 | _GEN_30521; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32281 = _GEN_31124 & _GEN_31132 | _GEN_30522; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32306 = _GEN_31124 & _GEN_31132 | _GEN_30523; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32331 = _GEN_31124 & _GEN_31132 | _GEN_30524; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  wire  _GEN_32356 = _GEN_31124 & _GEN_31132 | _GEN_30525; // @[sequencer-master.scala 438:47 sequencer-master.scala 188:42]
  reg  _T_2465; // @[sequencer-master.scala 444:24]
  wire  _T_2466 = v_0 & e_0_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2467 = v_1 & e_1_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2468 = v_2 & e_2_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2469 = v_3 & e_3_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2470 = v_4 & e_4_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2471 = v_5 & e_5_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2472 = v_6 & e_6_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2473 = v_7 & e_7_active_vcu; // @[sequencer-master.scala 446:59]
  wire  _T_2479 = _T_2466 | _T_2467 | _T_2468 | _T_2469 | _T_2470 | _T_2471 | _T_2472; // @[sequencer-master.scala 447:39]
  wire  _T_2486 = v_0 | v_1 | v_2 | v_3 | v_4 | v_5 | v_6; // @[sequencer-master.scala 448:36]
  wire  _T_2490 = e_0_active_vgu | e_0_active_vcu | e_0_active_vlu | e_0_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2491 = v_0 & _T_2490; // @[sequencer-master.scala 451:34]
  wire  _T_2494 = e_1_active_vgu | e_1_active_vcu | e_1_active_vlu | e_1_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2495 = v_1 & _T_2494; // @[sequencer-master.scala 451:34]
  wire  _T_2498 = e_2_active_vgu | e_2_active_vcu | e_2_active_vlu | e_2_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2499 = v_2 & _T_2498; // @[sequencer-master.scala 451:34]
  wire  _T_2502 = e_3_active_vgu | e_3_active_vcu | e_3_active_vlu | e_3_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2503 = v_3 & _T_2502; // @[sequencer-master.scala 451:34]
  wire  _T_2506 = e_4_active_vgu | e_4_active_vcu | e_4_active_vlu | e_4_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2507 = v_4 & _T_2506; // @[sequencer-master.scala 451:34]
  wire  _T_2510 = e_5_active_vgu | e_5_active_vcu | e_5_active_vlu | e_5_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2511 = v_5 & _T_2510; // @[sequencer-master.scala 451:34]
  wire  _T_2514 = e_6_active_vgu | e_6_active_vcu | e_6_active_vlu | e_6_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2515 = v_6 & _T_2514; // @[sequencer-master.scala 451:34]
  wire  _T_2518 = e_7_active_vgu | e_7_active_vcu | e_7_active_vlu | e_7_active_vsu; // @[sequencer-master.scala 452:57]
  wire  _T_2519 = v_7 & _T_2518; // @[sequencer-master.scala 451:34]
  wire [1:0] _T_2520 = _T_2491 + _T_2495; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2521 = _T_2499 + _T_2503; // @[Bitwise.scala 48:55]
  wire [2:0] _T_2522 = _T_2520 + _T_2521; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2523 = _T_2507 + _T_2511; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2524 = _T_2515 + _T_2519; // @[Bitwise.scala 48:55]
  wire [2:0] _T_2525 = _T_2523 + _T_2524; // @[Bitwise.scala 48:55]
  wire [3:0] _T_2526 = _T_2522 + _T_2525; // @[Bitwise.scala 48:55]
  wire  _T_2529 = e_0_active_viu | e_0_active_vimu | e_0_active_vidu | e_0_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2533 = _T_2529 | e_0_active_vfdu | e_0_active_vfcu | e_0_active_vfvu | e_0_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2534 = v_0 & _T_2533; // @[sequencer-master.scala 455:34]
  wire  _T_2537 = e_1_active_viu | e_1_active_vimu | e_1_active_vidu | e_1_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2541 = _T_2537 | e_1_active_vfdu | e_1_active_vfcu | e_1_active_vfvu | e_1_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2542 = v_1 & _T_2541; // @[sequencer-master.scala 455:34]
  wire  _T_2545 = e_2_active_viu | e_2_active_vimu | e_2_active_vidu | e_2_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2549 = _T_2545 | e_2_active_vfdu | e_2_active_vfcu | e_2_active_vfvu | e_2_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2550 = v_2 & _T_2549; // @[sequencer-master.scala 455:34]
  wire  _T_2553 = e_3_active_viu | e_3_active_vimu | e_3_active_vidu | e_3_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2557 = _T_2553 | e_3_active_vfdu | e_3_active_vfcu | e_3_active_vfvu | e_3_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2558 = v_3 & _T_2557; // @[sequencer-master.scala 455:34]
  wire  _T_2561 = e_4_active_viu | e_4_active_vimu | e_4_active_vidu | e_4_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2565 = _T_2561 | e_4_active_vfdu | e_4_active_vfcu | e_4_active_vfvu | e_4_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2566 = v_4 & _T_2565; // @[sequencer-master.scala 455:34]
  wire  _T_2569 = e_5_active_viu | e_5_active_vimu | e_5_active_vidu | e_5_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2573 = _T_2569 | e_5_active_vfdu | e_5_active_vfcu | e_5_active_vfvu | e_5_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2574 = v_5 & _T_2573; // @[sequencer-master.scala 455:34]
  wire  _T_2577 = e_6_active_viu | e_6_active_vimu | e_6_active_vidu | e_6_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2581 = _T_2577 | e_6_active_vfdu | e_6_active_vfcu | e_6_active_vfvu | e_6_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2582 = v_6 & _T_2581; // @[sequencer-master.scala 455:34]
  wire  _T_2585 = e_7_active_viu | e_7_active_vimu | e_7_active_vidu | e_7_active_vfmu; // @[sequencer-master.scala 456:59]
  wire  _T_2589 = _T_2585 | e_7_active_vfdu | e_7_active_vfcu | e_7_active_vfvu | e_7_active_vqu; // @[sequencer-master.scala 457:76]
  wire  _T_2590 = v_7 & _T_2589; // @[sequencer-master.scala 455:34]
  wire [1:0] _T_2591 = _T_2534 + _T_2542; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2592 = _T_2550 + _T_2558; // @[Bitwise.scala 48:55]
  wire [2:0] _T_2593 = _T_2591 + _T_2592; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2594 = _T_2566 + _T_2574; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2595 = _T_2582 + _T_2590; // @[Bitwise.scala 48:55]
  wire [2:0] _T_2596 = _T_2594 + _T_2595; // @[Bitwise.scala 48:55]
  wire [3:0] _T_2597 = _T_2593 + _T_2596; // @[Bitwise.scala 48:55]
  wire  _T_2598 = e_0_active_vpu | e_0_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2599 = v_0 & _T_2598; // @[sequencer-master.scala 461:34]
  wire  _T_2600 = e_1_active_vpu | e_1_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2601 = v_1 & _T_2600; // @[sequencer-master.scala 461:34]
  wire  _T_2602 = e_2_active_vpu | e_2_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2603 = v_2 & _T_2602; // @[sequencer-master.scala 461:34]
  wire  _T_2604 = e_3_active_vpu | e_3_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2605 = v_3 & _T_2604; // @[sequencer-master.scala 461:34]
  wire  _T_2606 = e_4_active_vpu | e_4_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2607 = v_4 & _T_2606; // @[sequencer-master.scala 461:34]
  wire  _T_2608 = e_5_active_vpu | e_5_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2609 = v_5 & _T_2608; // @[sequencer-master.scala 461:34]
  wire  _T_2610 = e_6_active_vpu | e_6_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2611 = v_6 & _T_2610; // @[sequencer-master.scala 461:34]
  wire  _T_2612 = e_7_active_vpu | e_7_active_vipu; // @[sequencer-master.scala 462:25]
  wire  _T_2613 = v_7 & _T_2612; // @[sequencer-master.scala 461:34]
  wire [1:0] _T_2614 = _T_2599 + _T_2601; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2615 = _T_2603 + _T_2605; // @[Bitwise.scala 48:55]
  wire [2:0] _T_2616 = _T_2614 + _T_2615; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2617 = _T_2607 + _T_2609; // @[Bitwise.scala 48:55]
  wire [1:0] _T_2618 = _T_2611 + _T_2613; // @[Bitwise.scala 48:55]
  wire [2:0] _T_2619 = _T_2617 + _T_2618; // @[Bitwise.scala 48:55]
  wire [3:0] _T_2620 = _T_2616 + _T_2619; // @[Bitwise.scala 48:55]
  wire  new_DoPrim0 = _T_2433 | _T_2435;
  wire  new_DoPrim594 = _T_1752 & _GEN_30116;
  wire  new_DoPrim595 = _T_1752 & _GEN_30117;
  wire  new_DoPrim596 = _T_1752 & _GEN_30118;
  wire  new_DoPrim597 = _T_1752 & _GEN_30119;
  wire  new_DoPrim598 = _T_1752 & _GEN_30120;
  wire  new_DoPrim599 = _T_1752 & _GEN_30121;
  wire  new_DoPrim600 = _T_1752 & _GEN_30122;
  wire  new_DoPrim601 = _T_1752 & _GEN_30123;
  wire  new_DoPrim1056402 = _T_2479 | _T_2473;
  wire  new_DoPrim1056403 = _T_2486 | v_7;
  wire [2:0] new_DoPrim1056405 = _T_2526[2:0];
  wire [2:0] new_DoPrim1056406 = _T_2597[2:0];
  wire [2:0] new_DoPrim1056407 = _T_2620[2:0];
  wire [3:0] new_DoPrim1056411 = {_T_2411,_T_2413};
  wire  _GEN_38872 = _T_1752 & io_op_bits_active_vidiv; // @[sequencer-master.scala 298:15]
  wire  _GEN_38878 = _T_1752 & io_op_bits_active_vfdiv; // @[sequencer-master.scala 298:15]
  assign io_op_ready = new_DoPrim0; // @[sequencer-master.scala 399:66]
  assign io_master_state_valid_0 = v_0; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_1 = v_1; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_2 = v_2; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_3 = v_3; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_4 = v_4; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_5 = v_5; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_6 = v_6; // @[sequencer-master.scala 115:25]
  assign io_master_state_valid_7 = v_7; // @[sequencer-master.scala 115:25]
  assign io_master_state_e_0_fn_union = e_0_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_sreg_ss1 = e_0_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_sreg_ss2 = e_0_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_sreg_ss3 = e_0_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vp_id = e_0_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vp_valid = e_0_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vp_scalar = e_0_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vp_pred = e_0_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs1_id = e_0_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs1_valid = e_0_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs1_scalar = e_0_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs1_pred = e_0_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs1_prec = e_0_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs2_id = e_0_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs2_valid = e_0_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs2_scalar = e_0_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs2_pred = e_0_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs2_prec = e_0_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs3_id = e_0_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs3_valid = e_0_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs3_scalar = e_0_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs3_pred = e_0_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vs3_prec = e_0_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vd_id = e_0_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vd_valid = e_0_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vd_scalar = e_0_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vd_pred = e_0_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_base_vd_prec = e_0_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_viu = e_0_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vipu = e_0_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vimu = e_0_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vidu = e_0_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vfmu = e_0_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vfdu = e_0_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vfcu = e_0_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vfvu = e_0_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vpu = e_0_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vgu = e_0_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vcu = e_0_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vlu = e_0_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vsu = e_0_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_active_vqu = e_0_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_0 = e_0_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_1 = e_0_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_2 = e_0_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_3 = e_0_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_4 = e_0_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_5 = e_0_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_6 = e_0_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_raw_7 = e_0_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_0 = e_0_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_1 = e_0_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_2 = e_0_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_3 = e_0_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_4 = e_0_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_5 = e_0_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_6 = e_0_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_war_7 = e_0_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_0 = e_0_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_1 = e_0_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_2 = e_0_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_3 = e_0_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_4 = e_0_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_5 = e_0_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_6 = e_0_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_waw_7 = e_0_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_last = e_0_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_rports = e_0_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_wport_sram = e_0_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_0_wport_pred = e_0_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_fn_union = e_1_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_sreg_ss1 = e_1_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_sreg_ss2 = e_1_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_sreg_ss3 = e_1_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vp_id = e_1_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vp_valid = e_1_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vp_scalar = e_1_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vp_pred = e_1_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs1_id = e_1_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs1_valid = e_1_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs1_scalar = e_1_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs1_pred = e_1_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs1_prec = e_1_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs2_id = e_1_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs2_valid = e_1_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs2_scalar = e_1_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs2_pred = e_1_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs2_prec = e_1_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs3_id = e_1_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs3_valid = e_1_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs3_scalar = e_1_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs3_pred = e_1_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vs3_prec = e_1_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vd_id = e_1_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vd_valid = e_1_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vd_scalar = e_1_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vd_pred = e_1_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_base_vd_prec = e_1_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_viu = e_1_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vipu = e_1_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vimu = e_1_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vidu = e_1_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vfmu = e_1_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vfdu = e_1_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vfcu = e_1_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vfvu = e_1_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vpu = e_1_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vgu = e_1_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vcu = e_1_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vlu = e_1_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vsu = e_1_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_active_vqu = e_1_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_0 = e_1_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_1 = e_1_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_2 = e_1_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_3 = e_1_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_4 = e_1_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_5 = e_1_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_6 = e_1_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_raw_7 = e_1_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_0 = e_1_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_1 = e_1_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_2 = e_1_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_3 = e_1_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_4 = e_1_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_5 = e_1_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_6 = e_1_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_war_7 = e_1_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_0 = e_1_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_1 = e_1_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_2 = e_1_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_3 = e_1_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_4 = e_1_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_5 = e_1_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_6 = e_1_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_waw_7 = e_1_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_last = e_1_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_rports = e_1_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_wport_sram = e_1_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_1_wport_pred = e_1_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_fn_union = e_2_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_sreg_ss1 = e_2_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_sreg_ss2 = e_2_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_sreg_ss3 = e_2_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vp_id = e_2_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vp_valid = e_2_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vp_scalar = e_2_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vp_pred = e_2_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs1_id = e_2_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs1_valid = e_2_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs1_scalar = e_2_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs1_pred = e_2_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs1_prec = e_2_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs2_id = e_2_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs2_valid = e_2_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs2_scalar = e_2_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs2_pred = e_2_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs2_prec = e_2_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs3_id = e_2_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs3_valid = e_2_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs3_scalar = e_2_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs3_pred = e_2_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vs3_prec = e_2_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vd_id = e_2_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vd_valid = e_2_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vd_scalar = e_2_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vd_pred = e_2_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_base_vd_prec = e_2_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_viu = e_2_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vipu = e_2_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vimu = e_2_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vidu = e_2_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vfmu = e_2_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vfdu = e_2_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vfcu = e_2_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vfvu = e_2_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vpu = e_2_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vgu = e_2_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vcu = e_2_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vlu = e_2_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vsu = e_2_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_active_vqu = e_2_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_0 = e_2_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_1 = e_2_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_2 = e_2_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_3 = e_2_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_4 = e_2_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_5 = e_2_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_6 = e_2_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_raw_7 = e_2_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_0 = e_2_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_1 = e_2_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_2 = e_2_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_3 = e_2_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_4 = e_2_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_5 = e_2_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_6 = e_2_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_war_7 = e_2_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_0 = e_2_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_1 = e_2_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_2 = e_2_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_3 = e_2_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_4 = e_2_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_5 = e_2_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_6 = e_2_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_waw_7 = e_2_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_last = e_2_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_rports = e_2_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_wport_sram = e_2_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_2_wport_pred = e_2_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_fn_union = e_3_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_sreg_ss1 = e_3_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_sreg_ss2 = e_3_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_sreg_ss3 = e_3_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vp_id = e_3_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vp_valid = e_3_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vp_scalar = e_3_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vp_pred = e_3_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs1_id = e_3_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs1_valid = e_3_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs1_scalar = e_3_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs1_pred = e_3_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs1_prec = e_3_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs2_id = e_3_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs2_valid = e_3_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs2_scalar = e_3_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs2_pred = e_3_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs2_prec = e_3_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs3_id = e_3_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs3_valid = e_3_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs3_scalar = e_3_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs3_pred = e_3_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vs3_prec = e_3_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vd_id = e_3_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vd_valid = e_3_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vd_scalar = e_3_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vd_pred = e_3_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_base_vd_prec = e_3_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_viu = e_3_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vipu = e_3_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vimu = e_3_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vidu = e_3_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vfmu = e_3_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vfdu = e_3_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vfcu = e_3_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vfvu = e_3_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vpu = e_3_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vgu = e_3_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vcu = e_3_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vlu = e_3_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vsu = e_3_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_active_vqu = e_3_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_0 = e_3_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_1 = e_3_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_2 = e_3_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_3 = e_3_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_4 = e_3_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_5 = e_3_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_6 = e_3_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_raw_7 = e_3_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_0 = e_3_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_1 = e_3_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_2 = e_3_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_3 = e_3_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_4 = e_3_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_5 = e_3_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_6 = e_3_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_war_7 = e_3_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_0 = e_3_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_1 = e_3_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_2 = e_3_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_3 = e_3_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_4 = e_3_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_5 = e_3_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_6 = e_3_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_waw_7 = e_3_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_last = e_3_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_rports = e_3_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_wport_sram = e_3_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_3_wport_pred = e_3_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_fn_union = e_4_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_sreg_ss1 = e_4_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_sreg_ss2 = e_4_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_sreg_ss3 = e_4_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vp_id = e_4_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vp_valid = e_4_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vp_scalar = e_4_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vp_pred = e_4_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs1_id = e_4_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs1_valid = e_4_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs1_scalar = e_4_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs1_pred = e_4_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs1_prec = e_4_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs2_id = e_4_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs2_valid = e_4_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs2_scalar = e_4_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs2_pred = e_4_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs2_prec = e_4_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs3_id = e_4_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs3_valid = e_4_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs3_scalar = e_4_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs3_pred = e_4_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vs3_prec = e_4_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vd_id = e_4_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vd_valid = e_4_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vd_scalar = e_4_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vd_pred = e_4_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_base_vd_prec = e_4_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_viu = e_4_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vipu = e_4_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vimu = e_4_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vidu = e_4_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vfmu = e_4_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vfdu = e_4_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vfcu = e_4_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vfvu = e_4_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vpu = e_4_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vgu = e_4_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vcu = e_4_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vlu = e_4_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vsu = e_4_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_active_vqu = e_4_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_0 = e_4_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_1 = e_4_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_2 = e_4_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_3 = e_4_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_4 = e_4_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_5 = e_4_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_6 = e_4_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_raw_7 = e_4_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_0 = e_4_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_1 = e_4_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_2 = e_4_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_3 = e_4_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_4 = e_4_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_5 = e_4_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_6 = e_4_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_war_7 = e_4_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_0 = e_4_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_1 = e_4_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_2 = e_4_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_3 = e_4_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_4 = e_4_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_5 = e_4_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_6 = e_4_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_waw_7 = e_4_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_last = e_4_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_rports = e_4_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_wport_sram = e_4_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_4_wport_pred = e_4_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_fn_union = e_5_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_sreg_ss1 = e_5_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_sreg_ss2 = e_5_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_sreg_ss3 = e_5_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vp_id = e_5_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vp_valid = e_5_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vp_scalar = e_5_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vp_pred = e_5_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs1_id = e_5_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs1_valid = e_5_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs1_scalar = e_5_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs1_pred = e_5_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs1_prec = e_5_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs2_id = e_5_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs2_valid = e_5_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs2_scalar = e_5_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs2_pred = e_5_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs2_prec = e_5_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs3_id = e_5_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs3_valid = e_5_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs3_scalar = e_5_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs3_pred = e_5_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vs3_prec = e_5_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vd_id = e_5_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vd_valid = e_5_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vd_scalar = e_5_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vd_pred = e_5_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_base_vd_prec = e_5_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_viu = e_5_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vipu = e_5_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vimu = e_5_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vidu = e_5_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vfmu = e_5_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vfdu = e_5_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vfcu = e_5_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vfvu = e_5_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vpu = e_5_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vgu = e_5_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vcu = e_5_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vlu = e_5_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vsu = e_5_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_active_vqu = e_5_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_0 = e_5_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_1 = e_5_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_2 = e_5_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_3 = e_5_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_4 = e_5_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_5 = e_5_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_6 = e_5_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_raw_7 = e_5_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_0 = e_5_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_1 = e_5_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_2 = e_5_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_3 = e_5_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_4 = e_5_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_5 = e_5_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_6 = e_5_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_war_7 = e_5_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_0 = e_5_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_1 = e_5_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_2 = e_5_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_3 = e_5_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_4 = e_5_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_5 = e_5_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_6 = e_5_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_waw_7 = e_5_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_last = e_5_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_rports = e_5_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_wport_sram = e_5_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_5_wport_pred = e_5_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_fn_union = e_6_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_sreg_ss1 = e_6_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_sreg_ss2 = e_6_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_sreg_ss3 = e_6_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vp_id = e_6_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vp_valid = e_6_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vp_scalar = e_6_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vp_pred = e_6_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs1_id = e_6_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs1_valid = e_6_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs1_scalar = e_6_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs1_pred = e_6_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs1_prec = e_6_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs2_id = e_6_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs2_valid = e_6_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs2_scalar = e_6_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs2_pred = e_6_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs2_prec = e_6_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs3_id = e_6_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs3_valid = e_6_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs3_scalar = e_6_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs3_pred = e_6_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vs3_prec = e_6_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vd_id = e_6_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vd_valid = e_6_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vd_scalar = e_6_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vd_pred = e_6_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_base_vd_prec = e_6_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_viu = e_6_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vipu = e_6_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vimu = e_6_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vidu = e_6_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vfmu = e_6_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vfdu = e_6_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vfcu = e_6_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vfvu = e_6_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vpu = e_6_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vgu = e_6_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vcu = e_6_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vlu = e_6_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vsu = e_6_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_active_vqu = e_6_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_0 = e_6_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_1 = e_6_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_2 = e_6_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_3 = e_6_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_4 = e_6_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_5 = e_6_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_6 = e_6_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_raw_7 = e_6_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_0 = e_6_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_1 = e_6_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_2 = e_6_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_3 = e_6_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_4 = e_6_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_5 = e_6_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_6 = e_6_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_war_7 = e_6_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_0 = e_6_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_1 = e_6_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_2 = e_6_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_3 = e_6_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_4 = e_6_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_5 = e_6_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_6 = e_6_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_waw_7 = e_6_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_last = e_6_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_rports = e_6_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_wport_sram = e_6_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_6_wport_pred = e_6_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_fn_union = e_7_fn_union; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_sreg_ss1 = e_7_sreg_ss1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_sreg_ss2 = e_7_sreg_ss2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_sreg_ss3 = e_7_sreg_ss3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vp_id = e_7_base_vp_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vp_valid = e_7_base_vp_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vp_scalar = e_7_base_vp_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vp_pred = e_7_base_vp_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs1_id = e_7_base_vs1_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs1_valid = e_7_base_vs1_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs1_scalar = e_7_base_vs1_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs1_pred = e_7_base_vs1_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs1_prec = e_7_base_vs1_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs2_id = e_7_base_vs2_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs2_valid = e_7_base_vs2_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs2_scalar = e_7_base_vs2_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs2_pred = e_7_base_vs2_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs2_prec = e_7_base_vs2_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs3_id = e_7_base_vs3_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs3_valid = e_7_base_vs3_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs3_scalar = e_7_base_vs3_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs3_pred = e_7_base_vs3_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vs3_prec = e_7_base_vs3_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vd_id = e_7_base_vd_id; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vd_valid = e_7_base_vd_valid; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vd_scalar = e_7_base_vd_scalar; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vd_pred = e_7_base_vd_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_base_vd_prec = e_7_base_vd_prec; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_rate = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_viu = e_7_active_viu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vipu = e_7_active_vipu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vimu = e_7_active_vimu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vidu = e_7_active_vidu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vfmu = e_7_active_vfmu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vfdu = e_7_active_vfdu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vfcu = e_7_active_vfcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vfvu = e_7_active_vfvu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vrpu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vrfu = 1'h0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vpu = e_7_active_vpu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vgu = e_7_active_vgu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vcu = e_7_active_vcu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vlu = e_7_active_vlu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vsu = e_7_active_vsu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_active_vqu = e_7_active_vqu; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_0 = e_7_raw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_1 = e_7_raw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_2 = e_7_raw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_3 = e_7_raw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_4 = e_7_raw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_5 = e_7_raw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_6 = e_7_raw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_raw_7 = e_7_raw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_0 = e_7_war_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_1 = e_7_war_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_2 = e_7_war_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_3 = e_7_war_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_4 = e_7_war_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_5 = e_7_war_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_6 = e_7_war_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_war_7 = e_7_war_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_0 = e_7_waw_0; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_1 = e_7_waw_1; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_2 = e_7_waw_2; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_3 = e_7_waw_3; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_4 = e_7_waw_4; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_5 = e_7_waw_5; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_6 = e_7_waw_6; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_waw_7 = e_7_waw_7; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_last = e_7_last; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_rports = e_7_rports; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_wport_sram = e_7_wport_sram; // @[sequencer-master.scala 116:21]
  assign io_master_state_e_7_wport_pred = e_7_wport_pred; // @[sequencer-master.scala 116:21]
  assign io_master_state_head = head; // @[sequencer-master.scala 117:24]
  assign io_master_update_valid_0 = new_DoPrim594; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_1 = new_DoPrim595; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_2 = new_DoPrim596; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_3 = new_DoPrim597; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_4 = new_DoPrim598; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_5 = new_DoPrim599; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_6 = new_DoPrim600; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_valid_7 = new_DoPrim601; // @[sequencer-master.scala 639:27 sequencer-master.scala 410:35]
  assign io_master_update_reg_0_vp_id = _T_1752 ? _GEN_30372 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_0_vs1_id = _T_1752 ? _GEN_30452 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_0_vs2_id = _T_1752 ? _GEN_14532 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_0_vs3_id = _T_1752 ? _GEN_10224 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_0_vd_id = _T_1752 ? _GEN_28410 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_1_vp_id = _T_1752 ? _GEN_30373 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_1_vs1_id = _T_1752 ? _GEN_30453 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_1_vs2_id = _T_1752 ? _GEN_14533 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_1_vs3_id = _T_1752 ? _GEN_10225 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_1_vd_id = _T_1752 ? _GEN_28411 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_2_vp_id = _T_1752 ? _GEN_30374 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_2_vs1_id = _T_1752 ? _GEN_30454 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_2_vs2_id = _T_1752 ? _GEN_14534 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_2_vs3_id = _T_1752 ? _GEN_10226 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_2_vd_id = _T_1752 ? _GEN_28412 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_3_vp_id = _T_1752 ? _GEN_30375 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_3_vs1_id = _T_1752 ? _GEN_30455 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_3_vs2_id = _T_1752 ? _GEN_14535 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_3_vs3_id = _T_1752 ? _GEN_10227 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_3_vd_id = _T_1752 ? _GEN_28413 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_4_vp_id = _T_1752 ? _GEN_30376 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_4_vs1_id = _T_1752 ? _GEN_30456 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_4_vs2_id = _T_1752 ? _GEN_14536 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_4_vs3_id = _T_1752 ? _GEN_10228 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_4_vd_id = _T_1752 ? _GEN_28414 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_5_vp_id = _T_1752 ? _GEN_30377 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_5_vs1_id = _T_1752 ? _GEN_30457 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_5_vs2_id = _T_1752 ? _GEN_14537 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_5_vs3_id = _T_1752 ? _GEN_10229 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_5_vd_id = _T_1752 ? _GEN_28415 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_6_vp_id = _T_1752 ? _GEN_30378 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_6_vs1_id = _T_1752 ? _GEN_30458 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_6_vs2_id = _T_1752 ? _GEN_14538 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_6_vs3_id = _T_1752 ? _GEN_10230 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_6_vd_id = _T_1752 ? _GEN_28416 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_7_vp_id = _T_1752 ? _GEN_30379 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_7_vs1_id = _T_1752 ? _GEN_30459 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_7_vs2_id = _T_1752 ? _GEN_14539 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_7_vs3_id = _T_1752 ? _GEN_10231 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_master_update_reg_7_vd_id = _T_1752 ? _GEN_28417 : 8'h0; // @[sequencer-master.scala 639:27 sequencer-master.scala 411:33]
  assign io_pending_mem = new_DoPrim1056402; // @[sequencer-master.scala 447:39]
  assign io_pending_all = new_DoPrim1056403; // @[sequencer-master.scala 448:36]
  assign io_vf_last = _T_2465; // @[sequencer-master.scala 444:18]
  assign io_counters_memoryUOps = new_DoPrim1056405; // @[sequencer-master.scala 450:30]
  assign io_counters_arithUOps = new_DoPrim1056406; // @[sequencer-master.scala 454:29]
  assign io_counters_predUOps = new_DoPrim1056407; // @[sequencer-master.scala 460:28]
  assign io_debug_head = head; // @[sequencer-master.scala 478:21]
  assign io_debug_tail = tail; // @[sequencer-master.scala 479:21]
  assign io_debug_maybe_full = maybe_full; // @[sequencer-master.scala 477:27]
  assign io_debug_empty = new_DoPrim1056411; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_0 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_0 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 372:35]
        v_0 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_0 <= _GEN_30462;
      end
    end else begin
      v_0 <= _GEN_30462;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_1 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_1 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 372:35]
        v_1 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_1 <= _GEN_30463;
      end
    end else begin
      v_1 <= _GEN_30463;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_2 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_2 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 372:35]
        v_2 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_2 <= _GEN_30464;
      end
    end else begin
      v_2 <= _GEN_30464;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_3 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_3 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 372:35]
        v_3 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_3 <= _GEN_30465;
      end
    end else begin
      v_3 <= _GEN_30465;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_4 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_4 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 372:35]
        v_4 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_4 <= _GEN_30466;
      end
    end else begin
      v_4 <= _GEN_30466;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_5 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_5 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 372:35]
        v_5 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_5 <= _GEN_30467;
      end
    end else begin
      v_5 <= _GEN_30467;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_6 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_6 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 372:35]
        v_6 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_6 <= _GEN_30468;
      end
    end else begin
      v_6 <= _GEN_30468;
    end
    if (reset) begin // @[sequencer-master.scala 107:14]
      v_7 <= 1'h0; // @[sequencer-master.scala 107:14]
    end else if (reset) begin // @[sequencer-master.scala 468:20]
      v_7 <= 1'h0; // @[sequencer-master.scala 372:35]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 372:35]
        v_7 <= 1'h0; // @[sequencer-master.scala 372:35]
      end else begin
        v_7 <= _GEN_30469;
      end
    end else begin
      v_7 <= _GEN_30469;
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_0_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_0_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_0_fn_union <= _GEN_28700;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_0_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_0_fn_union <= _GEN_27066;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_fn_union <= _GEN_25328;
      end else begin
        e_0_fn_union <= _GEN_23798;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_0_sreg_ss1 <= _GEN_24512;
          end else begin
            e_0_sreg_ss1 <= _GEN_23878;
          end
        end else begin
          e_0_sreg_ss1 <= _GEN_23878;
        end
      end else begin
        e_0_sreg_ss1 <= _GEN_23878;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_0_sreg_ss2 <= _GEN_13524;
          end else begin
            e_0_sreg_ss2 <= _GEN_12650;
          end
        end else begin
          e_0_sreg_ss2 <= _GEN_12650;
        end
      end else begin
        e_0_sreg_ss2 <= _GEN_12650;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_0_sreg_ss3 <= _GEN_9168;
          end else begin
            e_0_sreg_ss3 <= _GEN_3746;
          end
        end else begin
          e_0_sreg_ss3 <= _GEN_3746;
        end
      end else begin
        e_0_sreg_ss3 <= _GEN_3746;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_0_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_0_base_vp_id <= _GEN_28748;
          end
        end else begin
          e_0_base_vp_id <= _GEN_28748;
        end
      end else begin
        e_0_base_vp_id <= _GEN_28306;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_0_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_0_base_vp_valid <= _GEN_29268;
          end
        end else begin
          e_0_base_vp_valid <= _GEN_29268;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_0_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_0_base_vp_valid <= _GEN_26802;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_base_vp_valid <= _GEN_25384;
      end else begin
        e_0_base_vp_valid <= _GEN_23534;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_0_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_0_base_vp_scalar <= _GEN_28764;
          end
        end else begin
          e_0_base_vp_scalar <= _GEN_28764;
        end
      end else begin
        e_0_base_vp_scalar <= _GEN_28314;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_0_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_0_base_vp_pred <= _GEN_28772;
          end
        end else begin
          e_0_base_vp_pred <= _GEN_28772;
        end
      end else begin
        e_0_base_vp_pred <= _GEN_28322;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_0_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_0_base_vs1_id <= _GEN_26176;
          end
        end else begin
          e_0_base_vs1_id <= _GEN_26176;
        end
      end else begin
        e_0_base_vs1_id <= _GEN_26176;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_0_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_0_base_vs1_valid <= _GEN_29276;
          end
        end else begin
          e_0_base_vs1_valid <= _GEN_29276;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_0_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_0_base_vs1_valid <= _GEN_26810;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_base_vs1_valid <= _GEN_25600;
      end else begin
        e_0_base_vs1_valid <= _GEN_23542;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_0_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_0_base_vs1_scalar <= _GEN_26184;
          end
        end else begin
          e_0_base_vs1_scalar <= _GEN_26184;
        end
      end else begin
        e_0_base_vs1_scalar <= _GEN_26184;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_0_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_0_base_vs1_pred <= _GEN_26192;
          end
        end else begin
          e_0_base_vs1_pred <= _GEN_26192;
        end
      end else begin
        e_0_base_vs1_pred <= _GEN_26192;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_0_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_0_base_vs1_prec <= _GEN_26200;
          end
        end else begin
          e_0_base_vs1_prec <= _GEN_26200;
        end
      end else begin
        e_0_base_vs1_prec <= _GEN_26200;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs2_id <= _GEN_12610;
          end
        end else begin
          e_0_base_vs2_id <= _GEN_12610;
        end
      end else begin
        e_0_base_vs2_id <= _GEN_12610;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_0_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_0_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_0_base_vs2_valid <= _GEN_28452;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_0_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_0_base_vs2_valid <= _GEN_26818;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_base_vs2_valid <= _GEN_25080;
      end else begin
        e_0_base_vs2_valid <= _GEN_23550;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs2_scalar <= _GEN_12618;
          end
        end else begin
          e_0_base_vs2_scalar <= _GEN_12618;
        end
      end else begin
        e_0_base_vs2_scalar <= _GEN_12618;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs2_pred <= _GEN_12626;
          end
        end else begin
          e_0_base_vs2_pred <= _GEN_12626;
        end
      end else begin
        e_0_base_vs2_pred <= _GEN_12626;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs2_prec <= _GEN_12634;
          end
        end else begin
          e_0_base_vs2_prec <= _GEN_12634;
        end
      end else begin
        e_0_base_vs2_prec <= _GEN_12634;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs3_id <= _GEN_3706;
          end
        end else begin
          e_0_base_vs3_id <= _GEN_3706;
        end
      end else begin
        e_0_base_vs3_id <= _GEN_3706;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_0_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_0_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_0_base_vs3_valid <= _GEN_28460;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_0_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_0_base_vs3_valid <= _GEN_26826;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_base_vs3_valid <= _GEN_25088;
      end else begin
        e_0_base_vs3_valid <= _GEN_23558;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs3_scalar <= _GEN_3714;
          end
        end else begin
          e_0_base_vs3_scalar <= _GEN_3714;
        end
      end else begin
        e_0_base_vs3_scalar <= _GEN_3714;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs3_pred <= _GEN_3722;
          end
        end else begin
          e_0_base_vs3_pred <= _GEN_3722;
        end
      end else begin
        e_0_base_vs3_pred <= _GEN_3722;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h0 == tail) begin // @[sequencer-master.scala 329:29]
            e_0_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_0_base_vs3_prec <= _GEN_3730;
          end
        end else begin
          e_0_base_vs3_prec <= _GEN_3730;
        end
      end else begin
        e_0_base_vs3_prec <= _GEN_3730;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_0_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_0_base_vd_id <= _GEN_23926;
          end
        end else begin
          e_0_base_vd_id <= _GEN_23926;
        end
      end else begin
        e_0_base_vd_id <= _GEN_23926;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_0_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_0_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_0_base_vd_valid <= _GEN_28468;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_0_base_vd_valid <= _GEN_27650;
        end else begin
          e_0_base_vd_valid <= _GEN_27402;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_base_vd_valid <= _GEN_25096;
      end else begin
        e_0_base_vd_valid <= _GEN_23566;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_0_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_0_base_vd_scalar <= _GEN_23934;
          end
        end else begin
          e_0_base_vd_scalar <= _GEN_23934;
        end
      end else begin
        e_0_base_vd_scalar <= _GEN_23934;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_0_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_0_base_vd_pred <= _GEN_23942;
          end
        end else begin
          e_0_base_vd_pred <= _GEN_23942;
        end
      end else begin
        e_0_base_vd_pred <= _GEN_23942;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h0 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_0_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_0_base_vd_prec <= _GEN_23950;
          end
        end else begin
          e_0_base_vd_prec <= _GEN_23950;
        end
      end else begin
        e_0_base_vd_prec <= _GEN_23950;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_viu <= _GEN_30734;
      end
    end else begin
      e_0_active_viu <= _GEN_30734;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vipu <= _GEN_30944;
      end
    end else begin
      e_0_active_vipu <= _GEN_30944;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vimu <= _GEN_31000;
      end
    end else begin
      e_0_active_vimu <= _GEN_31000;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vidu <= _GEN_31016;
      end
    end else begin
      e_0_active_vidu <= _GEN_31016;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vfmu <= _GEN_31024;
      end
    end else begin
      e_0_active_vfmu <= _GEN_31024;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vfdu <= _GEN_31032;
      end
    end else begin
      e_0_active_vfdu <= _GEN_31032;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vfcu <= _GEN_31040;
      end
    end else begin
      e_0_active_vfcu <= _GEN_31040;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vfvu <= _GEN_31048;
      end
    end else begin
      e_0_active_vfvu <= _GEN_31048;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vpu <= _GEN_31088;
      end
    end else begin
      e_0_active_vpu <= _GEN_31088;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vgu <= _GEN_31056;
      end
    end else begin
      e_0_active_vgu <= _GEN_31056;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vcu <= _GEN_31064;
      end
    end else begin
      e_0_active_vcu <= _GEN_31064;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vlu <= _GEN_31080;
      end
    end else begin
      e_0_active_vlu <= _GEN_31080;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vsu <= _GEN_31072;
      end
    end else begin
      e_0_active_vsu <= _GEN_31072;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_0_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h0 == head) begin // @[sequencer-master.scala 373:43]
        e_0_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_0_active_vqu <= _GEN_31008;
      end
    end else begin
      e_0_active_vqu <= _GEN_31008;
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_0 <= _GEN_30526;
        end
      end else begin
        e_0_raw_0 <= _GEN_30526;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_1 <= _GEN_30550;
        end
      end else begin
        e_0_raw_1 <= _GEN_30550;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_2 <= _GEN_30574;
        end
      end else begin
        e_0_raw_2 <= _GEN_30574;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_3 <= _GEN_30598;
        end
      end else begin
        e_0_raw_3 <= _GEN_30598;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_4 <= _GEN_30622;
        end
      end else begin
        e_0_raw_4 <= _GEN_30622;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_5 <= _GEN_30646;
        end
      end else begin
        e_0_raw_5 <= _GEN_30646;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_6 <= _GEN_30670;
        end
      end else begin
        e_0_raw_6 <= _GEN_30670;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_0_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_0_raw_7 <= _GEN_30694;
        end
      end else begin
        e_0_raw_7 <= _GEN_30694;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_0 <= _GEN_30534;
        end
      end else begin
        e_0_war_0 <= _GEN_30534;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_1 <= _GEN_30558;
        end
      end else begin
        e_0_war_1 <= _GEN_30558;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_2 <= _GEN_30582;
        end
      end else begin
        e_0_war_2 <= _GEN_30582;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_3 <= _GEN_30606;
        end
      end else begin
        e_0_war_3 <= _GEN_30606;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_4 <= _GEN_30630;
        end
      end else begin
        e_0_war_4 <= _GEN_30630;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_5 <= _GEN_30654;
        end
      end else begin
        e_0_war_5 <= _GEN_30654;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_6 <= _GEN_30678;
        end
      end else begin
        e_0_war_6 <= _GEN_30678;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_0_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_0_war_7 <= _GEN_30702;
        end
      end else begin
        e_0_war_7 <= _GEN_30702;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_0 <= _GEN_30542;
        end
      end else begin
        e_0_waw_0 <= _GEN_30542;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_1 <= _GEN_30566;
        end
      end else begin
        e_0_waw_1 <= _GEN_30566;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_2 <= _GEN_30590;
        end
      end else begin
        e_0_waw_2 <= _GEN_30590;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_3 <= _GEN_30614;
        end
      end else begin
        e_0_waw_3 <= _GEN_30614;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_4 <= _GEN_30638;
        end
      end else begin
        e_0_waw_4 <= _GEN_30638;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_5 <= _GEN_30662;
        end
      end else begin
        e_0_waw_5 <= _GEN_30662;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_6 <= _GEN_30686;
        end
      end else begin
        e_0_waw_6 <= _GEN_30686;
      end
    end
    if (_GEN_32181) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_0_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_0_waw_7 <= _GEN_30710;
        end
      end else begin
        e_0_waw_7 <= _GEN_30710;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_0_last <= _GEN_31100;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_0_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_0_last <= _GEN_29196;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_0_last <= _GEN_27610;
      end else begin
        e_0_last <= _GEN_26112;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_0_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_0_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_0_rports <= _GEN_28916;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_0_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_0_rports <= _GEN_27074;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_rports <= _GEN_25768;
      end else begin
        e_0_rports <= _GEN_23886;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_0_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_0_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_0_wport_sram <= _GEN_28924;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_0_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_0_wport_sram <= _GEN_27082;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_wport_sram <= _GEN_25776;
      end else begin
        e_0_wport_sram <= _GEN_23894;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_0_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h0 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_0_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_0_wport_pred <= _GEN_28932;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h0 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_0_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_0_wport_pred <= _GEN_27090;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_0_wport_pred <= _GEN_25784;
      end else begin
        e_0_wport_pred <= _GEN_23902;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_1_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_1_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_1_fn_union <= _GEN_28701;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_1_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_1_fn_union <= _GEN_27067;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_fn_union <= _GEN_25329;
      end else begin
        e_1_fn_union <= _GEN_23799;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_1_sreg_ss1 <= _GEN_24513;
          end else begin
            e_1_sreg_ss1 <= _GEN_23879;
          end
        end else begin
          e_1_sreg_ss1 <= _GEN_23879;
        end
      end else begin
        e_1_sreg_ss1 <= _GEN_23879;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_1_sreg_ss2 <= _GEN_13525;
          end else begin
            e_1_sreg_ss2 <= _GEN_12651;
          end
        end else begin
          e_1_sreg_ss2 <= _GEN_12651;
        end
      end else begin
        e_1_sreg_ss2 <= _GEN_12651;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_1_sreg_ss3 <= _GEN_9169;
          end else begin
            e_1_sreg_ss3 <= _GEN_3747;
          end
        end else begin
          e_1_sreg_ss3 <= _GEN_3747;
        end
      end else begin
        e_1_sreg_ss3 <= _GEN_3747;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_1_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_1_base_vp_id <= _GEN_28749;
          end
        end else begin
          e_1_base_vp_id <= _GEN_28749;
        end
      end else begin
        e_1_base_vp_id <= _GEN_28307;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_1_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_1_base_vp_valid <= _GEN_29269;
          end
        end else begin
          e_1_base_vp_valid <= _GEN_29269;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_1_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_1_base_vp_valid <= _GEN_26803;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_base_vp_valid <= _GEN_25385;
      end else begin
        e_1_base_vp_valid <= _GEN_23535;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_1_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_1_base_vp_scalar <= _GEN_28765;
          end
        end else begin
          e_1_base_vp_scalar <= _GEN_28765;
        end
      end else begin
        e_1_base_vp_scalar <= _GEN_28315;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_1_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_1_base_vp_pred <= _GEN_28773;
          end
        end else begin
          e_1_base_vp_pred <= _GEN_28773;
        end
      end else begin
        e_1_base_vp_pred <= _GEN_28323;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_1_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_1_base_vs1_id <= _GEN_26177;
          end
        end else begin
          e_1_base_vs1_id <= _GEN_26177;
        end
      end else begin
        e_1_base_vs1_id <= _GEN_26177;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_1_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_1_base_vs1_valid <= _GEN_29277;
          end
        end else begin
          e_1_base_vs1_valid <= _GEN_29277;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_1_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_1_base_vs1_valid <= _GEN_26811;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_base_vs1_valid <= _GEN_25601;
      end else begin
        e_1_base_vs1_valid <= _GEN_23543;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_1_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_1_base_vs1_scalar <= _GEN_26185;
          end
        end else begin
          e_1_base_vs1_scalar <= _GEN_26185;
        end
      end else begin
        e_1_base_vs1_scalar <= _GEN_26185;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_1_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_1_base_vs1_pred <= _GEN_26193;
          end
        end else begin
          e_1_base_vs1_pred <= _GEN_26193;
        end
      end else begin
        e_1_base_vs1_pred <= _GEN_26193;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_1_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_1_base_vs1_prec <= _GEN_26201;
          end
        end else begin
          e_1_base_vs1_prec <= _GEN_26201;
        end
      end else begin
        e_1_base_vs1_prec <= _GEN_26201;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs2_id <= _GEN_12611;
          end
        end else begin
          e_1_base_vs2_id <= _GEN_12611;
        end
      end else begin
        e_1_base_vs2_id <= _GEN_12611;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_1_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_1_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_1_base_vs2_valid <= _GEN_28453;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_1_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_1_base_vs2_valid <= _GEN_26819;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_base_vs2_valid <= _GEN_25081;
      end else begin
        e_1_base_vs2_valid <= _GEN_23551;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs2_scalar <= _GEN_12619;
          end
        end else begin
          e_1_base_vs2_scalar <= _GEN_12619;
        end
      end else begin
        e_1_base_vs2_scalar <= _GEN_12619;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs2_pred <= _GEN_12627;
          end
        end else begin
          e_1_base_vs2_pred <= _GEN_12627;
        end
      end else begin
        e_1_base_vs2_pred <= _GEN_12627;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs2_prec <= _GEN_12635;
          end
        end else begin
          e_1_base_vs2_prec <= _GEN_12635;
        end
      end else begin
        e_1_base_vs2_prec <= _GEN_12635;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs3_id <= _GEN_3707;
          end
        end else begin
          e_1_base_vs3_id <= _GEN_3707;
        end
      end else begin
        e_1_base_vs3_id <= _GEN_3707;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_1_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_1_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_1_base_vs3_valid <= _GEN_28461;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_1_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_1_base_vs3_valid <= _GEN_26827;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_base_vs3_valid <= _GEN_25089;
      end else begin
        e_1_base_vs3_valid <= _GEN_23559;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs3_scalar <= _GEN_3715;
          end
        end else begin
          e_1_base_vs3_scalar <= _GEN_3715;
        end
      end else begin
        e_1_base_vs3_scalar <= _GEN_3715;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs3_pred <= _GEN_3723;
          end
        end else begin
          e_1_base_vs3_pred <= _GEN_3723;
        end
      end else begin
        e_1_base_vs3_pred <= _GEN_3723;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h1 == tail) begin // @[sequencer-master.scala 329:29]
            e_1_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_1_base_vs3_prec <= _GEN_3731;
          end
        end else begin
          e_1_base_vs3_prec <= _GEN_3731;
        end
      end else begin
        e_1_base_vs3_prec <= _GEN_3731;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_1_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_1_base_vd_id <= _GEN_23927;
          end
        end else begin
          e_1_base_vd_id <= _GEN_23927;
        end
      end else begin
        e_1_base_vd_id <= _GEN_23927;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_1_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_1_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_1_base_vd_valid <= _GEN_28469;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_1_base_vd_valid <= _GEN_27651;
        end else begin
          e_1_base_vd_valid <= _GEN_27403;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_base_vd_valid <= _GEN_25097;
      end else begin
        e_1_base_vd_valid <= _GEN_23567;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_1_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_1_base_vd_scalar <= _GEN_23935;
          end
        end else begin
          e_1_base_vd_scalar <= _GEN_23935;
        end
      end else begin
        e_1_base_vd_scalar <= _GEN_23935;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_1_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_1_base_vd_pred <= _GEN_23943;
          end
        end else begin
          e_1_base_vd_pred <= _GEN_23943;
        end
      end else begin
        e_1_base_vd_pred <= _GEN_23943;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h1 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_1_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_1_base_vd_prec <= _GEN_23951;
          end
        end else begin
          e_1_base_vd_prec <= _GEN_23951;
        end
      end else begin
        e_1_base_vd_prec <= _GEN_23951;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_viu <= _GEN_30735;
      end
    end else begin
      e_1_active_viu <= _GEN_30735;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vipu <= _GEN_30945;
      end
    end else begin
      e_1_active_vipu <= _GEN_30945;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vimu <= _GEN_31001;
      end
    end else begin
      e_1_active_vimu <= _GEN_31001;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vidu <= _GEN_31017;
      end
    end else begin
      e_1_active_vidu <= _GEN_31017;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vfmu <= _GEN_31025;
      end
    end else begin
      e_1_active_vfmu <= _GEN_31025;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vfdu <= _GEN_31033;
      end
    end else begin
      e_1_active_vfdu <= _GEN_31033;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vfcu <= _GEN_31041;
      end
    end else begin
      e_1_active_vfcu <= _GEN_31041;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vfvu <= _GEN_31049;
      end
    end else begin
      e_1_active_vfvu <= _GEN_31049;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vpu <= _GEN_31089;
      end
    end else begin
      e_1_active_vpu <= _GEN_31089;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vgu <= _GEN_31057;
      end
    end else begin
      e_1_active_vgu <= _GEN_31057;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vcu <= _GEN_31065;
      end
    end else begin
      e_1_active_vcu <= _GEN_31065;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vlu <= _GEN_31081;
      end
    end else begin
      e_1_active_vlu <= _GEN_31081;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vsu <= _GEN_31073;
      end
    end else begin
      e_1_active_vsu <= _GEN_31073;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_1_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h1 == head) begin // @[sequencer-master.scala 373:43]
        e_1_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_1_active_vqu <= _GEN_31009;
      end
    end else begin
      e_1_active_vqu <= _GEN_31009;
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_0 <= _GEN_30527;
        end
      end else begin
        e_1_raw_0 <= _GEN_30527;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_1 <= _GEN_30551;
        end
      end else begin
        e_1_raw_1 <= _GEN_30551;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_2 <= _GEN_30575;
        end
      end else begin
        e_1_raw_2 <= _GEN_30575;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_3 <= _GEN_30599;
        end
      end else begin
        e_1_raw_3 <= _GEN_30599;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_4 <= _GEN_30623;
        end
      end else begin
        e_1_raw_4 <= _GEN_30623;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_5 <= _GEN_30647;
        end
      end else begin
        e_1_raw_5 <= _GEN_30647;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_6 <= _GEN_30671;
        end
      end else begin
        e_1_raw_6 <= _GEN_30671;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_1_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_1_raw_7 <= _GEN_30695;
        end
      end else begin
        e_1_raw_7 <= _GEN_30695;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_0 <= _GEN_30535;
        end
      end else begin
        e_1_war_0 <= _GEN_30535;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_1 <= _GEN_30559;
        end
      end else begin
        e_1_war_1 <= _GEN_30559;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_2 <= _GEN_30583;
        end
      end else begin
        e_1_war_2 <= _GEN_30583;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_3 <= _GEN_30607;
        end
      end else begin
        e_1_war_3 <= _GEN_30607;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_4 <= _GEN_30631;
        end
      end else begin
        e_1_war_4 <= _GEN_30631;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_5 <= _GEN_30655;
        end
      end else begin
        e_1_war_5 <= _GEN_30655;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_6 <= _GEN_30679;
        end
      end else begin
        e_1_war_6 <= _GEN_30679;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_1_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_1_war_7 <= _GEN_30703;
        end
      end else begin
        e_1_war_7 <= _GEN_30703;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_0 <= _GEN_30543;
        end
      end else begin
        e_1_waw_0 <= _GEN_30543;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_1 <= _GEN_30567;
        end
      end else begin
        e_1_waw_1 <= _GEN_30567;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_2 <= _GEN_30591;
        end
      end else begin
        e_1_waw_2 <= _GEN_30591;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_3 <= _GEN_30615;
        end
      end else begin
        e_1_waw_3 <= _GEN_30615;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_4 <= _GEN_30639;
        end
      end else begin
        e_1_waw_4 <= _GEN_30639;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_5 <= _GEN_30663;
        end
      end else begin
        e_1_waw_5 <= _GEN_30663;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_6 <= _GEN_30687;
        end
      end else begin
        e_1_waw_6 <= _GEN_30687;
      end
    end
    if (_GEN_32206) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_1_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_1_waw_7 <= _GEN_30711;
        end
      end else begin
        e_1_waw_7 <= _GEN_30711;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_1_last <= _GEN_31101;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_1_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_1_last <= _GEN_29197;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_1_last <= _GEN_27611;
      end else begin
        e_1_last <= _GEN_26113;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_1_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_1_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_1_rports <= _GEN_28917;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_1_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_1_rports <= _GEN_27075;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_rports <= _GEN_25769;
      end else begin
        e_1_rports <= _GEN_23887;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_1_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_1_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_1_wport_sram <= _GEN_28925;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_1_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_1_wport_sram <= _GEN_27083;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_wport_sram <= _GEN_25777;
      end else begin
        e_1_wport_sram <= _GEN_23895;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_1_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h1 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_1_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_1_wport_pred <= _GEN_28933;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h1 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_1_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_1_wport_pred <= _GEN_27091;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_1_wport_pred <= _GEN_25785;
      end else begin
        e_1_wport_pred <= _GEN_23903;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_2_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_2_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_2_fn_union <= _GEN_28702;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_2_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_2_fn_union <= _GEN_27068;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_fn_union <= _GEN_25330;
      end else begin
        e_2_fn_union <= _GEN_23800;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_2_sreg_ss1 <= _GEN_24514;
          end else begin
            e_2_sreg_ss1 <= _GEN_23880;
          end
        end else begin
          e_2_sreg_ss1 <= _GEN_23880;
        end
      end else begin
        e_2_sreg_ss1 <= _GEN_23880;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_2_sreg_ss2 <= _GEN_13526;
          end else begin
            e_2_sreg_ss2 <= _GEN_12652;
          end
        end else begin
          e_2_sreg_ss2 <= _GEN_12652;
        end
      end else begin
        e_2_sreg_ss2 <= _GEN_12652;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_2_sreg_ss3 <= _GEN_9170;
          end else begin
            e_2_sreg_ss3 <= _GEN_3748;
          end
        end else begin
          e_2_sreg_ss3 <= _GEN_3748;
        end
      end else begin
        e_2_sreg_ss3 <= _GEN_3748;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_2_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_2_base_vp_id <= _GEN_28750;
          end
        end else begin
          e_2_base_vp_id <= _GEN_28750;
        end
      end else begin
        e_2_base_vp_id <= _GEN_28308;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_2_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_2_base_vp_valid <= _GEN_29270;
          end
        end else begin
          e_2_base_vp_valid <= _GEN_29270;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_2_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_2_base_vp_valid <= _GEN_26804;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_base_vp_valid <= _GEN_25386;
      end else begin
        e_2_base_vp_valid <= _GEN_23536;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_2_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_2_base_vp_scalar <= _GEN_28766;
          end
        end else begin
          e_2_base_vp_scalar <= _GEN_28766;
        end
      end else begin
        e_2_base_vp_scalar <= _GEN_28316;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_2_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_2_base_vp_pred <= _GEN_28774;
          end
        end else begin
          e_2_base_vp_pred <= _GEN_28774;
        end
      end else begin
        e_2_base_vp_pred <= _GEN_28324;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_2_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_2_base_vs1_id <= _GEN_26178;
          end
        end else begin
          e_2_base_vs1_id <= _GEN_26178;
        end
      end else begin
        e_2_base_vs1_id <= _GEN_26178;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_2_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_2_base_vs1_valid <= _GEN_29278;
          end
        end else begin
          e_2_base_vs1_valid <= _GEN_29278;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_2_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_2_base_vs1_valid <= _GEN_26812;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_base_vs1_valid <= _GEN_25602;
      end else begin
        e_2_base_vs1_valid <= _GEN_23544;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_2_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_2_base_vs1_scalar <= _GEN_26186;
          end
        end else begin
          e_2_base_vs1_scalar <= _GEN_26186;
        end
      end else begin
        e_2_base_vs1_scalar <= _GEN_26186;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_2_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_2_base_vs1_pred <= _GEN_26194;
          end
        end else begin
          e_2_base_vs1_pred <= _GEN_26194;
        end
      end else begin
        e_2_base_vs1_pred <= _GEN_26194;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_2_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_2_base_vs1_prec <= _GEN_26202;
          end
        end else begin
          e_2_base_vs1_prec <= _GEN_26202;
        end
      end else begin
        e_2_base_vs1_prec <= _GEN_26202;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs2_id <= _GEN_12612;
          end
        end else begin
          e_2_base_vs2_id <= _GEN_12612;
        end
      end else begin
        e_2_base_vs2_id <= _GEN_12612;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_2_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_2_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_2_base_vs2_valid <= _GEN_28454;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_2_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_2_base_vs2_valid <= _GEN_26820;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_base_vs2_valid <= _GEN_25082;
      end else begin
        e_2_base_vs2_valid <= _GEN_23552;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs2_scalar <= _GEN_12620;
          end
        end else begin
          e_2_base_vs2_scalar <= _GEN_12620;
        end
      end else begin
        e_2_base_vs2_scalar <= _GEN_12620;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs2_pred <= _GEN_12628;
          end
        end else begin
          e_2_base_vs2_pred <= _GEN_12628;
        end
      end else begin
        e_2_base_vs2_pred <= _GEN_12628;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs2_prec <= _GEN_12636;
          end
        end else begin
          e_2_base_vs2_prec <= _GEN_12636;
        end
      end else begin
        e_2_base_vs2_prec <= _GEN_12636;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs3_id <= _GEN_3708;
          end
        end else begin
          e_2_base_vs3_id <= _GEN_3708;
        end
      end else begin
        e_2_base_vs3_id <= _GEN_3708;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_2_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_2_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_2_base_vs3_valid <= _GEN_28462;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_2_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_2_base_vs3_valid <= _GEN_26828;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_base_vs3_valid <= _GEN_25090;
      end else begin
        e_2_base_vs3_valid <= _GEN_23560;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs3_scalar <= _GEN_3716;
          end
        end else begin
          e_2_base_vs3_scalar <= _GEN_3716;
        end
      end else begin
        e_2_base_vs3_scalar <= _GEN_3716;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs3_pred <= _GEN_3724;
          end
        end else begin
          e_2_base_vs3_pred <= _GEN_3724;
        end
      end else begin
        e_2_base_vs3_pred <= _GEN_3724;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h2 == tail) begin // @[sequencer-master.scala 329:29]
            e_2_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_2_base_vs3_prec <= _GEN_3732;
          end
        end else begin
          e_2_base_vs3_prec <= _GEN_3732;
        end
      end else begin
        e_2_base_vs3_prec <= _GEN_3732;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_2_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_2_base_vd_id <= _GEN_23928;
          end
        end else begin
          e_2_base_vd_id <= _GEN_23928;
        end
      end else begin
        e_2_base_vd_id <= _GEN_23928;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_2_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_2_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_2_base_vd_valid <= _GEN_28470;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_2_base_vd_valid <= _GEN_27652;
        end else begin
          e_2_base_vd_valid <= _GEN_27404;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_base_vd_valid <= _GEN_25098;
      end else begin
        e_2_base_vd_valid <= _GEN_23568;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_2_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_2_base_vd_scalar <= _GEN_23936;
          end
        end else begin
          e_2_base_vd_scalar <= _GEN_23936;
        end
      end else begin
        e_2_base_vd_scalar <= _GEN_23936;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_2_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_2_base_vd_pred <= _GEN_23944;
          end
        end else begin
          e_2_base_vd_pred <= _GEN_23944;
        end
      end else begin
        e_2_base_vd_pred <= _GEN_23944;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h2 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_2_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_2_base_vd_prec <= _GEN_23952;
          end
        end else begin
          e_2_base_vd_prec <= _GEN_23952;
        end
      end else begin
        e_2_base_vd_prec <= _GEN_23952;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_viu <= _GEN_30736;
      end
    end else begin
      e_2_active_viu <= _GEN_30736;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vipu <= _GEN_30946;
      end
    end else begin
      e_2_active_vipu <= _GEN_30946;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vimu <= _GEN_31002;
      end
    end else begin
      e_2_active_vimu <= _GEN_31002;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vidu <= _GEN_31018;
      end
    end else begin
      e_2_active_vidu <= _GEN_31018;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vfmu <= _GEN_31026;
      end
    end else begin
      e_2_active_vfmu <= _GEN_31026;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vfdu <= _GEN_31034;
      end
    end else begin
      e_2_active_vfdu <= _GEN_31034;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vfcu <= _GEN_31042;
      end
    end else begin
      e_2_active_vfcu <= _GEN_31042;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vfvu <= _GEN_31050;
      end
    end else begin
      e_2_active_vfvu <= _GEN_31050;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vpu <= _GEN_31090;
      end
    end else begin
      e_2_active_vpu <= _GEN_31090;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vgu <= _GEN_31058;
      end
    end else begin
      e_2_active_vgu <= _GEN_31058;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vcu <= _GEN_31066;
      end
    end else begin
      e_2_active_vcu <= _GEN_31066;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vlu <= _GEN_31082;
      end
    end else begin
      e_2_active_vlu <= _GEN_31082;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vsu <= _GEN_31074;
      end
    end else begin
      e_2_active_vsu <= _GEN_31074;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_2_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h2 == head) begin // @[sequencer-master.scala 373:43]
        e_2_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_2_active_vqu <= _GEN_31010;
      end
    end else begin
      e_2_active_vqu <= _GEN_31010;
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_0 <= _GEN_30528;
        end
      end else begin
        e_2_raw_0 <= _GEN_30528;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_1 <= _GEN_30552;
        end
      end else begin
        e_2_raw_1 <= _GEN_30552;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_2 <= _GEN_30576;
        end
      end else begin
        e_2_raw_2 <= _GEN_30576;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_3 <= _GEN_30600;
        end
      end else begin
        e_2_raw_3 <= _GEN_30600;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_4 <= _GEN_30624;
        end
      end else begin
        e_2_raw_4 <= _GEN_30624;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_5 <= _GEN_30648;
        end
      end else begin
        e_2_raw_5 <= _GEN_30648;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_6 <= _GEN_30672;
        end
      end else begin
        e_2_raw_6 <= _GEN_30672;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_2_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_2_raw_7 <= _GEN_30696;
        end
      end else begin
        e_2_raw_7 <= _GEN_30696;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_0 <= _GEN_30536;
        end
      end else begin
        e_2_war_0 <= _GEN_30536;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_1 <= _GEN_30560;
        end
      end else begin
        e_2_war_1 <= _GEN_30560;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_2 <= _GEN_30584;
        end
      end else begin
        e_2_war_2 <= _GEN_30584;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_3 <= _GEN_30608;
        end
      end else begin
        e_2_war_3 <= _GEN_30608;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_4 <= _GEN_30632;
        end
      end else begin
        e_2_war_4 <= _GEN_30632;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_5 <= _GEN_30656;
        end
      end else begin
        e_2_war_5 <= _GEN_30656;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_6 <= _GEN_30680;
        end
      end else begin
        e_2_war_6 <= _GEN_30680;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_2_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_2_war_7 <= _GEN_30704;
        end
      end else begin
        e_2_war_7 <= _GEN_30704;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_0 <= _GEN_30544;
        end
      end else begin
        e_2_waw_0 <= _GEN_30544;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_1 <= _GEN_30568;
        end
      end else begin
        e_2_waw_1 <= _GEN_30568;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_2 <= _GEN_30592;
        end
      end else begin
        e_2_waw_2 <= _GEN_30592;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_3 <= _GEN_30616;
        end
      end else begin
        e_2_waw_3 <= _GEN_30616;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_4 <= _GEN_30640;
        end
      end else begin
        e_2_waw_4 <= _GEN_30640;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_5 <= _GEN_30664;
        end
      end else begin
        e_2_waw_5 <= _GEN_30664;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_6 <= _GEN_30688;
        end
      end else begin
        e_2_waw_6 <= _GEN_30688;
      end
    end
    if (_GEN_32231) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_2_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_2_waw_7 <= _GEN_30712;
        end
      end else begin
        e_2_waw_7 <= _GEN_30712;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_2_last <= _GEN_31102;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_2_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_2_last <= _GEN_29198;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_2_last <= _GEN_27612;
      end else begin
        e_2_last <= _GEN_26114;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_2_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_2_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_2_rports <= _GEN_28918;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_2_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_2_rports <= _GEN_27076;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_rports <= _GEN_25770;
      end else begin
        e_2_rports <= _GEN_23888;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_2_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_2_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_2_wport_sram <= _GEN_28926;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_2_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_2_wport_sram <= _GEN_27084;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_wport_sram <= _GEN_25778;
      end else begin
        e_2_wport_sram <= _GEN_23896;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_2_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h2 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_2_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_2_wport_pred <= _GEN_28934;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h2 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_2_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_2_wport_pred <= _GEN_27092;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_2_wport_pred <= _GEN_25786;
      end else begin
        e_2_wport_pred <= _GEN_23904;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_3_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_3_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_3_fn_union <= _GEN_28703;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_3_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_3_fn_union <= _GEN_27069;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_fn_union <= _GEN_25331;
      end else begin
        e_3_fn_union <= _GEN_23801;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_3_sreg_ss1 <= _GEN_24515;
          end else begin
            e_3_sreg_ss1 <= _GEN_23881;
          end
        end else begin
          e_3_sreg_ss1 <= _GEN_23881;
        end
      end else begin
        e_3_sreg_ss1 <= _GEN_23881;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_3_sreg_ss2 <= _GEN_13527;
          end else begin
            e_3_sreg_ss2 <= _GEN_12653;
          end
        end else begin
          e_3_sreg_ss2 <= _GEN_12653;
        end
      end else begin
        e_3_sreg_ss2 <= _GEN_12653;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_3_sreg_ss3 <= _GEN_9171;
          end else begin
            e_3_sreg_ss3 <= _GEN_3749;
          end
        end else begin
          e_3_sreg_ss3 <= _GEN_3749;
        end
      end else begin
        e_3_sreg_ss3 <= _GEN_3749;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_3_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_3_base_vp_id <= _GEN_28751;
          end
        end else begin
          e_3_base_vp_id <= _GEN_28751;
        end
      end else begin
        e_3_base_vp_id <= _GEN_28309;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_3_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_3_base_vp_valid <= _GEN_29271;
          end
        end else begin
          e_3_base_vp_valid <= _GEN_29271;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_3_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_3_base_vp_valid <= _GEN_26805;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_base_vp_valid <= _GEN_25387;
      end else begin
        e_3_base_vp_valid <= _GEN_23537;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_3_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_3_base_vp_scalar <= _GEN_28767;
          end
        end else begin
          e_3_base_vp_scalar <= _GEN_28767;
        end
      end else begin
        e_3_base_vp_scalar <= _GEN_28317;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_3_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_3_base_vp_pred <= _GEN_28775;
          end
        end else begin
          e_3_base_vp_pred <= _GEN_28775;
        end
      end else begin
        e_3_base_vp_pred <= _GEN_28325;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_3_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_3_base_vs1_id <= _GEN_26179;
          end
        end else begin
          e_3_base_vs1_id <= _GEN_26179;
        end
      end else begin
        e_3_base_vs1_id <= _GEN_26179;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_3_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_3_base_vs1_valid <= _GEN_29279;
          end
        end else begin
          e_3_base_vs1_valid <= _GEN_29279;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_3_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_3_base_vs1_valid <= _GEN_26813;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_base_vs1_valid <= _GEN_25603;
      end else begin
        e_3_base_vs1_valid <= _GEN_23545;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_3_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_3_base_vs1_scalar <= _GEN_26187;
          end
        end else begin
          e_3_base_vs1_scalar <= _GEN_26187;
        end
      end else begin
        e_3_base_vs1_scalar <= _GEN_26187;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_3_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_3_base_vs1_pred <= _GEN_26195;
          end
        end else begin
          e_3_base_vs1_pred <= _GEN_26195;
        end
      end else begin
        e_3_base_vs1_pred <= _GEN_26195;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_3_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_3_base_vs1_prec <= _GEN_26203;
          end
        end else begin
          e_3_base_vs1_prec <= _GEN_26203;
        end
      end else begin
        e_3_base_vs1_prec <= _GEN_26203;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs2_id <= _GEN_12613;
          end
        end else begin
          e_3_base_vs2_id <= _GEN_12613;
        end
      end else begin
        e_3_base_vs2_id <= _GEN_12613;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_3_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_3_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_3_base_vs2_valid <= _GEN_28455;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_3_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_3_base_vs2_valid <= _GEN_26821;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_base_vs2_valid <= _GEN_25083;
      end else begin
        e_3_base_vs2_valid <= _GEN_23553;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs2_scalar <= _GEN_12621;
          end
        end else begin
          e_3_base_vs2_scalar <= _GEN_12621;
        end
      end else begin
        e_3_base_vs2_scalar <= _GEN_12621;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs2_pred <= _GEN_12629;
          end
        end else begin
          e_3_base_vs2_pred <= _GEN_12629;
        end
      end else begin
        e_3_base_vs2_pred <= _GEN_12629;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs2_prec <= _GEN_12637;
          end
        end else begin
          e_3_base_vs2_prec <= _GEN_12637;
        end
      end else begin
        e_3_base_vs2_prec <= _GEN_12637;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs3_id <= _GEN_3709;
          end
        end else begin
          e_3_base_vs3_id <= _GEN_3709;
        end
      end else begin
        e_3_base_vs3_id <= _GEN_3709;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_3_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_3_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_3_base_vs3_valid <= _GEN_28463;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_3_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_3_base_vs3_valid <= _GEN_26829;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_base_vs3_valid <= _GEN_25091;
      end else begin
        e_3_base_vs3_valid <= _GEN_23561;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs3_scalar <= _GEN_3717;
          end
        end else begin
          e_3_base_vs3_scalar <= _GEN_3717;
        end
      end else begin
        e_3_base_vs3_scalar <= _GEN_3717;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs3_pred <= _GEN_3725;
          end
        end else begin
          e_3_base_vs3_pred <= _GEN_3725;
        end
      end else begin
        e_3_base_vs3_pred <= _GEN_3725;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h3 == tail) begin // @[sequencer-master.scala 329:29]
            e_3_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_3_base_vs3_prec <= _GEN_3733;
          end
        end else begin
          e_3_base_vs3_prec <= _GEN_3733;
        end
      end else begin
        e_3_base_vs3_prec <= _GEN_3733;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_3_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_3_base_vd_id <= _GEN_23929;
          end
        end else begin
          e_3_base_vd_id <= _GEN_23929;
        end
      end else begin
        e_3_base_vd_id <= _GEN_23929;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_3_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_3_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_3_base_vd_valid <= _GEN_28471;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_3_base_vd_valid <= _GEN_27653;
        end else begin
          e_3_base_vd_valid <= _GEN_27405;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_base_vd_valid <= _GEN_25099;
      end else begin
        e_3_base_vd_valid <= _GEN_23569;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_3_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_3_base_vd_scalar <= _GEN_23937;
          end
        end else begin
          e_3_base_vd_scalar <= _GEN_23937;
        end
      end else begin
        e_3_base_vd_scalar <= _GEN_23937;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_3_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_3_base_vd_pred <= _GEN_23945;
          end
        end else begin
          e_3_base_vd_pred <= _GEN_23945;
        end
      end else begin
        e_3_base_vd_pred <= _GEN_23945;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h3 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_3_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_3_base_vd_prec <= _GEN_23953;
          end
        end else begin
          e_3_base_vd_prec <= _GEN_23953;
        end
      end else begin
        e_3_base_vd_prec <= _GEN_23953;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_viu <= _GEN_30737;
      end
    end else begin
      e_3_active_viu <= _GEN_30737;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vipu <= _GEN_30947;
      end
    end else begin
      e_3_active_vipu <= _GEN_30947;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vimu <= _GEN_31003;
      end
    end else begin
      e_3_active_vimu <= _GEN_31003;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vidu <= _GEN_31019;
      end
    end else begin
      e_3_active_vidu <= _GEN_31019;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vfmu <= _GEN_31027;
      end
    end else begin
      e_3_active_vfmu <= _GEN_31027;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vfdu <= _GEN_31035;
      end
    end else begin
      e_3_active_vfdu <= _GEN_31035;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vfcu <= _GEN_31043;
      end
    end else begin
      e_3_active_vfcu <= _GEN_31043;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vfvu <= _GEN_31051;
      end
    end else begin
      e_3_active_vfvu <= _GEN_31051;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vpu <= _GEN_31091;
      end
    end else begin
      e_3_active_vpu <= _GEN_31091;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vgu <= _GEN_31059;
      end
    end else begin
      e_3_active_vgu <= _GEN_31059;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vcu <= _GEN_31067;
      end
    end else begin
      e_3_active_vcu <= _GEN_31067;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vlu <= _GEN_31083;
      end
    end else begin
      e_3_active_vlu <= _GEN_31083;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vsu <= _GEN_31075;
      end
    end else begin
      e_3_active_vsu <= _GEN_31075;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_3_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h3 == head) begin // @[sequencer-master.scala 373:43]
        e_3_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_3_active_vqu <= _GEN_31011;
      end
    end else begin
      e_3_active_vqu <= _GEN_31011;
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_0 <= _GEN_30529;
        end
      end else begin
        e_3_raw_0 <= _GEN_30529;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_1 <= _GEN_30553;
        end
      end else begin
        e_3_raw_1 <= _GEN_30553;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_2 <= _GEN_30577;
        end
      end else begin
        e_3_raw_2 <= _GEN_30577;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_3 <= _GEN_30601;
        end
      end else begin
        e_3_raw_3 <= _GEN_30601;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_4 <= _GEN_30625;
        end
      end else begin
        e_3_raw_4 <= _GEN_30625;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_5 <= _GEN_30649;
        end
      end else begin
        e_3_raw_5 <= _GEN_30649;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_6 <= _GEN_30673;
        end
      end else begin
        e_3_raw_6 <= _GEN_30673;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_3_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_3_raw_7 <= _GEN_30697;
        end
      end else begin
        e_3_raw_7 <= _GEN_30697;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_0 <= _GEN_30537;
        end
      end else begin
        e_3_war_0 <= _GEN_30537;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_1 <= _GEN_30561;
        end
      end else begin
        e_3_war_1 <= _GEN_30561;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_2 <= _GEN_30585;
        end
      end else begin
        e_3_war_2 <= _GEN_30585;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_3 <= _GEN_30609;
        end
      end else begin
        e_3_war_3 <= _GEN_30609;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_4 <= _GEN_30633;
        end
      end else begin
        e_3_war_4 <= _GEN_30633;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_5 <= _GEN_30657;
        end
      end else begin
        e_3_war_5 <= _GEN_30657;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_6 <= _GEN_30681;
        end
      end else begin
        e_3_war_6 <= _GEN_30681;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_3_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_3_war_7 <= _GEN_30705;
        end
      end else begin
        e_3_war_7 <= _GEN_30705;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_0 <= _GEN_30545;
        end
      end else begin
        e_3_waw_0 <= _GEN_30545;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_1 <= _GEN_30569;
        end
      end else begin
        e_3_waw_1 <= _GEN_30569;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_2 <= _GEN_30593;
        end
      end else begin
        e_3_waw_2 <= _GEN_30593;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_3 <= _GEN_30617;
        end
      end else begin
        e_3_waw_3 <= _GEN_30617;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_4 <= _GEN_30641;
        end
      end else begin
        e_3_waw_4 <= _GEN_30641;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_5 <= _GEN_30665;
        end
      end else begin
        e_3_waw_5 <= _GEN_30665;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_6 <= _GEN_30689;
        end
      end else begin
        e_3_waw_6 <= _GEN_30689;
      end
    end
    if (_GEN_32256) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_3_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_3_waw_7 <= _GEN_30713;
        end
      end else begin
        e_3_waw_7 <= _GEN_30713;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_3_last <= _GEN_31103;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_3_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_3_last <= _GEN_29199;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_3_last <= _GEN_27613;
      end else begin
        e_3_last <= _GEN_26115;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_3_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_3_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_3_rports <= _GEN_28919;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_3_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_3_rports <= _GEN_27077;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_rports <= _GEN_25771;
      end else begin
        e_3_rports <= _GEN_23889;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_3_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_3_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_3_wport_sram <= _GEN_28927;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_3_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_3_wport_sram <= _GEN_27085;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_wport_sram <= _GEN_25779;
      end else begin
        e_3_wport_sram <= _GEN_23897;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_3_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h3 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_3_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_3_wport_pred <= _GEN_28935;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h3 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_3_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_3_wport_pred <= _GEN_27093;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_3_wport_pred <= _GEN_25787;
      end else begin
        e_3_wport_pred <= _GEN_23905;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_4_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_4_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_4_fn_union <= _GEN_28704;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_4_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_4_fn_union <= _GEN_27070;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_fn_union <= _GEN_25332;
      end else begin
        e_4_fn_union <= _GEN_23802;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_4_sreg_ss1 <= _GEN_24516;
          end else begin
            e_4_sreg_ss1 <= _GEN_23882;
          end
        end else begin
          e_4_sreg_ss1 <= _GEN_23882;
        end
      end else begin
        e_4_sreg_ss1 <= _GEN_23882;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_4_sreg_ss2 <= _GEN_13528;
          end else begin
            e_4_sreg_ss2 <= _GEN_12654;
          end
        end else begin
          e_4_sreg_ss2 <= _GEN_12654;
        end
      end else begin
        e_4_sreg_ss2 <= _GEN_12654;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_4_sreg_ss3 <= _GEN_9172;
          end else begin
            e_4_sreg_ss3 <= _GEN_3750;
          end
        end else begin
          e_4_sreg_ss3 <= _GEN_3750;
        end
      end else begin
        e_4_sreg_ss3 <= _GEN_3750;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_4_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_4_base_vp_id <= _GEN_28752;
          end
        end else begin
          e_4_base_vp_id <= _GEN_28752;
        end
      end else begin
        e_4_base_vp_id <= _GEN_28310;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_4_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_4_base_vp_valid <= _GEN_29272;
          end
        end else begin
          e_4_base_vp_valid <= _GEN_29272;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_4_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_4_base_vp_valid <= _GEN_26806;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_base_vp_valid <= _GEN_25388;
      end else begin
        e_4_base_vp_valid <= _GEN_23538;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_4_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_4_base_vp_scalar <= _GEN_28768;
          end
        end else begin
          e_4_base_vp_scalar <= _GEN_28768;
        end
      end else begin
        e_4_base_vp_scalar <= _GEN_28318;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_4_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_4_base_vp_pred <= _GEN_28776;
          end
        end else begin
          e_4_base_vp_pred <= _GEN_28776;
        end
      end else begin
        e_4_base_vp_pred <= _GEN_28326;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_4_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_4_base_vs1_id <= _GEN_26180;
          end
        end else begin
          e_4_base_vs1_id <= _GEN_26180;
        end
      end else begin
        e_4_base_vs1_id <= _GEN_26180;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_4_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_4_base_vs1_valid <= _GEN_29280;
          end
        end else begin
          e_4_base_vs1_valid <= _GEN_29280;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_4_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_4_base_vs1_valid <= _GEN_26814;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_base_vs1_valid <= _GEN_25604;
      end else begin
        e_4_base_vs1_valid <= _GEN_23546;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_4_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_4_base_vs1_scalar <= _GEN_26188;
          end
        end else begin
          e_4_base_vs1_scalar <= _GEN_26188;
        end
      end else begin
        e_4_base_vs1_scalar <= _GEN_26188;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_4_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_4_base_vs1_pred <= _GEN_26196;
          end
        end else begin
          e_4_base_vs1_pred <= _GEN_26196;
        end
      end else begin
        e_4_base_vs1_pred <= _GEN_26196;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_4_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_4_base_vs1_prec <= _GEN_26204;
          end
        end else begin
          e_4_base_vs1_prec <= _GEN_26204;
        end
      end else begin
        e_4_base_vs1_prec <= _GEN_26204;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs2_id <= _GEN_12614;
          end
        end else begin
          e_4_base_vs2_id <= _GEN_12614;
        end
      end else begin
        e_4_base_vs2_id <= _GEN_12614;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_4_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_4_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_4_base_vs2_valid <= _GEN_28456;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_4_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_4_base_vs2_valid <= _GEN_26822;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_base_vs2_valid <= _GEN_25084;
      end else begin
        e_4_base_vs2_valid <= _GEN_23554;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs2_scalar <= _GEN_12622;
          end
        end else begin
          e_4_base_vs2_scalar <= _GEN_12622;
        end
      end else begin
        e_4_base_vs2_scalar <= _GEN_12622;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs2_pred <= _GEN_12630;
          end
        end else begin
          e_4_base_vs2_pred <= _GEN_12630;
        end
      end else begin
        e_4_base_vs2_pred <= _GEN_12630;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs2_prec <= _GEN_12638;
          end
        end else begin
          e_4_base_vs2_prec <= _GEN_12638;
        end
      end else begin
        e_4_base_vs2_prec <= _GEN_12638;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs3_id <= _GEN_3710;
          end
        end else begin
          e_4_base_vs3_id <= _GEN_3710;
        end
      end else begin
        e_4_base_vs3_id <= _GEN_3710;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_4_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_4_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_4_base_vs3_valid <= _GEN_28464;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_4_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_4_base_vs3_valid <= _GEN_26830;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_base_vs3_valid <= _GEN_25092;
      end else begin
        e_4_base_vs3_valid <= _GEN_23562;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs3_scalar <= _GEN_3718;
          end
        end else begin
          e_4_base_vs3_scalar <= _GEN_3718;
        end
      end else begin
        e_4_base_vs3_scalar <= _GEN_3718;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs3_pred <= _GEN_3726;
          end
        end else begin
          e_4_base_vs3_pred <= _GEN_3726;
        end
      end else begin
        e_4_base_vs3_pred <= _GEN_3726;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h4 == tail) begin // @[sequencer-master.scala 329:29]
            e_4_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_4_base_vs3_prec <= _GEN_3734;
          end
        end else begin
          e_4_base_vs3_prec <= _GEN_3734;
        end
      end else begin
        e_4_base_vs3_prec <= _GEN_3734;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_4_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_4_base_vd_id <= _GEN_23930;
          end
        end else begin
          e_4_base_vd_id <= _GEN_23930;
        end
      end else begin
        e_4_base_vd_id <= _GEN_23930;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_4_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_4_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_4_base_vd_valid <= _GEN_28472;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_4_base_vd_valid <= _GEN_27654;
        end else begin
          e_4_base_vd_valid <= _GEN_27406;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_base_vd_valid <= _GEN_25100;
      end else begin
        e_4_base_vd_valid <= _GEN_23570;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_4_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_4_base_vd_scalar <= _GEN_23938;
          end
        end else begin
          e_4_base_vd_scalar <= _GEN_23938;
        end
      end else begin
        e_4_base_vd_scalar <= _GEN_23938;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_4_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_4_base_vd_pred <= _GEN_23946;
          end
        end else begin
          e_4_base_vd_pred <= _GEN_23946;
        end
      end else begin
        e_4_base_vd_pred <= _GEN_23946;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h4 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_4_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_4_base_vd_prec <= _GEN_23954;
          end
        end else begin
          e_4_base_vd_prec <= _GEN_23954;
        end
      end else begin
        e_4_base_vd_prec <= _GEN_23954;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_viu <= _GEN_30738;
      end
    end else begin
      e_4_active_viu <= _GEN_30738;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vipu <= _GEN_30948;
      end
    end else begin
      e_4_active_vipu <= _GEN_30948;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vimu <= _GEN_31004;
      end
    end else begin
      e_4_active_vimu <= _GEN_31004;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vidu <= _GEN_31020;
      end
    end else begin
      e_4_active_vidu <= _GEN_31020;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vfmu <= _GEN_31028;
      end
    end else begin
      e_4_active_vfmu <= _GEN_31028;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vfdu <= _GEN_31036;
      end
    end else begin
      e_4_active_vfdu <= _GEN_31036;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vfcu <= _GEN_31044;
      end
    end else begin
      e_4_active_vfcu <= _GEN_31044;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vfvu <= _GEN_31052;
      end
    end else begin
      e_4_active_vfvu <= _GEN_31052;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vpu <= _GEN_31092;
      end
    end else begin
      e_4_active_vpu <= _GEN_31092;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vgu <= _GEN_31060;
      end
    end else begin
      e_4_active_vgu <= _GEN_31060;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vcu <= _GEN_31068;
      end
    end else begin
      e_4_active_vcu <= _GEN_31068;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vlu <= _GEN_31084;
      end
    end else begin
      e_4_active_vlu <= _GEN_31084;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vsu <= _GEN_31076;
      end
    end else begin
      e_4_active_vsu <= _GEN_31076;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_4_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h4 == head) begin // @[sequencer-master.scala 373:43]
        e_4_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_4_active_vqu <= _GEN_31012;
      end
    end else begin
      e_4_active_vqu <= _GEN_31012;
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_0 <= _GEN_30530;
        end
      end else begin
        e_4_raw_0 <= _GEN_30530;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_1 <= _GEN_30554;
        end
      end else begin
        e_4_raw_1 <= _GEN_30554;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_2 <= _GEN_30578;
        end
      end else begin
        e_4_raw_2 <= _GEN_30578;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_3 <= _GEN_30602;
        end
      end else begin
        e_4_raw_3 <= _GEN_30602;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_4 <= _GEN_30626;
        end
      end else begin
        e_4_raw_4 <= _GEN_30626;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_5 <= _GEN_30650;
        end
      end else begin
        e_4_raw_5 <= _GEN_30650;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_6 <= _GEN_30674;
        end
      end else begin
        e_4_raw_6 <= _GEN_30674;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_4_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_4_raw_7 <= _GEN_30698;
        end
      end else begin
        e_4_raw_7 <= _GEN_30698;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_0 <= _GEN_30538;
        end
      end else begin
        e_4_war_0 <= _GEN_30538;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_1 <= _GEN_30562;
        end
      end else begin
        e_4_war_1 <= _GEN_30562;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_2 <= _GEN_30586;
        end
      end else begin
        e_4_war_2 <= _GEN_30586;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_3 <= _GEN_30610;
        end
      end else begin
        e_4_war_3 <= _GEN_30610;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_4 <= _GEN_30634;
        end
      end else begin
        e_4_war_4 <= _GEN_30634;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_5 <= _GEN_30658;
        end
      end else begin
        e_4_war_5 <= _GEN_30658;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_6 <= _GEN_30682;
        end
      end else begin
        e_4_war_6 <= _GEN_30682;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_4_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_4_war_7 <= _GEN_30706;
        end
      end else begin
        e_4_war_7 <= _GEN_30706;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_0 <= _GEN_30546;
        end
      end else begin
        e_4_waw_0 <= _GEN_30546;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_1 <= _GEN_30570;
        end
      end else begin
        e_4_waw_1 <= _GEN_30570;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_2 <= _GEN_30594;
        end
      end else begin
        e_4_waw_2 <= _GEN_30594;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_3 <= _GEN_30618;
        end
      end else begin
        e_4_waw_3 <= _GEN_30618;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_4 <= _GEN_30642;
        end
      end else begin
        e_4_waw_4 <= _GEN_30642;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_5 <= _GEN_30666;
        end
      end else begin
        e_4_waw_5 <= _GEN_30666;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_6 <= _GEN_30690;
        end
      end else begin
        e_4_waw_6 <= _GEN_30690;
      end
    end
    if (_GEN_32281) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_4_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_4_waw_7 <= _GEN_30714;
        end
      end else begin
        e_4_waw_7 <= _GEN_30714;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_4_last <= _GEN_31104;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_4_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_4_last <= _GEN_29200;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_4_last <= _GEN_27614;
      end else begin
        e_4_last <= _GEN_26116;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_4_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_4_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_4_rports <= _GEN_28920;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_4_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_4_rports <= _GEN_27078;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_rports <= _GEN_25772;
      end else begin
        e_4_rports <= _GEN_23890;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_4_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_4_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_4_wport_sram <= _GEN_28928;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_4_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_4_wport_sram <= _GEN_27086;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_wport_sram <= _GEN_25780;
      end else begin
        e_4_wport_sram <= _GEN_23898;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_4_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h4 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_4_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_4_wport_pred <= _GEN_28936;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h4 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_4_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_4_wport_pred <= _GEN_27094;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_4_wport_pred <= _GEN_25788;
      end else begin
        e_4_wport_pred <= _GEN_23906;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_5_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_5_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_5_fn_union <= _GEN_28705;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_5_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_5_fn_union <= _GEN_27071;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_fn_union <= _GEN_25333;
      end else begin
        e_5_fn_union <= _GEN_23803;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_5_sreg_ss1 <= _GEN_24517;
          end else begin
            e_5_sreg_ss1 <= _GEN_23883;
          end
        end else begin
          e_5_sreg_ss1 <= _GEN_23883;
        end
      end else begin
        e_5_sreg_ss1 <= _GEN_23883;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_5_sreg_ss2 <= _GEN_13529;
          end else begin
            e_5_sreg_ss2 <= _GEN_12655;
          end
        end else begin
          e_5_sreg_ss2 <= _GEN_12655;
        end
      end else begin
        e_5_sreg_ss2 <= _GEN_12655;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_5_sreg_ss3 <= _GEN_9173;
          end else begin
            e_5_sreg_ss3 <= _GEN_3751;
          end
        end else begin
          e_5_sreg_ss3 <= _GEN_3751;
        end
      end else begin
        e_5_sreg_ss3 <= _GEN_3751;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_5_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_5_base_vp_id <= _GEN_28753;
          end
        end else begin
          e_5_base_vp_id <= _GEN_28753;
        end
      end else begin
        e_5_base_vp_id <= _GEN_28311;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_5_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_5_base_vp_valid <= _GEN_29273;
          end
        end else begin
          e_5_base_vp_valid <= _GEN_29273;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_5_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_5_base_vp_valid <= _GEN_26807;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_base_vp_valid <= _GEN_25389;
      end else begin
        e_5_base_vp_valid <= _GEN_23539;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_5_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_5_base_vp_scalar <= _GEN_28769;
          end
        end else begin
          e_5_base_vp_scalar <= _GEN_28769;
        end
      end else begin
        e_5_base_vp_scalar <= _GEN_28319;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_5_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_5_base_vp_pred <= _GEN_28777;
          end
        end else begin
          e_5_base_vp_pred <= _GEN_28777;
        end
      end else begin
        e_5_base_vp_pred <= _GEN_28327;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_5_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_5_base_vs1_id <= _GEN_26181;
          end
        end else begin
          e_5_base_vs1_id <= _GEN_26181;
        end
      end else begin
        e_5_base_vs1_id <= _GEN_26181;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_5_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_5_base_vs1_valid <= _GEN_29281;
          end
        end else begin
          e_5_base_vs1_valid <= _GEN_29281;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_5_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_5_base_vs1_valid <= _GEN_26815;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_base_vs1_valid <= _GEN_25605;
      end else begin
        e_5_base_vs1_valid <= _GEN_23547;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_5_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_5_base_vs1_scalar <= _GEN_26189;
          end
        end else begin
          e_5_base_vs1_scalar <= _GEN_26189;
        end
      end else begin
        e_5_base_vs1_scalar <= _GEN_26189;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_5_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_5_base_vs1_pred <= _GEN_26197;
          end
        end else begin
          e_5_base_vs1_pred <= _GEN_26197;
        end
      end else begin
        e_5_base_vs1_pred <= _GEN_26197;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_5_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_5_base_vs1_prec <= _GEN_26205;
          end
        end else begin
          e_5_base_vs1_prec <= _GEN_26205;
        end
      end else begin
        e_5_base_vs1_prec <= _GEN_26205;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs2_id <= _GEN_12615;
          end
        end else begin
          e_5_base_vs2_id <= _GEN_12615;
        end
      end else begin
        e_5_base_vs2_id <= _GEN_12615;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_5_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_5_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_5_base_vs2_valid <= _GEN_28457;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_5_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_5_base_vs2_valid <= _GEN_26823;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_base_vs2_valid <= _GEN_25085;
      end else begin
        e_5_base_vs2_valid <= _GEN_23555;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs2_scalar <= _GEN_12623;
          end
        end else begin
          e_5_base_vs2_scalar <= _GEN_12623;
        end
      end else begin
        e_5_base_vs2_scalar <= _GEN_12623;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs2_pred <= _GEN_12631;
          end
        end else begin
          e_5_base_vs2_pred <= _GEN_12631;
        end
      end else begin
        e_5_base_vs2_pred <= _GEN_12631;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs2_prec <= _GEN_12639;
          end
        end else begin
          e_5_base_vs2_prec <= _GEN_12639;
        end
      end else begin
        e_5_base_vs2_prec <= _GEN_12639;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs3_id <= _GEN_3711;
          end
        end else begin
          e_5_base_vs3_id <= _GEN_3711;
        end
      end else begin
        e_5_base_vs3_id <= _GEN_3711;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_5_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_5_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_5_base_vs3_valid <= _GEN_28465;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_5_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_5_base_vs3_valid <= _GEN_26831;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_base_vs3_valid <= _GEN_25093;
      end else begin
        e_5_base_vs3_valid <= _GEN_23563;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs3_scalar <= _GEN_3719;
          end
        end else begin
          e_5_base_vs3_scalar <= _GEN_3719;
        end
      end else begin
        e_5_base_vs3_scalar <= _GEN_3719;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs3_pred <= _GEN_3727;
          end
        end else begin
          e_5_base_vs3_pred <= _GEN_3727;
        end
      end else begin
        e_5_base_vs3_pred <= _GEN_3727;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h5 == tail) begin // @[sequencer-master.scala 329:29]
            e_5_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_5_base_vs3_prec <= _GEN_3735;
          end
        end else begin
          e_5_base_vs3_prec <= _GEN_3735;
        end
      end else begin
        e_5_base_vs3_prec <= _GEN_3735;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_5_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_5_base_vd_id <= _GEN_23931;
          end
        end else begin
          e_5_base_vd_id <= _GEN_23931;
        end
      end else begin
        e_5_base_vd_id <= _GEN_23931;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_5_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_5_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_5_base_vd_valid <= _GEN_28473;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_5_base_vd_valid <= _GEN_27655;
        end else begin
          e_5_base_vd_valid <= _GEN_27407;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_base_vd_valid <= _GEN_25101;
      end else begin
        e_5_base_vd_valid <= _GEN_23571;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_5_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_5_base_vd_scalar <= _GEN_23939;
          end
        end else begin
          e_5_base_vd_scalar <= _GEN_23939;
        end
      end else begin
        e_5_base_vd_scalar <= _GEN_23939;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_5_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_5_base_vd_pred <= _GEN_23947;
          end
        end else begin
          e_5_base_vd_pred <= _GEN_23947;
        end
      end else begin
        e_5_base_vd_pred <= _GEN_23947;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h5 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_5_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_5_base_vd_prec <= _GEN_23955;
          end
        end else begin
          e_5_base_vd_prec <= _GEN_23955;
        end
      end else begin
        e_5_base_vd_prec <= _GEN_23955;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_viu <= _GEN_30739;
      end
    end else begin
      e_5_active_viu <= _GEN_30739;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vipu <= _GEN_30949;
      end
    end else begin
      e_5_active_vipu <= _GEN_30949;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vimu <= _GEN_31005;
      end
    end else begin
      e_5_active_vimu <= _GEN_31005;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vidu <= _GEN_31021;
      end
    end else begin
      e_5_active_vidu <= _GEN_31021;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vfmu <= _GEN_31029;
      end
    end else begin
      e_5_active_vfmu <= _GEN_31029;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vfdu <= _GEN_31037;
      end
    end else begin
      e_5_active_vfdu <= _GEN_31037;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vfcu <= _GEN_31045;
      end
    end else begin
      e_5_active_vfcu <= _GEN_31045;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vfvu <= _GEN_31053;
      end
    end else begin
      e_5_active_vfvu <= _GEN_31053;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vpu <= _GEN_31093;
      end
    end else begin
      e_5_active_vpu <= _GEN_31093;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vgu <= _GEN_31061;
      end
    end else begin
      e_5_active_vgu <= _GEN_31061;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vcu <= _GEN_31069;
      end
    end else begin
      e_5_active_vcu <= _GEN_31069;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vlu <= _GEN_31085;
      end
    end else begin
      e_5_active_vlu <= _GEN_31085;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vsu <= _GEN_31077;
      end
    end else begin
      e_5_active_vsu <= _GEN_31077;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_5_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h5 == head) begin // @[sequencer-master.scala 373:43]
        e_5_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_5_active_vqu <= _GEN_31013;
      end
    end else begin
      e_5_active_vqu <= _GEN_31013;
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_0 <= _GEN_30531;
        end
      end else begin
        e_5_raw_0 <= _GEN_30531;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_1 <= _GEN_30555;
        end
      end else begin
        e_5_raw_1 <= _GEN_30555;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_2 <= _GEN_30579;
        end
      end else begin
        e_5_raw_2 <= _GEN_30579;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_3 <= _GEN_30603;
        end
      end else begin
        e_5_raw_3 <= _GEN_30603;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_4 <= _GEN_30627;
        end
      end else begin
        e_5_raw_4 <= _GEN_30627;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_5 <= _GEN_30651;
        end
      end else begin
        e_5_raw_5 <= _GEN_30651;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_6 <= _GEN_30675;
        end
      end else begin
        e_5_raw_6 <= _GEN_30675;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_5_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_5_raw_7 <= _GEN_30699;
        end
      end else begin
        e_5_raw_7 <= _GEN_30699;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_0 <= _GEN_30539;
        end
      end else begin
        e_5_war_0 <= _GEN_30539;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_1 <= _GEN_30563;
        end
      end else begin
        e_5_war_1 <= _GEN_30563;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_2 <= _GEN_30587;
        end
      end else begin
        e_5_war_2 <= _GEN_30587;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_3 <= _GEN_30611;
        end
      end else begin
        e_5_war_3 <= _GEN_30611;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_4 <= _GEN_30635;
        end
      end else begin
        e_5_war_4 <= _GEN_30635;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_5 <= _GEN_30659;
        end
      end else begin
        e_5_war_5 <= _GEN_30659;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_6 <= _GEN_30683;
        end
      end else begin
        e_5_war_6 <= _GEN_30683;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_5_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_5_war_7 <= _GEN_30707;
        end
      end else begin
        e_5_war_7 <= _GEN_30707;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_0 <= _GEN_30547;
        end
      end else begin
        e_5_waw_0 <= _GEN_30547;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_1 <= _GEN_30571;
        end
      end else begin
        e_5_waw_1 <= _GEN_30571;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_2 <= _GEN_30595;
        end
      end else begin
        e_5_waw_2 <= _GEN_30595;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_3 <= _GEN_30619;
        end
      end else begin
        e_5_waw_3 <= _GEN_30619;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_4 <= _GEN_30643;
        end
      end else begin
        e_5_waw_4 <= _GEN_30643;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_5 <= _GEN_30667;
        end
      end else begin
        e_5_waw_5 <= _GEN_30667;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_6 <= _GEN_30691;
        end
      end else begin
        e_5_waw_6 <= _GEN_30691;
      end
    end
    if (_GEN_32306) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_5_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_5_waw_7 <= _GEN_30715;
        end
      end else begin
        e_5_waw_7 <= _GEN_30715;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_5_last <= _GEN_31105;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_5_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_5_last <= _GEN_29201;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_5_last <= _GEN_27615;
      end else begin
        e_5_last <= _GEN_26117;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_5_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_5_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_5_rports <= _GEN_28921;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_5_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_5_rports <= _GEN_27079;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_rports <= _GEN_25773;
      end else begin
        e_5_rports <= _GEN_23891;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_5_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_5_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_5_wport_sram <= _GEN_28929;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_5_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_5_wport_sram <= _GEN_27087;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_wport_sram <= _GEN_25781;
      end else begin
        e_5_wport_sram <= _GEN_23899;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_5_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h5 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_5_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_5_wport_pred <= _GEN_28937;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h5 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_5_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_5_wport_pred <= _GEN_27095;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_5_wport_pred <= _GEN_25789;
      end else begin
        e_5_wport_pred <= _GEN_23907;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_6_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_6_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_6_fn_union <= _GEN_28706;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_6_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_6_fn_union <= _GEN_27072;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_fn_union <= _GEN_25334;
      end else begin
        e_6_fn_union <= _GEN_23804;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_6_sreg_ss1 <= _GEN_24518;
          end else begin
            e_6_sreg_ss1 <= _GEN_23884;
          end
        end else begin
          e_6_sreg_ss1 <= _GEN_23884;
        end
      end else begin
        e_6_sreg_ss1 <= _GEN_23884;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_6_sreg_ss2 <= _GEN_13530;
          end else begin
            e_6_sreg_ss2 <= _GEN_12656;
          end
        end else begin
          e_6_sreg_ss2 <= _GEN_12656;
        end
      end else begin
        e_6_sreg_ss2 <= _GEN_12656;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_6_sreg_ss3 <= _GEN_9174;
          end else begin
            e_6_sreg_ss3 <= _GEN_3752;
          end
        end else begin
          e_6_sreg_ss3 <= _GEN_3752;
        end
      end else begin
        e_6_sreg_ss3 <= _GEN_3752;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_6_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_6_base_vp_id <= _GEN_28754;
          end
        end else begin
          e_6_base_vp_id <= _GEN_28754;
        end
      end else begin
        e_6_base_vp_id <= _GEN_28312;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_6_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_6_base_vp_valid <= _GEN_29274;
          end
        end else begin
          e_6_base_vp_valid <= _GEN_29274;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_6_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_6_base_vp_valid <= _GEN_26808;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_base_vp_valid <= _GEN_25390;
      end else begin
        e_6_base_vp_valid <= _GEN_23540;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_6_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_6_base_vp_scalar <= _GEN_28770;
          end
        end else begin
          e_6_base_vp_scalar <= _GEN_28770;
        end
      end else begin
        e_6_base_vp_scalar <= _GEN_28320;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_6_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_6_base_vp_pred <= _GEN_28778;
          end
        end else begin
          e_6_base_vp_pred <= _GEN_28778;
        end
      end else begin
        e_6_base_vp_pred <= _GEN_28328;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_6_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_6_base_vs1_id <= _GEN_26182;
          end
        end else begin
          e_6_base_vs1_id <= _GEN_26182;
        end
      end else begin
        e_6_base_vs1_id <= _GEN_26182;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_6_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_6_base_vs1_valid <= _GEN_29282;
          end
        end else begin
          e_6_base_vs1_valid <= _GEN_29282;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_6_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_6_base_vs1_valid <= _GEN_26816;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_base_vs1_valid <= _GEN_25606;
      end else begin
        e_6_base_vs1_valid <= _GEN_23548;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_6_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_6_base_vs1_scalar <= _GEN_26190;
          end
        end else begin
          e_6_base_vs1_scalar <= _GEN_26190;
        end
      end else begin
        e_6_base_vs1_scalar <= _GEN_26190;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_6_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_6_base_vs1_pred <= _GEN_26198;
          end
        end else begin
          e_6_base_vs1_pred <= _GEN_26198;
        end
      end else begin
        e_6_base_vs1_pred <= _GEN_26198;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_6_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_6_base_vs1_prec <= _GEN_26206;
          end
        end else begin
          e_6_base_vs1_prec <= _GEN_26206;
        end
      end else begin
        e_6_base_vs1_prec <= _GEN_26206;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs2_id <= _GEN_12616;
          end
        end else begin
          e_6_base_vs2_id <= _GEN_12616;
        end
      end else begin
        e_6_base_vs2_id <= _GEN_12616;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_6_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_6_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_6_base_vs2_valid <= _GEN_28458;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_6_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_6_base_vs2_valid <= _GEN_26824;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_base_vs2_valid <= _GEN_25086;
      end else begin
        e_6_base_vs2_valid <= _GEN_23556;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs2_scalar <= _GEN_12624;
          end
        end else begin
          e_6_base_vs2_scalar <= _GEN_12624;
        end
      end else begin
        e_6_base_vs2_scalar <= _GEN_12624;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs2_pred <= _GEN_12632;
          end
        end else begin
          e_6_base_vs2_pred <= _GEN_12632;
        end
      end else begin
        e_6_base_vs2_pred <= _GEN_12632;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs2_prec <= _GEN_12640;
          end
        end else begin
          e_6_base_vs2_prec <= _GEN_12640;
        end
      end else begin
        e_6_base_vs2_prec <= _GEN_12640;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs3_id <= _GEN_3712;
          end
        end else begin
          e_6_base_vs3_id <= _GEN_3712;
        end
      end else begin
        e_6_base_vs3_id <= _GEN_3712;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_6_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_6_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_6_base_vs3_valid <= _GEN_28466;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_6_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_6_base_vs3_valid <= _GEN_26832;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_base_vs3_valid <= _GEN_25094;
      end else begin
        e_6_base_vs3_valid <= _GEN_23564;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs3_scalar <= _GEN_3720;
          end
        end else begin
          e_6_base_vs3_scalar <= _GEN_3720;
        end
      end else begin
        e_6_base_vs3_scalar <= _GEN_3720;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs3_pred <= _GEN_3728;
          end
        end else begin
          e_6_base_vs3_pred <= _GEN_3728;
        end
      end else begin
        e_6_base_vs3_pred <= _GEN_3728;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h6 == tail) begin // @[sequencer-master.scala 329:29]
            e_6_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_6_base_vs3_prec <= _GEN_3736;
          end
        end else begin
          e_6_base_vs3_prec <= _GEN_3736;
        end
      end else begin
        e_6_base_vs3_prec <= _GEN_3736;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_6_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_6_base_vd_id <= _GEN_23932;
          end
        end else begin
          e_6_base_vd_id <= _GEN_23932;
        end
      end else begin
        e_6_base_vd_id <= _GEN_23932;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_6_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_6_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_6_base_vd_valid <= _GEN_28474;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_6_base_vd_valid <= _GEN_27656;
        end else begin
          e_6_base_vd_valid <= _GEN_27408;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_base_vd_valid <= _GEN_25102;
      end else begin
        e_6_base_vd_valid <= _GEN_23572;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_6_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_6_base_vd_scalar <= _GEN_23940;
          end
        end else begin
          e_6_base_vd_scalar <= _GEN_23940;
        end
      end else begin
        e_6_base_vd_scalar <= _GEN_23940;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_6_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_6_base_vd_pred <= _GEN_23948;
          end
        end else begin
          e_6_base_vd_pred <= _GEN_23948;
        end
      end else begin
        e_6_base_vd_pred <= _GEN_23948;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h6 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_6_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_6_base_vd_prec <= _GEN_23956;
          end
        end else begin
          e_6_base_vd_prec <= _GEN_23956;
        end
      end else begin
        e_6_base_vd_prec <= _GEN_23956;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_viu <= _GEN_30740;
      end
    end else begin
      e_6_active_viu <= _GEN_30740;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vipu <= _GEN_30950;
      end
    end else begin
      e_6_active_vipu <= _GEN_30950;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vimu <= _GEN_31006;
      end
    end else begin
      e_6_active_vimu <= _GEN_31006;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vidu <= _GEN_31022;
      end
    end else begin
      e_6_active_vidu <= _GEN_31022;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vfmu <= _GEN_31030;
      end
    end else begin
      e_6_active_vfmu <= _GEN_31030;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vfdu <= _GEN_31038;
      end
    end else begin
      e_6_active_vfdu <= _GEN_31038;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vfcu <= _GEN_31046;
      end
    end else begin
      e_6_active_vfcu <= _GEN_31046;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vfvu <= _GEN_31054;
      end
    end else begin
      e_6_active_vfvu <= _GEN_31054;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vpu <= _GEN_31094;
      end
    end else begin
      e_6_active_vpu <= _GEN_31094;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vgu <= _GEN_31062;
      end
    end else begin
      e_6_active_vgu <= _GEN_31062;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vcu <= _GEN_31070;
      end
    end else begin
      e_6_active_vcu <= _GEN_31070;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vlu <= _GEN_31086;
      end
    end else begin
      e_6_active_vlu <= _GEN_31086;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vsu <= _GEN_31078;
      end
    end else begin
      e_6_active_vsu <= _GEN_31078;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_6_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h6 == head) begin // @[sequencer-master.scala 373:43]
        e_6_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_6_active_vqu <= _GEN_31014;
      end
    end else begin
      e_6_active_vqu <= _GEN_31014;
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_0 <= _GEN_30532;
        end
      end else begin
        e_6_raw_0 <= _GEN_30532;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_1 <= _GEN_30556;
        end
      end else begin
        e_6_raw_1 <= _GEN_30556;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_2 <= _GEN_30580;
        end
      end else begin
        e_6_raw_2 <= _GEN_30580;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_3 <= _GEN_30604;
        end
      end else begin
        e_6_raw_3 <= _GEN_30604;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_4 <= _GEN_30628;
        end
      end else begin
        e_6_raw_4 <= _GEN_30628;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_5 <= _GEN_30652;
        end
      end else begin
        e_6_raw_5 <= _GEN_30652;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_6 <= _GEN_30676;
        end
      end else begin
        e_6_raw_6 <= _GEN_30676;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_6_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_6_raw_7 <= _GEN_30700;
        end
      end else begin
        e_6_raw_7 <= _GEN_30700;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_0 <= _GEN_30540;
        end
      end else begin
        e_6_war_0 <= _GEN_30540;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_1 <= _GEN_30564;
        end
      end else begin
        e_6_war_1 <= _GEN_30564;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_2 <= _GEN_30588;
        end
      end else begin
        e_6_war_2 <= _GEN_30588;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_3 <= _GEN_30612;
        end
      end else begin
        e_6_war_3 <= _GEN_30612;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_4 <= _GEN_30636;
        end
      end else begin
        e_6_war_4 <= _GEN_30636;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_5 <= _GEN_30660;
        end
      end else begin
        e_6_war_5 <= _GEN_30660;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_6 <= _GEN_30684;
        end
      end else begin
        e_6_war_6 <= _GEN_30684;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_6_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_6_war_7 <= _GEN_30708;
        end
      end else begin
        e_6_war_7 <= _GEN_30708;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_0 <= _GEN_30548;
        end
      end else begin
        e_6_waw_0 <= _GEN_30548;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_1 <= _GEN_30572;
        end
      end else begin
        e_6_waw_1 <= _GEN_30572;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_2 <= _GEN_30596;
        end
      end else begin
        e_6_waw_2 <= _GEN_30596;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_3 <= _GEN_30620;
        end
      end else begin
        e_6_waw_3 <= _GEN_30620;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_4 <= _GEN_30644;
        end
      end else begin
        e_6_waw_4 <= _GEN_30644;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_5 <= _GEN_30668;
        end
      end else begin
        e_6_waw_5 <= _GEN_30668;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_6 <= _GEN_30692;
        end
      end else begin
        e_6_waw_6 <= _GEN_30692;
      end
    end
    if (_GEN_32331) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_6_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_6_waw_7 <= _GEN_30716;
        end
      end else begin
        e_6_waw_7 <= _GEN_30716;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_6_last <= _GEN_31106;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_6_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_6_last <= _GEN_29202;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_6_last <= _GEN_27616;
      end else begin
        e_6_last <= _GEN_26118;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_6_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_6_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_6_rports <= _GEN_28922;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_6_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_6_rports <= _GEN_27080;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_rports <= _GEN_25774;
      end else begin
        e_6_rports <= _GEN_23892;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_6_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_6_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_6_wport_sram <= _GEN_28930;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_6_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_6_wport_sram <= _GEN_27088;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_wport_sram <= _GEN_25782;
      end else begin
        e_6_wport_sram <= _GEN_23900;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_6_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h6 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_6_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_6_wport_pred <= _GEN_28938;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h6 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_6_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_6_wport_pred <= _GEN_27096;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_6_wport_pred <= _GEN_25790;
      end else begin
        e_6_wport_pred <= _GEN_23908;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_7_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 289:23]
          e_7_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_7_fn_union <= _GEN_28707;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 289:23]
          e_7_fn_union <= io_op_bits_fn_union; // @[sequencer-master.scala 289:23]
        end else begin
          e_7_fn_union <= _GEN_27073;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_fn_union <= _GEN_25335;
      end else begin
        e_7_fn_union <= _GEN_23805;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_7_sreg_ss1 <= _GEN_24519;
          end else begin
            e_7_sreg_ss1 <= _GEN_23885;
          end
        end else begin
          e_7_sreg_ss1 <= _GEN_23885;
        end
      end else begin
        e_7_sreg_ss1 <= _GEN_23885;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_366) begin // @[sequencer-master.scala 331:55]
            e_7_sreg_ss2 <= _GEN_13531;
          end else begin
            e_7_sreg_ss2 <= _GEN_12657;
          end
        end else begin
          e_7_sreg_ss2 <= _GEN_12657;
        end
      end else begin
        e_7_sreg_ss2 <= _GEN_12657;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (_T_543) begin // @[sequencer-master.scala 331:55]
            e_7_sreg_ss3 <= _GEN_9175;
          end else begin
            e_7_sreg_ss3 <= _GEN_3753;
          end
        end else begin
          e_7_sreg_ss3 <= _GEN_3753;
        end
      end else begin
        e_7_sreg_ss3 <= _GEN_3753;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_7_base_vp_id <= io_op_bits_base_vp_id; // @[sequencer-master.scala 321:24]
          end else begin
            e_7_base_vp_id <= _GEN_28755;
          end
        end else begin
          e_7_base_vp_id <= _GEN_28755;
        end
      end else begin
        e_7_base_vp_id <= _GEN_28313;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_7_base_vp_valid <= io_op_bits_base_vp_valid; // @[sequencer-master.scala 321:24]
          end else begin
            e_7_base_vp_valid <= _GEN_29275;
          end
        end else begin
          e_7_base_vp_valid <= _GEN_29275;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 272:28]
          e_7_base_vp_valid <= 1'h0; // @[sequencer-master.scala 272:28]
        end else begin
          e_7_base_vp_valid <= _GEN_26809;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_base_vp_valid <= _GEN_25391;
      end else begin
        e_7_base_vp_valid <= _GEN_23541;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_7_base_vp_scalar <= io_op_bits_base_vp_scalar; // @[sequencer-master.scala 321:24]
          end else begin
            e_7_base_vp_scalar <= _GEN_28771;
          end
        end else begin
          e_7_base_vp_scalar <= _GEN_28771;
        end
      end else begin
        e_7_base_vp_scalar <= _GEN_28321;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vp_valid) begin // @[sequencer-master.scala 320:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 321:24]
            e_7_base_vp_pred <= io_op_bits_base_vp_pred; // @[sequencer-master.scala 321:24]
          end else begin
            e_7_base_vp_pred <= _GEN_28779;
          end
        end else begin
          e_7_base_vp_pred <= _GEN_28779;
        end
      end else begin
        e_7_base_vp_pred <= _GEN_28329;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_7_base_vs1_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 355:25]
          end else begin
            e_7_base_vs1_id <= _GEN_26183;
          end
        end else begin
          e_7_base_vs1_id <= _GEN_26183;
        end
      end else begin
        e_7_base_vs1_id <= _GEN_26183;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_7_base_vs1_valid <= io_op_bits_base_vd_valid; // @[sequencer-master.scala 355:25]
          end else begin
            e_7_base_vs1_valid <= _GEN_29283;
          end
        end else begin
          e_7_base_vs1_valid <= _GEN_29283;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 273:29]
          e_7_base_vs1_valid <= 1'h0; // @[sequencer-master.scala 273:29]
        end else begin
          e_7_base_vs1_valid <= _GEN_26817;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_base_vs1_valid <= _GEN_25607;
      end else begin
        e_7_base_vs1_valid <= _GEN_23549;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_7_base_vs1_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 355:25]
          end else begin
            e_7_base_vs1_scalar <= _GEN_26191;
          end
        end else begin
          e_7_base_vs1_scalar <= _GEN_26191;
        end
      end else begin
        e_7_base_vs1_scalar <= _GEN_26191;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_7_base_vs1_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 355:25]
          end else begin
            e_7_base_vs1_pred <= _GEN_26199;
          end
        end else begin
          e_7_base_vs1_pred <= _GEN_26199;
        end
      end else begin
        e_7_base_vs1_pred <= _GEN_26199;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 354:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 355:25]
            e_7_base_vs1_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 355:25]
          end else begin
            e_7_base_vs1_prec <= _GEN_26207;
          end
        end else begin
          e_7_base_vs1_prec <= _GEN_26207;
        end
      end else begin
        e_7_base_vs1_prec <= _GEN_26207;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs2_id <= io_op_bits_base_vs2_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs2_id <= _GEN_12617;
          end
        end else begin
          e_7_base_vs2_id <= _GEN_12617;
        end
      end else begin
        e_7_base_vs2_id <= _GEN_12617;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_7_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 274:29]
          e_7_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_7_base_vs2_valid <= _GEN_28459;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 274:29]
          e_7_base_vs2_valid <= 1'h0; // @[sequencer-master.scala 274:29]
        end else begin
          e_7_base_vs2_valid <= _GEN_26825;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_base_vs2_valid <= _GEN_25087;
      end else begin
        e_7_base_vs2_valid <= _GEN_23557;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs2_scalar <= io_op_bits_base_vs2_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs2_scalar <= _GEN_12625;
          end
        end else begin
          e_7_base_vs2_scalar <= _GEN_12625;
        end
      end else begin
        e_7_base_vs2_scalar <= _GEN_12625;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs2_pred <= io_op_bits_base_vs2_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs2_pred <= _GEN_12633;
          end
        end else begin
          e_7_base_vs2_pred <= _GEN_12633;
        end
      end else begin
        e_7_base_vs2_pred <= _GEN_12633;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfcmp) begin // @[sequencer-master.scala 646:40]
        if (io_op_bits_base_vs2_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs2_prec <= io_op_bits_base_vs2_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs2_prec <= _GEN_12641;
          end
        end else begin
          e_7_base_vs2_prec <= _GEN_12641;
        end
      end else begin
        e_7_base_vs2_prec <= _GEN_12641;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs3_id <= io_op_bits_base_vs3_id; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs3_id <= _GEN_3713;
          end
        end else begin
          e_7_base_vs3_id <= _GEN_3713;
        end
      end else begin
        e_7_base_vs3_id <= _GEN_3713;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_7_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 275:29]
          e_7_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_7_base_vs3_valid <= _GEN_28467;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 275:29]
          e_7_base_vs3_valid <= 1'h0; // @[sequencer-master.scala 275:29]
        end else begin
          e_7_base_vs3_valid <= _GEN_26833;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_base_vs3_valid <= _GEN_25095;
      end else begin
        e_7_base_vs3_valid <= _GEN_23565;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs3_scalar <= io_op_bits_base_vs3_scalar; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs3_scalar <= _GEN_3721;
          end
        end else begin
          e_7_base_vs3_scalar <= _GEN_3721;
        end
      end else begin
        e_7_base_vs3_scalar <= _GEN_3721;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs3_pred <= io_op_bits_base_vs3_pred; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs3_pred <= _GEN_3729;
          end
        end else begin
          e_7_base_vs3_pred <= _GEN_3729;
        end
      end else begin
        e_7_base_vs3_pred <= _GEN_3729;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vfma) begin // @[sequencer-master.scala 644:39]
        if (io_op_bits_base_vs3_valid) begin // @[sequencer-master.scala 328:47]
          if (3'h7 == tail) begin // @[sequencer-master.scala 329:29]
            e_7_base_vs3_prec <= io_op_bits_base_vs3_prec; // @[sequencer-master.scala 329:29]
          end else begin
            e_7_base_vs3_prec <= _GEN_3737;
          end
        end else begin
          e_7_base_vs3_prec <= _GEN_3737;
        end
      end else begin
        e_7_base_vs3_prec <= _GEN_3737;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_7_base_vd_id <= io_op_bits_base_vd_id; // @[sequencer-master.scala 363:24]
          end else begin
            e_7_base_vd_id <= _GEN_23933;
          end
        end else begin
          e_7_base_vd_id <= _GEN_23933;
        end
      end else begin
        e_7_base_vd_id <= _GEN_23933;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 276:28]
          e_7_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 276:28]
          e_7_base_vd_valid <= 1'h0; // @[sequencer-master.scala 276:28]
        end else begin
          e_7_base_vd_valid <= _GEN_28475;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          e_7_base_vd_valid <= _GEN_27657;
        end else begin
          e_7_base_vd_valid <= _GEN_27409;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_base_vd_valid <= _GEN_25103;
      end else begin
        e_7_base_vd_valid <= _GEN_23573;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_7_base_vd_scalar <= io_op_bits_base_vd_scalar; // @[sequencer-master.scala 363:24]
          end else begin
            e_7_base_vd_scalar <= _GEN_23941;
          end
        end else begin
          e_7_base_vd_scalar <= _GEN_23941;
        end
      end else begin
        e_7_base_vd_scalar <= _GEN_23941;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_7_base_vd_pred <= io_op_bits_base_vd_pred; // @[sequencer-master.scala 363:24]
          end else begin
            e_7_base_vd_pred <= _GEN_23949;
          end
        end else begin
          e_7_base_vd_pred <= _GEN_23949;
        end
      end else begin
        e_7_base_vd_pred <= _GEN_23949;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (io_op_bits_base_vd_valid) begin // @[sequencer-master.scala 362:41]
          if (3'h7 == _T_1647) begin // @[sequencer-master.scala 363:24]
            e_7_base_vd_prec <= io_op_bits_base_vd_prec; // @[sequencer-master.scala 363:24]
          end else begin
            e_7_base_vd_prec <= _GEN_23957;
          end
        end else begin
          e_7_base_vd_prec <= _GEN_23957;
        end
      end else begin
        e_7_base_vd_prec <= _GEN_23957;
      end
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_viu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_viu <= _GEN_30741;
      end
    end else begin
      e_7_active_viu <= _GEN_30741;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vipu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vipu <= _GEN_30951;
      end
    end else begin
      e_7_active_vipu <= _GEN_30951;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vimu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vimu <= _GEN_31007;
      end
    end else begin
      e_7_active_vimu <= _GEN_31007;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vidu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vidu <= _GEN_31023;
      end
    end else begin
      e_7_active_vidu <= _GEN_31023;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vfmu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vfmu <= _GEN_31031;
      end
    end else begin
      e_7_active_vfmu <= _GEN_31031;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vfdu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vfdu <= _GEN_31039;
      end
    end else begin
      e_7_active_vfdu <= _GEN_31039;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vfcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vfcu <= _GEN_31047;
      end
    end else begin
      e_7_active_vfcu <= _GEN_31047;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vfvu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vfvu <= _GEN_31055;
      end
    end else begin
      e_7_active_vfvu <= _GEN_31055;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vpu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vpu <= _GEN_31095;
      end
    end else begin
      e_7_active_vpu <= _GEN_31095;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vgu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vgu <= _GEN_31063;
      end
    end else begin
      e_7_active_vgu <= _GEN_31063;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vcu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vcu <= _GEN_31071;
      end
    end else begin
      e_7_active_vcu <= _GEN_31071;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vlu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vlu <= _GEN_31087;
      end
    end else begin
      e_7_active_vlu <= _GEN_31087;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vsu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vsu <= _GEN_31079;
      end
    end else begin
      e_7_active_vsu <= _GEN_31079;
    end
    if (reset) begin // @[sequencer-master.scala 468:20]
      e_7_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
    end else if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      if (3'h7 == head) begin // @[sequencer-master.scala 373:43]
        e_7_active_vqu <= 1'h0; // @[sequencer-master.scala 373:43]
      end else begin
        e_7_active_vqu <= _GEN_31015;
      end
    end else begin
      e_7_active_vqu <= _GEN_31015;
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_0 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_0 <= _GEN_30533;
        end
      end else begin
        e_7_raw_0 <= _GEN_30533;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_1 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_1 <= _GEN_30557;
        end
      end else begin
        e_7_raw_1 <= _GEN_30557;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_2 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_2 <= _GEN_30581;
        end
      end else begin
        e_7_raw_2 <= _GEN_30581;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_3 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_3 <= _GEN_30605;
        end
      end else begin
        e_7_raw_3 <= _GEN_30605;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_4 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_4 <= _GEN_30629;
        end
      end else begin
        e_7_raw_4 <= _GEN_30629;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_5 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_5 <= _GEN_30653;
        end
      end else begin
        e_7_raw_5 <= _GEN_30653;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_6 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_6 <= _GEN_30677;
        end
      end else begin
        e_7_raw_6 <= _GEN_30677;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 183:52]
          e_7_raw_7 <= 1'h0; // @[sequencer-master.scala 183:52]
        end else begin
          e_7_raw_7 <= _GEN_30701;
        end
      end else begin
        e_7_raw_7 <= _GEN_30701;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_0 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_0 <= _GEN_30541;
        end
      end else begin
        e_7_war_0 <= _GEN_30541;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_1 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_1 <= _GEN_30565;
        end
      end else begin
        e_7_war_1 <= _GEN_30565;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_2 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_2 <= _GEN_30589;
        end
      end else begin
        e_7_war_2 <= _GEN_30589;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_3 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_3 <= _GEN_30613;
        end
      end else begin
        e_7_war_3 <= _GEN_30613;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_4 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_4 <= _GEN_30637;
        end
      end else begin
        e_7_war_4 <= _GEN_30637;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_5 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_5 <= _GEN_30661;
        end
      end else begin
        e_7_war_5 <= _GEN_30661;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_6 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_6 <= _GEN_30685;
        end
      end else begin
        e_7_war_6 <= _GEN_30685;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 184:52]
          e_7_war_7 <= 1'h0; // @[sequencer-master.scala 184:52]
        end else begin
          e_7_war_7 <= _GEN_30709;
        end
      end else begin
        e_7_war_7 <= _GEN_30709;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h0 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_0 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_0 <= _GEN_30549;
        end
      end else begin
        e_7_waw_0 <= _GEN_30549;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h1 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_1 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_1 <= _GEN_30573;
        end
      end else begin
        e_7_waw_1 <= _GEN_30573;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h2 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_2 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_2 <= _GEN_30597;
        end
      end else begin
        e_7_waw_2 <= _GEN_30597;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h3 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_3 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_3 <= _GEN_30621;
        end
      end else begin
        e_7_waw_3 <= _GEN_30621;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h4 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_4 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_4 <= _GEN_30645;
        end
      end else begin
        e_7_waw_4 <= _GEN_30645;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h5 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_5 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_5 <= _GEN_30669;
        end
      end else begin
        e_7_waw_5 <= _GEN_30669;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h6 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_6 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_6 <= _GEN_30693;
        end
      end else begin
        e_7_waw_6 <= _GEN_30693;
      end
    end
    if (_GEN_32356) begin // @[sequencer-master.scala 203:31]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        if (3'h7 == head) begin // @[sequencer-master.scala 185:52]
          e_7_waw_7 <= 1'h0; // @[sequencer-master.scala 185:52]
        end else begin
          e_7_waw_7 <= _GEN_30717;
        end
      end else begin
        e_7_waw_7 <= _GEN_30717;
      end
    end
    if (io_vf_stop) begin // @[sequencer-master.scala 433:25]
      e_7_last <= _GEN_31107;
    end else if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 283:19]
          e_7_last <= 1'h0; // @[sequencer-master.scala 283:19]
        end else begin
          e_7_last <= _GEN_29203;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        e_7_last <= _GEN_27617;
      end else begin
        e_7_last <= _GEN_26119;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_7_rports <= _e_T_1647_rports_1; // @[sequencer-master.scala 230:21]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 230:21]
          e_7_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_7_rports <= _GEN_28923;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 230:21]
          e_7_rports <= 2'h0; // @[sequencer-master.scala 230:21]
        end else begin
          e_7_rports <= _GEN_27081;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_rports <= _GEN_25775;
      end else begin
        e_7_rports <= _GEN_23893;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_7_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 231:25]
          e_7_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_7_wport_sram <= _GEN_28931;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 231:25]
          e_7_wport_sram <= 4'h0; // @[sequencer-master.scala 231:25]
        end else begin
          e_7_wport_sram <= _GEN_27089;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_wport_sram <= _GEN_25783;
      end else begin
        e_7_wport_sram <= _GEN_23901;
      end
    end
    if (_T_1752) begin // @[sequencer-master.scala 639:27]
      if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_7_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else if (3'h7 == _T_1645) begin // @[sequencer-master.scala 232:25]
          e_7_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_7_wport_pred <= _GEN_28939;
        end
      end else if (io_op_bits_active_vld) begin // @[sequencer-master.scala 653:38]
        if (3'h7 == _T_1647) begin // @[sequencer-master.scala 232:25]
          e_7_wport_pred <= 3'h0; // @[sequencer-master.scala 232:25]
        end else begin
          e_7_wport_pred <= _GEN_27097;
        end
      end else if (io_op_bits_active_vstx) begin // @[sequencer-master.scala 652:39]
        e_7_wport_pred <= _GEN_25791;
      end else begin
        e_7_wport_pred <= _GEN_23909;
      end
    end
    if (reset) begin // @[sequencer-master.scala 111:23]
      maybe_full <= 1'h0; // @[sequencer-master.scala 111:23]
    end else if (_T_2443) begin // @[sequencer-master.scala 422:26]
      maybe_full <= 1'h0; // @[sequencer-master.scala 424:20]
    end else begin
      maybe_full <= _GEN_31097;
    end
    if (reset) begin // @[sequencer-master.scala 112:17]
      head <= 3'h0; // @[sequencer-master.scala 112:17]
    end else if (_T_2443) begin // @[sequencer-master.scala 422:26]
      if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
        head <= _T_2440; // @[sequencer-master.scala 264:66]
      end
    end
    if (reset) begin // @[sequencer-master.scala 113:17]
      tail <= 3'h0; // @[sequencer-master.scala 113:17]
    end else if (_GEN_30942) begin // @[sequencer-master.scala 418:26]
      if (_T_1752) begin // @[sequencer-master.scala 639:27]
        if (io_op_bits_active_vst) begin // @[sequencer-master.scala 654:38]
          tail <= _T_1649; // @[sequencer-master.scala 265:66]
        end else begin
          tail <= _GEN_28419;
        end
      end
    end
    if (_GEN_31124 & _GEN_31132) begin // @[sequencer-master.scala 438:47]
      _T_2465 <= _GEN_32041 | io_vf_stop & _T_2440 == tail; // @[sequencer-master.scala 441:17]
    end else begin
      _T_2465 <= _GEN_31116;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vint & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vint & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vipred & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vipred & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vimul & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vimul & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vidiv & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n"
            ); // @[sequencer-master.scala 298:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vidiv & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fatal; // @[sequencer-master.scala 298:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_38872 & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_38872 & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfma & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfma & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfdiv & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n"
            ); // @[sequencer-master.scala 298:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfdiv & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fatal; // @[sequencer-master.scala 298:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_38878 & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_38878 & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfcmp & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfcmp & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfconv & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vfconv & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vrpred & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n"
            ); // @[sequencer-master.scala 298:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vrpred & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fatal; // @[sequencer-master.scala 298:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vrfirst & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n"
            ); // @[sequencer-master.scala 298:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vrfirst & ~(io_op_bits_active_vidiv | io_op_bits_active_vfdiv |
          io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset)) begin
          $fatal; // @[sequencer-master.scala 298:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vamo & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vamo & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vldx & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vldx & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vstx & _T_1764) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd_as_vs1: vd should always be vector\n    at sequencer-master.scala:353 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd_as_vs1: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 353:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vstx & _T_1764) begin
          $fatal; // @[sequencer-master.scala 353:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vld & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 361:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vld & ~(~io_op_bits_base_vd_valid | _T_721 | reset)) begin
          $fatal; // @[sequencer-master.scala 361:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vst & _T_1764) begin
          $fwrite(32'h80000002,
            "Assertion failed: iwindow.set.vd_as_vs1: vd should always be vector\n    at sequencer-master.scala:353 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd_as_vs1: vd should always be vector\")\n"
            ); // @[sequencer-master.scala 353:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1752 & io_op_bits_active_vst & _T_1764) begin
          $fatal; // @[sequencer-master.scala 353:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  v_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  v_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  v_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  v_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  v_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  v_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  v_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  v_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  e_0_fn_union = _RAND_8[9:0];
  _RAND_9 = {2{`RANDOM}};
  e_0_sreg_ss1 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  e_0_sreg_ss2 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  e_0_sreg_ss3 = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  e_0_base_vp_id = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  e_0_base_vp_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  e_0_base_vp_scalar = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  e_0_base_vp_pred = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  e_0_base_vs1_id = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  e_0_base_vs1_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  e_0_base_vs1_scalar = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  e_0_base_vs1_pred = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  e_0_base_vs1_prec = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  e_0_base_vs2_id = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  e_0_base_vs2_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  e_0_base_vs2_scalar = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  e_0_base_vs2_pred = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  e_0_base_vs2_prec = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  e_0_base_vs3_id = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  e_0_base_vs3_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  e_0_base_vs3_scalar = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  e_0_base_vs3_pred = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  e_0_base_vs3_prec = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  e_0_base_vd_id = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  e_0_base_vd_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  e_0_base_vd_scalar = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  e_0_base_vd_pred = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  e_0_base_vd_prec = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  e_0_active_viu = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  e_0_active_vipu = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  e_0_active_vimu = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  e_0_active_vidu = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  e_0_active_vfmu = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  e_0_active_vfdu = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  e_0_active_vfcu = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  e_0_active_vfvu = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  e_0_active_vpu = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  e_0_active_vgu = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  e_0_active_vcu = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  e_0_active_vlu = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  e_0_active_vsu = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  e_0_active_vqu = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  e_0_raw_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  e_0_raw_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  e_0_raw_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  e_0_raw_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  e_0_raw_4 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  e_0_raw_5 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  e_0_raw_6 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  e_0_raw_7 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  e_0_war_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  e_0_war_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  e_0_war_2 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  e_0_war_3 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  e_0_war_4 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  e_0_war_5 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  e_0_war_6 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  e_0_war_7 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  e_0_waw_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  e_0_waw_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  e_0_waw_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  e_0_waw_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  e_0_waw_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  e_0_waw_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  e_0_waw_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  e_0_waw_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  e_0_last = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  e_0_rports = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  e_0_wport_sram = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  e_0_wport_pred = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  e_1_fn_union = _RAND_78[9:0];
  _RAND_79 = {2{`RANDOM}};
  e_1_sreg_ss1 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  e_1_sreg_ss2 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  e_1_sreg_ss3 = _RAND_81[63:0];
  _RAND_82 = {1{`RANDOM}};
  e_1_base_vp_id = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  e_1_base_vp_valid = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  e_1_base_vp_scalar = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  e_1_base_vp_pred = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  e_1_base_vs1_id = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  e_1_base_vs1_valid = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  e_1_base_vs1_scalar = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  e_1_base_vs1_pred = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  e_1_base_vs1_prec = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  e_1_base_vs2_id = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  e_1_base_vs2_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  e_1_base_vs2_scalar = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  e_1_base_vs2_pred = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  e_1_base_vs2_prec = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  e_1_base_vs3_id = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  e_1_base_vs3_valid = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  e_1_base_vs3_scalar = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  e_1_base_vs3_pred = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  e_1_base_vs3_prec = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  e_1_base_vd_id = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  e_1_base_vd_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  e_1_base_vd_scalar = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  e_1_base_vd_pred = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  e_1_base_vd_prec = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  e_1_active_viu = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  e_1_active_vipu = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  e_1_active_vimu = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  e_1_active_vidu = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  e_1_active_vfmu = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  e_1_active_vfdu = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  e_1_active_vfcu = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  e_1_active_vfvu = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  e_1_active_vpu = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  e_1_active_vgu = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  e_1_active_vcu = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  e_1_active_vlu = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  e_1_active_vsu = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  e_1_active_vqu = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  e_1_raw_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  e_1_raw_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  e_1_raw_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  e_1_raw_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  e_1_raw_4 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  e_1_raw_5 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  e_1_raw_6 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  e_1_raw_7 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  e_1_war_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  e_1_war_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  e_1_war_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  e_1_war_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  e_1_war_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  e_1_war_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  e_1_war_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  e_1_war_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  e_1_waw_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  e_1_waw_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  e_1_waw_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  e_1_waw_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  e_1_waw_4 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  e_1_waw_5 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  e_1_waw_6 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  e_1_waw_7 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  e_1_last = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  e_1_rports = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  e_1_wport_sram = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  e_1_wport_pred = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  e_2_fn_union = _RAND_148[9:0];
  _RAND_149 = {2{`RANDOM}};
  e_2_sreg_ss1 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  e_2_sreg_ss2 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  e_2_sreg_ss3 = _RAND_151[63:0];
  _RAND_152 = {1{`RANDOM}};
  e_2_base_vp_id = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  e_2_base_vp_valid = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  e_2_base_vp_scalar = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  e_2_base_vp_pred = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  e_2_base_vs1_id = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  e_2_base_vs1_valid = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  e_2_base_vs1_scalar = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  e_2_base_vs1_pred = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  e_2_base_vs1_prec = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  e_2_base_vs2_id = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  e_2_base_vs2_valid = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  e_2_base_vs2_scalar = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  e_2_base_vs2_pred = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  e_2_base_vs2_prec = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  e_2_base_vs3_id = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  e_2_base_vs3_valid = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  e_2_base_vs3_scalar = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  e_2_base_vs3_pred = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  e_2_base_vs3_prec = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  e_2_base_vd_id = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  e_2_base_vd_valid = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  e_2_base_vd_scalar = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  e_2_base_vd_pred = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  e_2_base_vd_prec = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  e_2_active_viu = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  e_2_active_vipu = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  e_2_active_vimu = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  e_2_active_vidu = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  e_2_active_vfmu = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  e_2_active_vfdu = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  e_2_active_vfcu = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  e_2_active_vfvu = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  e_2_active_vpu = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  e_2_active_vgu = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  e_2_active_vcu = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  e_2_active_vlu = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  e_2_active_vsu = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  e_2_active_vqu = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  e_2_raw_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  e_2_raw_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  e_2_raw_2 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  e_2_raw_3 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  e_2_raw_4 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  e_2_raw_5 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  e_2_raw_6 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  e_2_raw_7 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  e_2_war_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  e_2_war_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  e_2_war_2 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  e_2_war_3 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  e_2_war_4 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  e_2_war_5 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  e_2_war_6 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  e_2_war_7 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  e_2_waw_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  e_2_waw_1 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  e_2_waw_2 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  e_2_waw_3 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  e_2_waw_4 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  e_2_waw_5 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  e_2_waw_6 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  e_2_waw_7 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  e_2_last = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  e_2_rports = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  e_2_wport_sram = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  e_2_wport_pred = _RAND_217[2:0];
  _RAND_218 = {1{`RANDOM}};
  e_3_fn_union = _RAND_218[9:0];
  _RAND_219 = {2{`RANDOM}};
  e_3_sreg_ss1 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  e_3_sreg_ss2 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  e_3_sreg_ss3 = _RAND_221[63:0];
  _RAND_222 = {1{`RANDOM}};
  e_3_base_vp_id = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  e_3_base_vp_valid = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  e_3_base_vp_scalar = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  e_3_base_vp_pred = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  e_3_base_vs1_id = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  e_3_base_vs1_valid = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  e_3_base_vs1_scalar = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  e_3_base_vs1_pred = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  e_3_base_vs1_prec = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  e_3_base_vs2_id = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  e_3_base_vs2_valid = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  e_3_base_vs2_scalar = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  e_3_base_vs2_pred = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  e_3_base_vs2_prec = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  e_3_base_vs3_id = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  e_3_base_vs3_valid = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  e_3_base_vs3_scalar = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  e_3_base_vs3_pred = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  e_3_base_vs3_prec = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  e_3_base_vd_id = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  e_3_base_vd_valid = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  e_3_base_vd_scalar = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  e_3_base_vd_pred = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  e_3_base_vd_prec = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  e_3_active_viu = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  e_3_active_vipu = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  e_3_active_vimu = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  e_3_active_vidu = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  e_3_active_vfmu = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  e_3_active_vfdu = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  e_3_active_vfcu = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  e_3_active_vfvu = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  e_3_active_vpu = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  e_3_active_vgu = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  e_3_active_vcu = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  e_3_active_vlu = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  e_3_active_vsu = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  e_3_active_vqu = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  e_3_raw_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  e_3_raw_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  e_3_raw_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  e_3_raw_3 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  e_3_raw_4 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  e_3_raw_5 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  e_3_raw_6 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  e_3_raw_7 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  e_3_war_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  e_3_war_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  e_3_war_2 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  e_3_war_3 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  e_3_war_4 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  e_3_war_5 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  e_3_war_6 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  e_3_war_7 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  e_3_waw_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  e_3_waw_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  e_3_waw_2 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  e_3_waw_3 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  e_3_waw_4 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  e_3_waw_5 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  e_3_waw_6 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  e_3_waw_7 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  e_3_last = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  e_3_rports = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  e_3_wport_sram = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  e_3_wport_pred = _RAND_287[2:0];
  _RAND_288 = {1{`RANDOM}};
  e_4_fn_union = _RAND_288[9:0];
  _RAND_289 = {2{`RANDOM}};
  e_4_sreg_ss1 = _RAND_289[63:0];
  _RAND_290 = {2{`RANDOM}};
  e_4_sreg_ss2 = _RAND_290[63:0];
  _RAND_291 = {2{`RANDOM}};
  e_4_sreg_ss3 = _RAND_291[63:0];
  _RAND_292 = {1{`RANDOM}};
  e_4_base_vp_id = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  e_4_base_vp_valid = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  e_4_base_vp_scalar = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  e_4_base_vp_pred = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  e_4_base_vs1_id = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  e_4_base_vs1_valid = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  e_4_base_vs1_scalar = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  e_4_base_vs1_pred = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  e_4_base_vs1_prec = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  e_4_base_vs2_id = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  e_4_base_vs2_valid = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  e_4_base_vs2_scalar = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  e_4_base_vs2_pred = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  e_4_base_vs2_prec = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  e_4_base_vs3_id = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  e_4_base_vs3_valid = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  e_4_base_vs3_scalar = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  e_4_base_vs3_pred = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  e_4_base_vs3_prec = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  e_4_base_vd_id = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  e_4_base_vd_valid = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  e_4_base_vd_scalar = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  e_4_base_vd_pred = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  e_4_base_vd_prec = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  e_4_active_viu = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  e_4_active_vipu = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  e_4_active_vimu = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  e_4_active_vidu = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  e_4_active_vfmu = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  e_4_active_vfdu = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  e_4_active_vfcu = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  e_4_active_vfvu = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  e_4_active_vpu = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  e_4_active_vgu = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  e_4_active_vcu = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  e_4_active_vlu = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  e_4_active_vsu = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  e_4_active_vqu = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  e_4_raw_0 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  e_4_raw_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  e_4_raw_2 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  e_4_raw_3 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  e_4_raw_4 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  e_4_raw_5 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  e_4_raw_6 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  e_4_raw_7 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  e_4_war_0 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  e_4_war_1 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  e_4_war_2 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  e_4_war_3 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  e_4_war_4 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  e_4_war_5 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  e_4_war_6 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  e_4_war_7 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  e_4_waw_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  e_4_waw_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  e_4_waw_2 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  e_4_waw_3 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  e_4_waw_4 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  e_4_waw_5 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  e_4_waw_6 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  e_4_waw_7 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  e_4_last = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  e_4_rports = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  e_4_wport_sram = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  e_4_wport_pred = _RAND_357[2:0];
  _RAND_358 = {1{`RANDOM}};
  e_5_fn_union = _RAND_358[9:0];
  _RAND_359 = {2{`RANDOM}};
  e_5_sreg_ss1 = _RAND_359[63:0];
  _RAND_360 = {2{`RANDOM}};
  e_5_sreg_ss2 = _RAND_360[63:0];
  _RAND_361 = {2{`RANDOM}};
  e_5_sreg_ss3 = _RAND_361[63:0];
  _RAND_362 = {1{`RANDOM}};
  e_5_base_vp_id = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  e_5_base_vp_valid = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  e_5_base_vp_scalar = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  e_5_base_vp_pred = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  e_5_base_vs1_id = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  e_5_base_vs1_valid = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  e_5_base_vs1_scalar = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  e_5_base_vs1_pred = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  e_5_base_vs1_prec = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  e_5_base_vs2_id = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  e_5_base_vs2_valid = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  e_5_base_vs2_scalar = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  e_5_base_vs2_pred = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  e_5_base_vs2_prec = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  e_5_base_vs3_id = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  e_5_base_vs3_valid = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  e_5_base_vs3_scalar = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  e_5_base_vs3_pred = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  e_5_base_vs3_prec = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  e_5_base_vd_id = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  e_5_base_vd_valid = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  e_5_base_vd_scalar = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  e_5_base_vd_pred = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  e_5_base_vd_prec = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  e_5_active_viu = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  e_5_active_vipu = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  e_5_active_vimu = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  e_5_active_vidu = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  e_5_active_vfmu = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  e_5_active_vfdu = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  e_5_active_vfcu = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  e_5_active_vfvu = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  e_5_active_vpu = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  e_5_active_vgu = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  e_5_active_vcu = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  e_5_active_vlu = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  e_5_active_vsu = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  e_5_active_vqu = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  e_5_raw_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  e_5_raw_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  e_5_raw_2 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  e_5_raw_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  e_5_raw_4 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  e_5_raw_5 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  e_5_raw_6 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  e_5_raw_7 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  e_5_war_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  e_5_war_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  e_5_war_2 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  e_5_war_3 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  e_5_war_4 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  e_5_war_5 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  e_5_war_6 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  e_5_war_7 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  e_5_waw_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  e_5_waw_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  e_5_waw_2 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  e_5_waw_3 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  e_5_waw_4 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  e_5_waw_5 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  e_5_waw_6 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  e_5_waw_7 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  e_5_last = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  e_5_rports = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  e_5_wport_sram = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  e_5_wport_pred = _RAND_427[2:0];
  _RAND_428 = {1{`RANDOM}};
  e_6_fn_union = _RAND_428[9:0];
  _RAND_429 = {2{`RANDOM}};
  e_6_sreg_ss1 = _RAND_429[63:0];
  _RAND_430 = {2{`RANDOM}};
  e_6_sreg_ss2 = _RAND_430[63:0];
  _RAND_431 = {2{`RANDOM}};
  e_6_sreg_ss3 = _RAND_431[63:0];
  _RAND_432 = {1{`RANDOM}};
  e_6_base_vp_id = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  e_6_base_vp_valid = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  e_6_base_vp_scalar = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  e_6_base_vp_pred = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  e_6_base_vs1_id = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  e_6_base_vs1_valid = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  e_6_base_vs1_scalar = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  e_6_base_vs1_pred = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  e_6_base_vs1_prec = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  e_6_base_vs2_id = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  e_6_base_vs2_valid = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  e_6_base_vs2_scalar = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  e_6_base_vs2_pred = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  e_6_base_vs2_prec = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  e_6_base_vs3_id = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  e_6_base_vs3_valid = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  e_6_base_vs3_scalar = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  e_6_base_vs3_pred = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  e_6_base_vs3_prec = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  e_6_base_vd_id = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  e_6_base_vd_valid = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  e_6_base_vd_scalar = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  e_6_base_vd_pred = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  e_6_base_vd_prec = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  e_6_active_viu = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  e_6_active_vipu = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  e_6_active_vimu = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  e_6_active_vidu = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  e_6_active_vfmu = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  e_6_active_vfdu = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  e_6_active_vfcu = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  e_6_active_vfvu = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  e_6_active_vpu = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  e_6_active_vgu = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  e_6_active_vcu = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  e_6_active_vlu = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  e_6_active_vsu = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  e_6_active_vqu = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  e_6_raw_0 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  e_6_raw_1 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  e_6_raw_2 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  e_6_raw_3 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  e_6_raw_4 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  e_6_raw_5 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  e_6_raw_6 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  e_6_raw_7 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  e_6_war_0 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  e_6_war_1 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  e_6_war_2 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  e_6_war_3 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  e_6_war_4 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  e_6_war_5 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  e_6_war_6 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  e_6_war_7 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  e_6_waw_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  e_6_waw_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  e_6_waw_2 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  e_6_waw_3 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  e_6_waw_4 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  e_6_waw_5 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  e_6_waw_6 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  e_6_waw_7 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  e_6_last = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  e_6_rports = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  e_6_wport_sram = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  e_6_wport_pred = _RAND_497[2:0];
  _RAND_498 = {1{`RANDOM}};
  e_7_fn_union = _RAND_498[9:0];
  _RAND_499 = {2{`RANDOM}};
  e_7_sreg_ss1 = _RAND_499[63:0];
  _RAND_500 = {2{`RANDOM}};
  e_7_sreg_ss2 = _RAND_500[63:0];
  _RAND_501 = {2{`RANDOM}};
  e_7_sreg_ss3 = _RAND_501[63:0];
  _RAND_502 = {1{`RANDOM}};
  e_7_base_vp_id = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  e_7_base_vp_valid = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  e_7_base_vp_scalar = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  e_7_base_vp_pred = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  e_7_base_vs1_id = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  e_7_base_vs1_valid = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  e_7_base_vs1_scalar = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  e_7_base_vs1_pred = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  e_7_base_vs1_prec = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  e_7_base_vs2_id = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  e_7_base_vs2_valid = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  e_7_base_vs2_scalar = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  e_7_base_vs2_pred = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  e_7_base_vs2_prec = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  e_7_base_vs3_id = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  e_7_base_vs3_valid = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  e_7_base_vs3_scalar = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  e_7_base_vs3_pred = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  e_7_base_vs3_prec = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  e_7_base_vd_id = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  e_7_base_vd_valid = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  e_7_base_vd_scalar = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  e_7_base_vd_pred = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  e_7_base_vd_prec = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  e_7_active_viu = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  e_7_active_vipu = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  e_7_active_vimu = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  e_7_active_vidu = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  e_7_active_vfmu = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  e_7_active_vfdu = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  e_7_active_vfcu = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  e_7_active_vfvu = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  e_7_active_vpu = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  e_7_active_vgu = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  e_7_active_vcu = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  e_7_active_vlu = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  e_7_active_vsu = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  e_7_active_vqu = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  e_7_raw_0 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  e_7_raw_1 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  e_7_raw_2 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  e_7_raw_3 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  e_7_raw_4 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  e_7_raw_5 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  e_7_raw_6 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  e_7_raw_7 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  e_7_war_0 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  e_7_war_1 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  e_7_war_2 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  e_7_war_3 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  e_7_war_4 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  e_7_war_5 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  e_7_war_6 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  e_7_war_7 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  e_7_waw_0 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  e_7_waw_1 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  e_7_waw_2 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  e_7_waw_3 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  e_7_waw_4 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  e_7_waw_5 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  e_7_waw_6 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  e_7_waw_7 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  e_7_last = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  e_7_rports = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  e_7_wport_sram = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  e_7_wport_pred = _RAND_567[2:0];
  _RAND_568 = {1{`RANDOM}};
  maybe_full = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  head = _RAND_569[2:0];
  _RAND_570 = {1{`RANDOM}};
  tail = _RAND_570[2:0];
  _RAND_571 = {1{`RANDOM}};
  _T_2465 = _RAND_571[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
